`define INPUT_BITWIDTH 8
`define BITWIDTH 16
`define NUM_CYCLE 2
`define LOG_NUM_CYCLE 2
`define SIZE 100
`define NUMBER_UNIT 1
`define INST_BITWIDTH 3

`define SVM 1
//`define LINEAR 1
//`define LOGISTIC 1
//`define RECO 1
