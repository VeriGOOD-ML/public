
`timescale 1ns/1ps
module instruction_memory #(
    parameter integer addrLen = 5,
    parameter integer dataLen = 32,
    parameter integer peId  = 1
)(
    input clk,
    input rstn,
    
    input stall,
    input start,
    input restart,
    
    output reg [dataLen - 1: 0] data_out
);
//--------------------------------------------------------------------------------------
//reg [dataLen - 1: 0] mem  [0: (1 << addrLen) - 1];
reg [addrLen-1:0]        address;
reg enable;
reg [dataLen - 1: 0] rdata;
wire end_of_instruction;
always @(posedge clk or negedge rstn)
    if(~rstn)
        enable <= 1'b0;
    else if(start)
        enable <= 1'b1;
    else if(end_of_instruction)
       enable <= 1'b0;
always @(posedge clk or negedge rstn) begin
    if(~rstn)
        address <= {addrLen{1'b0}};
    else begin
        if(end_of_instruction)
            address <= {addrLen{1'b0}};
        else if(~stall && enable )
            address <= address + {{addrLen-1{1'b0}},1'b1};   
    end     
end
always @(posedge clk or negedge rstn) begin
    if(~rstn)
        data_out <= {1'b1,{dataLen-1{1'b0}}};
    else if((~stall && enable && ~end_of_instruction)||(end_of_instruction && start))
       data_out <= rdata;
end
    
assign end_of_instruction = (data_out[dataLen-1:dataLen-5] == 5'b0);
/****************************************************************************/
generate
if(peId == 0) begin
	always @(*) begin
		case(address)
			// PEs: 7 -> 8
			// srcs: (3, 0)(412) 3 --> (412) 3:PENB, pass, PUNB
			8'd0 : rdata = 43'b1100011011111110000000000000000001000000000;
			// PEs: 7 -> 8
			// srcs: (4, 1)(490) -4 --> (490) -4:PENB, pass, PUNB
			8'd1 : rdata = 43'b1100011011111110000000000000000001000000000;
			// PEs: 7 -> 8
			// srcs: (5, 2)(568) -1 --> (568) -1:PENB, pass, PUNB
			8'd2 : rdata = 43'b1100011011111110000000000000000001000000000;
			// PEs: 7 -> 24
			// srcs: (6, 16)(517) 0 --> (517) 0:PENB, pass, PUGB3
			8'd3 : rdata = 43'b1100011011111110000000000000000000000001011;
			// PEs: 1 -> 8
			// srcs: (9, 10)(495) -1 --> (495) -1:PEGB1, pass, PUNB
			8'd4 : rdata = 43'b1100011100000010000000000000000001000000000;
			// PEs: 2 -> 8
			// srcs: (10, 11)(498) 4 --> (498) 4:PEGB2, pass, PUNB
			8'd5 : rdata = 43'b1100011100000100000000000000000001000000000;
			// PEs: 4 -> 40
			// srcs: (11, 13)(504) 2 --> (504) 2:PEGB4, pass, PUGB5
			8'd6 : rdata = 43'b1100011100001000000000000000000000000001101;
			// PEs: 5 -> 56
			// srcs: (12, 14)(511) 4 --> (511) 4:PEGB5, pass, PUGB7
			8'd7 : rdata = 43'b1100011100001010000000000000000000000001111;
			// PEs: 6 -> 16
			// srcs: (13, 15)(514) -4 --> (514) -4:PEGB6, pass, PUGB2
			8'd8 : rdata = 43'b1100011100001100000000000000000000000001010;
			// PEs: 1 -> 48
			// srcs: (14, 3)(608) -4 --> (608) -4:PEGB1, pass, PUGB6
			8'd9 : rdata = 43'b1100011100000010000000000000000000000001110;
			// PEs: 4 -> 56
			// srcs: (15, 18)(759) 2 --> (759) 2:PEGB4, pass, PUGB7
			8'd10 : rdata = 43'b1100011100001000000000000000000000000001111;
			// PEs: 40 -> 0
			// srcs: (16, 5)(436) -1 --> (436) -1:PUGB5, pass, NI0
			8'd11 : rdata = 43'b1100011100001011000000000001000000000000000;
			// PEs: 7 -> 48
			// srcs: (17, 20)(607) -2 --> (607) -2:PENB, pass, PUGB6
			8'd12 : rdata = 43'b1100011011111110000000000000000000000001110;
			// PEs: 24 -> 1
			// srcs: (19, 4)(632) 2 --> (632) 2:PUGB3, pass, PENB
			8'd13 : rdata = 43'b1100011100000111000000000000000000100000000;
			// PEs: 0 -> 1
			// srcs: (26, 6)(436) -1 --> (436) -1:NI0, pass, PENB
			8'd14 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 56 -> 1
			// srcs: (27, 7)(678) -1 --> (678) -1:PUNB, pass, PENB
			8'd15 : rdata = 43'b1100011011111111000000000000000000100000000;
			// PEs: 56 -> 1
			// srcs: (28, 8)(486) 6 --> (486) 6:PUNB, pass, PENB
			8'd16 : rdata = 43'b1100011011111111000000000000000000100000000;
			// PEs: 56 -> 1
			// srcs: (29, 9)(489) -6 --> (489) -6:PUNB, pass, PENB
			8'd17 : rdata = 43'b1100011011111111000000000000000000100000000;
			// PEs: 8 -> 1
			// srcs: (30, 12)(695) 0 --> (695) 0:PUGB1, pass, PENB
			8'd18 : rdata = 43'b1100011100000011000000000000000000100000000;
			// PEs: 16 -> 1
			// srcs: (31, 17)(561) 2 --> (561) 2:PUGB2, pass, PENB
			8'd19 : rdata = 43'b1100011100000101000000000000000000100000000;
			// PEs: 1 -> 48
			// srcs: (33, 21)(633) 1 --> (633) 1:PEGB1, pass, PUGB6
			8'd20 : rdata = 43'b1100011100000010000000000000000000000001110;
			// PEs: 1 -> 8
			// srcs: (36, 25)(685) -4 --> (685) -4:PEGB1, pass, PUNB
			8'd21 : rdata = 43'b1100011100000010000000000000000001000000000;
			// PEs: 1 -> 16
			// srcs: (37, 26)(696) 9 --> (696) 9:PEGB1, pass, PUGB2
			8'd22 : rdata = 43'b1100011100000010000000000000000000000001010;
			// PEs: 2 -> 8
			// srcs: (44, 30)(683) -3 --> (683) -3:PEGB2, pass, PUNB
			8'd23 : rdata = 43'b1100011100000100000000000000000001000000000;
			// PEs: 16 -> 1
			// srcs: (47, 19)(567) 0 --> (567) 0:PUGB2, pass, PENB
			8'd24 : rdata = 43'b1100011100000101000000000000000000100000000;
			// PEs: 16 -> 0
			// srcs: (48, 22)(642) 12 --> (642) 12:PUGB2, pass, NI0
			8'd25 : rdata = 43'b1100011100000101000000000001000000000000000;
			// PEs: 48 -> 1
			// srcs: (49, 23)(644) 10 --> (644) 10:PUGB6, pass, PENB
			8'd26 : rdata = 43'b1100011100001101000000000000000000100000000;
			// PEs: 0 -> 1
			// srcs: (55, 24)(642) 12 --> (642) 12:NI0, pass, PENB
			8'd27 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 56 -> 1
			// srcs: (56, 27)(755) 16 --> (755) 16:PUNB, pass, PENB
			8'd28 : rdata = 43'b1100011011111111000000000000000000100000000;
			// PEs: 1 -> 48
			// srcs: (62, 29)(645) 22 --> (645) 22:PEGB1, pass, PUGB6
			8'd29 : rdata = 43'b1100011100000010000000000000000000000001110;
			// PEs: 56 -> 1
			// srcs: (65, 28)(760) -2 --> (760) -2:PUNB, pass, PENB
			8'd30 : rdata = 43'b1100011011111111000000000000000000100000000;
			// PEs: 32 -> 1
			// srcs: (106, 31)(775) 7 --> (775) 7:PUGB4, pass, PENB
			8'd31 : rdata = 43'b1100011100001001000000000000000000100000000;
			// PEs: 1 -> 48
			// srcs: (114, 32)(776) 21 --> (776) 21:PEGB1, pass, PUGB6
			8'd32 : rdata = 43'b1100011100000010000000000000000000000001110;
			// PEs: 24 -> 0
			// srcs: (146, 33)(703) 35 --> (703) 35:PUGB3, pass, NI0
			8'd33 : rdata = 43'b1100011100000111000000000001000000000000000;
			// PEs: 48 -> 1
			// srcs: (151, 34)(802) 57 --> (802) 57:PUGB6, pass, PENB
			8'd34 : rdata = 43'b1100011100001101000000000000000000100000000;
			// PEs: 0 -> 1
			// srcs: (158, 35)(703) 35 --> (703) 35:NI0, pass, PENB
			8'd35 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 1 -> 32
			// srcs: (165, 36)(803) 92 --> (803) 92:PEGB1, pass, PUGB4
			8'd36 : rdata = 43'b1100011100000010000000000000000000000001100;
			// PEs: 32 -> 1
			// srcs: (196, 37)(809) 0 --> (809) 0:PUGB4, pass, PENB
			8'd37 : rdata = 43'b1100011100001001000000000000000000100000000;
			// PEs: 32 -> 2
			// srcs: (200, 38)(809) 0 --> (809) 0:PUGB4, pass, PEGB2
			8'd38 : rdata = 43'b1100011100001001000000000000000000010100000;
			// PEs: 32 -> 3
			// srcs: (201, 39)(809) 0 --> (809) 0:PUGB4, pass, PEGB3
			8'd39 : rdata = 43'b1100011100001001000000000000000000010110000;
			// PEs: 32 -> 4
			// srcs: (202, 40)(809) 0 --> (809) 0:PUGB4, pass, PEGB4
			8'd40 : rdata = 43'b1100011100001001000000000000000000011000000;
			// PEs: 32 -> 5
			// srcs: (203, 41)(809) 0 --> (809) 0:PUGB4, pass, PEGB5
			8'd41 : rdata = 43'b1100011100001001000000000000000000011010000;
			// PEs: 32 -> 6
			// srcs: (204, 42)(809) 0 --> (809) 0:PUGB4, pass, PEGB6
			8'd42 : rdata = 43'b1100011100001001000000000000000000011100000;
			// PEs: 32 -> 7
			// srcs: (206, 43)(809) 0 --> (809) 0:PUGB4, pass, PEGB7
			8'd43 : rdata = 43'b1100011100001001000000000000000000011110000;
			// PEs: 32 -> 1
			// srcs: (275, 44)(809) 0 --> (809) 0:PUGB4, pass, PENB
			8'd44 : rdata = 43'b1100011100001001000000000000000000100000000;
			// PEs: 32 -> 2
			// srcs: (276, 45)(809) 0 --> (809) 0:PUGB4, pass, PEGB2
			8'd45 : rdata = 43'b1100011100001001000000000000000000010100000;
			// PEs: 32 -> 3
			// srcs: (277, 46)(809) 0 --> (809) 0:PUGB4, pass, PEGB3
			8'd46 : rdata = 43'b1100011100001001000000000000000000010110000;
			// PEs: 32 -> 4
			// srcs: (278, 47)(809) 0 --> (809) 0:PUGB4, pass, PEGB4
			8'd47 : rdata = 43'b1100011100001001000000000000000000011000000;
			// PEs: 32 -> 5
			// srcs: (280, 48)(809) 0 --> (809) 0:PUGB4, pass, PEGB5
			8'd48 : rdata = 43'b1100011100001001000000000000000000011010000;
			// PEs: 32 -> 6
			// srcs: (281, 49)(809) 0 --> (809) 0:PUGB4, pass, PEGB6
			8'd49 : rdata = 43'b1100011100001001000000000000000000011100000;
			// PEs: 32 -> 7
			// srcs: (283, 50)(809) 0 --> (809) 0:PUGB4, pass, PEGB7
			8'd50 : rdata = 43'b1100011100001001000000000000000000011110000;
			// PEs: 32 -> 1
			// srcs: (288, 51)(809) 0 --> (809) 0:PUGB4, pass, PENB
			8'd51 : rdata = 43'b1100011100001001000000000000000000100000000;
			// PEs: 32 -> 2
			// srcs: (291, 52)(809) 0 --> (809) 0:PUGB4, pass, PEGB2
			8'd52 : rdata = 43'b1100011100001001000000000000000000010100000;
			// PEs: 32 -> 3
			// srcs: (294, 53)(809) 0 --> (809) 0:PUGB4, pass, PEGB3
			8'd53 : rdata = 43'b1100011100001001000000000000000000010110000;
			// PEs: 32 -> 4
			// srcs: (297, 54)(809) 0 --> (809) 0:PUGB4, pass, PEGB4
			8'd54 : rdata = 43'b1100011100001001000000000000000000011000000;
			// PEs: 32 -> 5
			// srcs: (304, 55)(809) 0 --> (809) 0:PUGB4, pass, PEGB5
			8'd55 : rdata = 43'b1100011100001001000000000000000000011010000;
			// PEs: 32 -> 6
			// srcs: (307, 56)(809) 0 --> (809) 0:PUGB4, pass, PEGB6
			8'd56 : rdata = 43'b1100011100001001000000000000000000011100000;
			// PEs: 32 -> 7
			// srcs: (310, 57)(809) 0 --> (809) 0:PUGB4, pass, PEGB7
			8'd57 : rdata = 43'b1100011100001001000000000000000000011110000;
			// PEs: 32 -> 1
			// srcs: (352, 58)(809) 0 --> (809) 0:PUGB4, pass, PENB
			8'd58 : rdata = 43'b1100011100001001000000000000000000100000000;
			// PEs: 32 -> 2
			// srcs: (353, 59)(809) 0 --> (809) 0:PUGB4, pass, PEGB2
			8'd59 : rdata = 43'b1100011100001001000000000000000000010100000;
			// PEs: 32 -> 3
			// srcs: (355, 60)(809) 0 --> (809) 0:PUGB4, pass, PEGB3
			8'd60 : rdata = 43'b1100011100001001000000000000000000010110000;
			// PEs: 32 -> 4
			// srcs: (356, 61)(809) 0 --> (809) 0:PUGB4, pass, PEGB4
			8'd61 : rdata = 43'b1100011100001001000000000000000000011000000;
			// PEs: 32 -> 5
			// srcs: (358, 62)(809) 0 --> (809) 0:PUGB4, pass, PEGB5
			8'd62 : rdata = 43'b1100011100001001000000000000000000011010000;
			// PEs: 32 -> 6
			// srcs: (359, 63)(809) 0 --> (809) 0:PUGB4, pass, PEGB6
			8'd63 : rdata = 43'b1100011100001001000000000000000000011100000;
			// PEs: 32 -> 7
			// srcs: (361, 64)(809) 0 --> (809) 0:PUGB4, pass, PEGB7
			8'd64 : rdata = 43'b1100011100001001000000000000000000011110000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 1) begin
	always @(*) begin
		case(address)
			// PEs: 1, 1 -> 3
			// srcs: (1, 0)(4) 0, (205) 1 --> (405) 0:ND0, NW0, *, PEGB3
			8'd0 : rdata = 43'b0001101100000000010000000000000000010110000;
			// PEs: 1, 1 -> 2
			// srcs: (2, 1)(81) 0, (282) 0 --> (482) 0:ND1, NW1, *, PENB
			8'd1 : rdata = 43'b0001101100000001010000000010000000100000000;
			// PEs: 1, 1 -> 2
			// srcs: (3, 2)(158) -1, (359) -3 --> (559) 3:ND2, NW2, *, PENB
			8'd2 : rdata = 43'b0001101100000010010000000100000000100000000;
			// PEs: 1, 1 -> 0
			// srcs: (4, 3)(94) -1, (295) 1 --> (495) -1:ND3, NW3, *, PEGB0
			8'd3 : rdata = 43'b0001101100000011010000000110000000010000000;
			// PEs: 6 -> 
			// srcs: (6, 4)(410) -6 --> (410) -6:PEGB6, pass, 
			8'd4 : rdata = 43'b1100011100001100000000000000000000000000000;
			// PEs: 5, 1 -> 0
			// srcs: (9, 5)(409) 2, (410) -6 --> (608) -4:PEGB5, ALU, +, PEGB0
			8'd5 : rdata = 43'b0000111100001010001111111110000000010000000;
			// PEs: 0 -> 
			// srcs: (21, 6)(632) 2 --> (632) 2:PENB, pass, 
			8'd6 : rdata = 43'b1100011011111110000000000000000000000000000;
			// PEs: 1, 0 -> 0
			// srcs: (28, 7)(632) 2, (436) -1 --> (633) 1:ALU, PENB, +, PEGB0
			8'd7 : rdata = 43'b0000100111111111110111111100000000010000000;
			// PEs: 0, 2 -> 1
			// srcs: (29, 8)(678) -1, (679) -2 --> (680) -3:PENB, PEGB2, +, NI0
			8'd8 : rdata = 43'b0000111011111110111000001001000000000000000;
			// PEs: 4, 0 -> 2
			// srcs: (30, 9)(681) -6, (486) 6 --> (682) 0:PEGB4, PENB, +, PENB
			8'd9 : rdata = 43'b0000111100001000110111111100000000100000000;
			// PEs: 6, 0 -> 0
			// srcs: (31, 10)(684) 2, (489) -6 --> (685) -4:PEGB6, PENB, +, PEGB0
			8'd10 : rdata = 43'b0000111100001100110111111100000000010000000;
			// PEs: 0, 3 -> 0
			// srcs: (32, 11)(695) 0, (501) 9 --> (696) 9:PENB, PEGB3, +, PEGB0
			8'd11 : rdata = 43'b0000111011111110111000001100000000010000000;
			// PEs: 2, 0 -> 1
			// srcs: (33, 12)(756) 5, (561) 2 --> (757) 7:PEGB2, PENB, +, NI1
			8'd12 : rdata = 43'b0000111100000100110111111101010000000000000;
			// PEs: 1 -> 2
			// srcs: (37, 16)(680) -3 --> (680) -3:NI0, pass, PENB
			8'd13 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 6, 0 -> 1
			// srcs: (49, 13)(761) -7, (567) 0 --> (762) -7:PEGB6, PENB, +, NI0
			8'd14 : rdata = 43'b0000111100001100110111111101000000000000000;
			// PEs: 0 -> 
			// srcs: (51, 14)(644) 10 --> (644) 10:PENB, pass, 
			8'd15 : rdata = 43'b1100011011111110000000000000000000000000000;
			// PEs: 0, 1 -> 0
			// srcs: (57, 15)(642) 12, (644) 10 --> (645) 22:PENB, ALU, +, PEGB0
			8'd16 : rdata = 43'b0000111011111110001111111110000000010000000;
			// PEs: 0, 1 -> 1
			// srcs: (58, 17)(755) 16, (757) 7 --> (758) 23:PENB, NI1, +, NI2
			8'd17 : rdata = 43'b0000111011111110101000000011100000000000000;
			// PEs: 0, 1 -> 2
			// srcs: (68, 18)(760) -2, (762) -7 --> (763) -9:PENB, NI0, +, PENB
			8'd18 : rdata = 43'b0000111011111110101000000000000000100000000;
			// PEs: 1 -> 2
			// srcs: (75, 19)(758) 23 --> (758) 23:NI2, pass, PENB
			8'd19 : rdata = 43'b1100010100000010000000000000000000100000000;
			// PEs: 2, 0 -> 0
			// srcs: (109, 20)(764) 14, (775) 7 --> (776) 21:PEGB2, PENB, +, PEGB0
			8'd20 : rdata = 43'b0000111100000100110111111100000000010000000;
			// PEs: 0 -> 
			// srcs: (153, 21)(802) 57 --> (802) 57:PENB, pass, 
			8'd21 : rdata = 43'b1100011011111110000000000000000000000000000;
			// PEs: 0, 1 -> 0
			// srcs: (160, 22)(703) 35, (802) 57 --> (803) 92:PENB, ALU, +, PEGB0
			8'd22 : rdata = 43'b0000111011111110001111111110000000010000000;
			// PEs: 0, 1 -> 2
			// srcs: (199, 23)(809) 0, (4) 0 --> (810) 0:PENB, ND0, *, PENB
			8'd23 : rdata = 43'b0001111011111110011000000000000000100000000;
			// PEs: 1, 2 -> 1
			// srcs: (208, 27)(205) 1, (1010) 0 --> (1210) 1:NW0, PEGB2, -, NW0
			8'd24 : rdata = 43'b0001001000000000111000001000001000000000000;
			// PEs: 0, 1 -> 2
			// srcs: (277, 24)(809) 0, (81) 0 --> (887) 0:PENB, ND1, *, PENB
			8'd25 : rdata = 43'b0001111011111110011000000010000000100000000;
			// PEs: 1, 2 -> 1
			// srcs: (286, 28)(282) 0, (1087) 0 --> (1287) 0:NW1, PEGB2, -, NW1
			8'd26 : rdata = 43'b0001001000000001111000001000001010000000000;
			// PEs: 0, 1 -> 2
			// srcs: (290, 25)(809) 0, (94) -1 --> (900) 0:PENB, ND3, *, PENB
			8'd27 : rdata = 43'b0001111011111110011000000110000000100000000;
			// PEs: 1, 2 -> 1
			// srcs: (299, 29)(295) 1, (1100) 0 --> (1300) 1:NW3, PEGB2, -, NW3
			8'd28 : rdata = 43'b0001001000000011111000001000001110000000000;
			// PEs: 0, 1 -> 2
			// srcs: (354, 26)(809) 0, (158) -1 --> (964) 0:PENB, ND2, *, PENB
			8'd29 : rdata = 43'b0001111011111110011000000100000000100000000;
			// PEs: 1, 2 -> 1
			// srcs: (363, 30)(359) -3, (1164) 0 --> (1364) -3:NW2, PEGB2, -, NW2
			8'd30 : rdata = 43'b0001001000000010111000001000001100000000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 2) begin
	always @(*) begin
		case(address)
			// PEs: 2, 2 -> 3
			// srcs: (1, 0)(5) -3, (206) -1 --> (406) 3:ND0, NW0, *, PENB
			8'd0 : rdata = 43'b0001101100000000010000000000000000100000000;
			// PEs: 2, 2 -> 2
			// srcs: (2, 1)(82) -2, (283) 1 --> (483) -2:ND1, NW1, *, NI0
			8'd1 : rdata = 43'b0001101100000001010000000011000000000000000;
			// PEs: 2, 2 -> 2
			// srcs: (3, 2)(159) -2, (360) -1 --> (560) 2:ND2, NW2, *, NI1
			8'd2 : rdata = 43'b0001101100000010010000000101010000000000000;
			// PEs: 2, 2 -> 0
			// srcs: (4, 3)(97) -2, (298) -2 --> (498) 4:ND3, NW3, *, PEGB0
			8'd3 : rdata = 43'b0001101100000011010000000110000000010000000;
			// PEs: 1, 2 -> 1
			// srcs: (5, 5)(482) 0, (483) -2 --> (679) -2:PENB, NI0, +, PEGB1
			8'd4 : rdata = 43'b0000111011111110101000000000000000010010000;
			// PEs: 1, 2 -> 1
			// srcs: (6, 4)(559) 3, (560) 2 --> (756) 5:PENB, NI1, +, PEGB1
			8'd5 : rdata = 43'b0000111011111110101000000010000000010010000;
			// PEs: 1 -> 
			// srcs: (32, 6)(682) 0 --> (682) 0:PENB, pass, 
			8'd6 : rdata = 43'b1100011011111110000000000000000000000000000;
			// PEs: 1, 2 -> 0
			// srcs: (39, 7)(680) -3, (682) 0 --> (683) -3:PENB, ALU, +, PEGB0
			8'd7 : rdata = 43'b0000111011111110001111111110000000010000000;
			// PEs: 1 -> 
			// srcs: (70, 8)(763) -9 --> (763) -9:PENB, pass, 
			8'd8 : rdata = 43'b1100011011111110000000000000000000000000000;
			// PEs: 1, 2 -> 1
			// srcs: (77, 9)(758) 23, (763) -9 --> (764) 14:PENB, ALU, +, PEGB1
			8'd9 : rdata = 43'b0000111011111110001111111110000000010010000;
			// PEs: 2, 1 -> 1
			// srcs: (202, 14)(3) 1, (810) 0 --> (1010) 0:NM0, PENB, *, PEGB1
			8'd10 : rdata = 43'b0001110000000000110111111100000000010010000;
			// PEs: 0, 2 -> 3
			// srcs: (205, 10)(809) 0, (5) -3 --> (811) 0:PEGB0, ND0, *, PENB
			8'd11 : rdata = 43'b0001111100000000011000000000000000100000000;
			// PEs: 2, 3 -> 2
			// srcs: (214, 19)(206) -1, (1011) 0 --> (1211) -1:NW0, PEGB3, -, NW0
			8'd12 : rdata = 43'b0001001000000000111000001100001000000000000;
			// PEs: 2, 1 -> 1
			// srcs: (280, 15)(3) 1, (887) 0 --> (1087) 0:NM0, PENB, *, PEGB1
			8'd13 : rdata = 43'b0001110000000000110111111100000000010010000;
			// PEs: 0, 2 -> 3
			// srcs: (281, 11)(809) 0, (82) -2 --> (888) 0:PEGB0, ND1, *, PENB
			8'd14 : rdata = 43'b0001111100000000011000000010000000100000000;
			// PEs: 2, 3 -> 2
			// srcs: (290, 20)(283) 1, (1088) 0 --> (1288) 1:NW1, PEGB3, -, NW1
			8'd15 : rdata = 43'b0001001000000001111000001100001010000000000;
			// PEs: 2, 1 -> 1
			// srcs: (293, 16)(3) 1, (900) 0 --> (1100) 0:NM0, PENB, *, PEGB1
			8'd16 : rdata = 43'b0001110000000000110111111100000000010010000;
			// PEs: 0, 2 -> 
			// srcs: (296, 12)(809) 0, (97) -2 --> (903) 0:PEGB0, ND3, *, 
			8'd17 : rdata = 43'b0001111100000000011000000110000000000000000;
			// PEs: 2, 2 -> 
			// srcs: (299, 17)(3) 1, (903) 0 --> (1103) 0:NM0, ALU, *, 
			8'd18 : rdata = 43'b0001110000000000001111111110000000000000000;
			// PEs: 2, 2 -> 2
			// srcs: (302, 21)(298) -2, (1103) 0 --> (1303) -2:NW3, ALU, -, NW3
			8'd19 : rdata = 43'b0001001000000011001111111110001110000000000;
			// PEs: 2, 1 -> 1
			// srcs: (357, 18)(3) 1, (964) 0 --> (1164) 0:NM0, PENB, *, PEGB1
			8'd20 : rdata = 43'b0001110000000000110111111100000000010010000;
			// PEs: 0, 2 -> 3
			// srcs: (358, 13)(809) 0, (159) -2 --> (965) 0:PEGB0, ND2, *, PENB
			8'd21 : rdata = 43'b0001111100000000011000000100000000100000000;
			// PEs: 2, 3 -> 2
			// srcs: (367, 22)(360) -1, (1165) 0 --> (1365) -1:NW2, PEGB3, -, NW2
			8'd22 : rdata = 43'b0001001000000010111000001100001100000000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 3) begin
	always @(*) begin
		case(address)
			// PEs: 3, 3 -> 5
			// srcs: (1, 0)(6) -1, (207) 2 --> (407) -2:ND0, NW0, *, PEGB5
			8'd0 : rdata = 43'b0001101100000000010000000000000000011010000;
			// PEs: 3, 3 -> 4
			// srcs: (2, 1)(83) -2, (284) 2 --> (484) -4:ND1, NW1, *, PENB
			8'd1 : rdata = 43'b0001101100000001010000000010000000100000000;
			// PEs: 3, 3 -> 4
			// srcs: (3, 2)(161) 2, (362) 2 --> (562) 4:ND2, NW2, *, PENB
			8'd2 : rdata = 43'b0001101100000010010000000100000000100000000;
			// PEs: 3, 3 -> 1
			// srcs: (4, 3)(100) -3, (301) -3 --> (501) 9:ND3, NW3, *, PEGB1
			8'd3 : rdata = 43'b0001101100000011010000000110000000010010000;
			// PEs: 1, 2 -> 7
			// srcs: (7, 4)(405) 0, (406) 3 --> (605) 3:PEGB1, PENB, +, PEGB7
			8'd4 : rdata = 43'b0000111100000010110111111100000000011110000;
			// PEs: 0, 3 -> 3
			// srcs: (206, 5)(809) 0, (6) -1 --> (812) 0:PEGB0, ND0, *, NI0
			8'd5 : rdata = 43'b0001111100000000011000000001000000000000000;
			// PEs: 3, 2 -> 2
			// srcs: (208, 9)(3) 1, (811) 0 --> (1011) 0:NM0, PENB, *, PEGB2
			8'd6 : rdata = 43'b0001110000000000110111111100000000010100000;
			// PEs: 3, 3 -> 
			// srcs: (209, 10)(3) 1, (812) 0 --> (1012) 0:NM0, NI0, *, 
			8'd7 : rdata = 43'b0001110000000000101000000000000000000000000;
			// PEs: 3, 3 -> 3
			// srcs: (212, 14)(207) 2, (1012) 0 --> (1212) 2:NW0, ALU, -, NW0
			8'd8 : rdata = 43'b0001001000000000001111111110001000000000000;
			// PEs: 0, 3 -> 4
			// srcs: (282, 6)(809) 0, (83) -2 --> (889) 0:PEGB0, ND1, *, PENB
			8'd9 : rdata = 43'b0001111100000000011000000010000000100000000;
			// PEs: 3, 2 -> 2
			// srcs: (284, 11)(3) 1, (888) 0 --> (1088) 0:NM0, PENB, *, PEGB2
			8'd10 : rdata = 43'b0001110000000000110111111100000000010100000;
			// PEs: 3, 4 -> 3
			// srcs: (291, 15)(284) 2, (1089) 0 --> (1289) 2:NW1, PEGB4, -, NW1
			8'd11 : rdata = 43'b0001001000000001111000010000001010000000000;
			// PEs: 0, 3 -> 
			// srcs: (299, 7)(809) 0, (100) -3 --> (906) 0:PEGB0, ND3, *, 
			8'd12 : rdata = 43'b0001111100000000011000000110000000000000000;
			// PEs: 3, 3 -> 
			// srcs: (302, 12)(3) 1, (906) 0 --> (1106) 0:NM0, ALU, *, 
			8'd13 : rdata = 43'b0001110000000000001111111110000000000000000;
			// PEs: 3, 3 -> 3
			// srcs: (305, 16)(301) -3, (1106) 0 --> (1306) -3:NW3, ALU, -, NW3
			8'd14 : rdata = 43'b0001001000000011001111111110001110000000000;
			// PEs: 0, 3 -> 4
			// srcs: (360, 8)(809) 0, (161) 2 --> (967) 0:PEGB0, ND2, *, PENB
			8'd15 : rdata = 43'b0001111100000000011000000100000000100000000;
			// PEs: 3, 2 -> 2
			// srcs: (361, 13)(3) 1, (965) 0 --> (1165) 0:NM0, PENB, *, PEGB2
			8'd16 : rdata = 43'b0001110000000000110111111100000000010100000;
			// PEs: 3, 4 -> 3
			// srcs: (369, 17)(362) 2, (1167) 0 --> (1367) 2:NW2, PEGB4, -, NW2
			8'd17 : rdata = 43'b0001001000000010111000010000001100000000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 4) begin
	always @(*) begin
		case(address)
			// PEs: 4, 4 -> 5
			// srcs: (1, 0)(7) -3, (208) 1 --> (408) -3:ND0, NW0, *, PENB
			8'd0 : rdata = 43'b0001101100000000010000000000000000100000000;
			// PEs: 4, 4 -> 4
			// srcs: (2, 1)(84) 2, (285) -1 --> (485) -2:ND1, NW1, *, NI0
			8'd1 : rdata = 43'b0001101100000001010000000011000000000000000;
			// PEs: 4, 4 -> 4
			// srcs: (3, 2)(162) -1, (363) 2 --> (563) -2:ND2, NW2, *, NI1
			8'd2 : rdata = 43'b0001101100000010010000000101010000000000000;
			// PEs: 4, 4 -> 0
			// srcs: (4, 3)(103) -2, (304) -1 --> (504) 2:ND3, NW3, *, PEGB0
			8'd3 : rdata = 43'b0001101100000011010000000110000000010000000;
			// PEs: 3, 4 -> 1
			// srcs: (5, 4)(484) -4, (485) -2 --> (681) -6:PENB, NI0, +, PEGB1
			8'd4 : rdata = 43'b0000111011111110101000000000000000010010000;
			// PEs: 3, 4 -> 0
			// srcs: (6, 5)(562) 4, (563) -2 --> (759) 2:PENB, NI1, +, PEGB0
			8'd5 : rdata = 43'b0000111011111110101000000010000000010000000;
			// PEs: 0, 4 -> 5
			// srcs: (207, 6)(809) 0, (7) -3 --> (813) 0:PEGB0, ND0, *, PENB
			8'd6 : rdata = 43'b0001111100000000011000000000000000100000000;
			// PEs: 4, 5 -> 4
			// srcs: (216, 14)(208) 1, (1013) 0 --> (1213) 1:NW0, PEGB5, -, NW0
			8'd7 : rdata = 43'b0001001000000000111000010100001000000000000;
			// PEs: 0, 4 -> 4
			// srcs: (283, 7)(809) 0, (84) 2 --> (890) 0:PEGB0, ND1, *, NI0
			8'd8 : rdata = 43'b0001111100000000011000000011000000000000000;
			// PEs: 4, 3 -> 3
			// srcs: (285, 10)(3) 1, (889) 0 --> (1089) 0:NM0, PENB, *, PEGB3
			8'd9 : rdata = 43'b0001110000000000110111111100000000010110000;
			// PEs: 4, 4 -> 
			// srcs: (286, 11)(3) 1, (890) 0 --> (1090) 0:NM0, NI0, *, 
			8'd10 : rdata = 43'b0001110000000000101000000000000000000000000;
			// PEs: 4, 4 -> 4
			// srcs: (289, 15)(285) -1, (1090) 0 --> (1290) -1:NW1, ALU, -, NW1
			8'd11 : rdata = 43'b0001001000000001001111111110001010000000000;
			// PEs: 0, 4 -> 
			// srcs: (302, 8)(809) 0, (103) -2 --> (909) 0:PEGB0, ND3, *, 
			8'd12 : rdata = 43'b0001111100000000011000000110000000000000000;
			// PEs: 4, 4 -> 
			// srcs: (305, 12)(3) 1, (909) 0 --> (1109) 0:NM0, ALU, *, 
			8'd13 : rdata = 43'b0001110000000000001111111110000000000000000;
			// PEs: 4, 4 -> 4
			// srcs: (308, 16)(304) -1, (1109) 0 --> (1309) -1:NW3, ALU, -, NW3
			8'd14 : rdata = 43'b0001001000000011001111111110001110000000000;
			// PEs: 0, 4 -> 5
			// srcs: (361, 9)(809) 0, (162) -1 --> (968) 0:PEGB0, ND2, *, PENB
			8'd15 : rdata = 43'b0001111100000000011000000100000000100000000;
			// PEs: 4, 3 -> 3
			// srcs: (363, 13)(3) 1, (967) 0 --> (1167) 0:NM0, PENB, *, PEGB3
			8'd16 : rdata = 43'b0001110000000000110111111100000000010110000;
			// PEs: 4, 5 -> 4
			// srcs: (370, 17)(363) 2, (1168) 0 --> (1368) 2:NW2, PEGB5, -, NW2
			8'd17 : rdata = 43'b0001001000000010111000010100001100000000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 5) begin
	always @(*) begin
		case(address)
			// PEs: 5, 5 -> 1
			// srcs: (1, 0)(8) -2, (209) -1 --> (409) 2:ND0, NW0, *, PEGB1
			8'd0 : rdata = 43'b0001101100000000010000000000000000010010000;
			// PEs: 5, 5 -> 6
			// srcs: (2, 1)(86) 2, (287) 1 --> (487) 2:ND1, NW1, *, PENB
			8'd1 : rdata = 43'b0001101100000001010000000010000000100000000;
			// PEs: 5, 5 -> 6
			// srcs: (3, 2)(164) -2, (365) 2 --> (565) -4:ND2, NW2, *, PENB
			8'd2 : rdata = 43'b0001101100000010010000000100000000100000000;
			// PEs: 5, 5 -> 0
			// srcs: (4, 3)(110) 2, (311) 2 --> (511) 4:ND3, NW3, *, PEGB0
			8'd3 : rdata = 43'b0001101100000011010000000110000000010000000;
			// PEs: 3, 4 -> 7
			// srcs: (7, 4)(407) -2, (408) -3 --> (606) -5:PEGB3, PENB, +, PEGB7
			8'd4 : rdata = 43'b0000111100000110110111111100000000011110000;
			// PEs: 0, 5 -> 5
			// srcs: (208, 5)(809) 0, (8) -2 --> (814) 0:PEGB0, ND0, *, NI0
			8'd5 : rdata = 43'b0001111100000000011000000001000000000000000;
			// PEs: 5, 4 -> 4
			// srcs: (210, 9)(3) 1, (813) 0 --> (1013) 0:NM0, PENB, *, PEGB4
			8'd6 : rdata = 43'b0001110000000000110111111100000000011000000;
			// PEs: 5, 5 -> 
			// srcs: (211, 10)(3) 1, (814) 0 --> (1014) 0:NM0, NI0, *, 
			8'd7 : rdata = 43'b0001110000000000101000000000000000000000000;
			// PEs: 5, 5 -> 5
			// srcs: (214, 14)(209) -1, (1014) 0 --> (1214) -1:NW0, ALU, -, NW0
			8'd8 : rdata = 43'b0001001000000000001111111110001000000000000;
			// PEs: 0, 5 -> 
			// srcs: (285, 6)(809) 0, (86) 2 --> (892) 0:PEGB0, ND1, *, 
			8'd9 : rdata = 43'b0001111100000000011000000010000000000000000;
			// PEs: 5, 5 -> 
			// srcs: (288, 11)(3) 1, (892) 0 --> (1092) 0:NM0, ALU, *, 
			8'd10 : rdata = 43'b0001110000000000001111111110000000000000000;
			// PEs: 5, 5 -> 5
			// srcs: (291, 15)(287) 1, (1092) 0 --> (1292) 1:NW1, ALU, -, NW1
			8'd11 : rdata = 43'b0001001000000001001111111110001010000000000;
			// PEs: 0, 5 -> 
			// srcs: (309, 7)(809) 0, (110) 2 --> (916) 0:PEGB0, ND3, *, 
			8'd12 : rdata = 43'b0001111100000000011000000110000000000000000;
			// PEs: 5, 5 -> 
			// srcs: (312, 12)(3) 1, (916) 0 --> (1116) 0:NM0, ALU, *, 
			8'd13 : rdata = 43'b0001110000000000001111111110000000000000000;
			// PEs: 5, 5 -> 5
			// srcs: (315, 16)(311) 2, (1116) 0 --> (1316) 2:NW3, ALU, -, NW3
			8'd14 : rdata = 43'b0001001000000011001111111110001110000000000;
			// PEs: 0, 5 -> 6
			// srcs: (363, 8)(809) 0, (164) -2 --> (970) 0:PEGB0, ND2, *, PENB
			8'd15 : rdata = 43'b0001111100000000011000000100000000100000000;
			// PEs: 5, 4 -> 4
			// srcs: (364, 13)(3) 1, (968) 0 --> (1168) 0:NM0, PENB, *, PEGB4
			8'd16 : rdata = 43'b0001110000000000110111111100000000011000000;
			// PEs: 5, 6 -> 5
			// srcs: (372, 17)(365) 2, (1170) 0 --> (1370) 2:NW2, PEGB6, -, NW2
			8'd17 : rdata = 43'b0001001000000010111000011000001100000000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 6) begin
	always @(*) begin
		case(address)
			// PEs: 6, 6 -> 1
			// srcs: (1, 0)(9) 2, (210) -3 --> (410) -6:ND0, NW0, *, PEGB1
			8'd0 : rdata = 43'b0001101100000000010000000000000000010010000;
			// PEs: 6, 6 -> 6
			// srcs: (2, 1)(87) 0, (288) -1 --> (488) 0:ND1, NW1, *, NI0
			8'd1 : rdata = 43'b0001101100000001010000000011000000000000000;
			// PEs: 6, 6 -> 6
			// srcs: (3, 2)(165) -3, (366) 1 --> (566) -3:ND2, NW2, *, NI1
			8'd2 : rdata = 43'b0001101100000010010000000101010000000000000;
			// PEs: 6, 6 -> 0
			// srcs: (4, 3)(113) -2, (314) 2 --> (514) -4:ND3, NW3, *, PEGB0
			8'd3 : rdata = 43'b0001101100000011010000000110000000010000000;
			// PEs: 5, 6 -> 1
			// srcs: (5, 4)(487) 2, (488) 0 --> (684) 2:PENB, NI0, +, PEGB1
			8'd4 : rdata = 43'b0000111011111110101000000000000000010010000;
			// PEs: 5, 6 -> 1
			// srcs: (6, 5)(565) -4, (566) -3 --> (761) -7:PENB, NI1, +, PEGB1
			8'd5 : rdata = 43'b0000111011111110101000000010000000010010000;
			// PEs: 0, 6 -> 
			// srcs: (209, 6)(809) 0, (9) 2 --> (815) 0:PEGB0, ND0, *, 
			8'd6 : rdata = 43'b0001111100000000011000000000000000000000000;
			// PEs: 6, 6 -> 
			// srcs: (212, 10)(3) 1, (815) 0 --> (1015) 0:NM0, ALU, *, 
			8'd7 : rdata = 43'b0001110000000000001111111110000000000000000;
			// PEs: 6, 6 -> 6
			// srcs: (215, 14)(210) -3, (1015) 0 --> (1215) -3:NW0, ALU, -, NW0
			8'd8 : rdata = 43'b0001001000000000001111111110001000000000000;
			// PEs: 0, 6 -> 
			// srcs: (286, 7)(809) 0, (87) 0 --> (893) 0:PEGB0, ND1, *, 
			8'd9 : rdata = 43'b0001111100000000011000000010000000000000000;
			// PEs: 6, 6 -> 
			// srcs: (289, 11)(3) 1, (893) 0 --> (1093) 0:NM0, ALU, *, 
			8'd10 : rdata = 43'b0001110000000000001111111110000000000000000;
			// PEs: 6, 6 -> 6
			// srcs: (292, 15)(288) -1, (1093) 0 --> (1293) -1:NW1, ALU, -, NW1
			8'd11 : rdata = 43'b0001001000000001001111111110001010000000000;
			// PEs: 0, 6 -> 
			// srcs: (312, 8)(809) 0, (113) -2 --> (919) 0:PEGB0, ND3, *, 
			8'd12 : rdata = 43'b0001111100000000011000000110000000000000000;
			// PEs: 6, 6 -> 
			// srcs: (315, 12)(3) 1, (919) 0 --> (1119) 0:NM0, ALU, *, 
			8'd13 : rdata = 43'b0001110000000000001111111110000000000000000;
			// PEs: 6, 6 -> 6
			// srcs: (318, 16)(314) 2, (1119) 0 --> (1319) 2:NW3, ALU, -, NW3
			8'd14 : rdata = 43'b0001001000000011001111111110001110000000000;
			// PEs: 0, 6 -> 7
			// srcs: (364, 9)(809) 0, (165) -3 --> (971) 0:PEGB0, ND2, *, PENB
			8'd15 : rdata = 43'b0001111100000000011000000100000000100000000;
			// PEs: 6, 5 -> 5
			// srcs: (366, 13)(3) 1, (970) 0 --> (1170) 0:NM0, PENB, *, PEGB5
			8'd16 : rdata = 43'b0001110000000000110111111100000000011010000;
			// PEs: 6, 7 -> 6
			// srcs: (373, 17)(366) 1, (1171) 0 --> (1371) 1:NW2, PEGB7, -, NW2
			8'd17 : rdata = 43'b0001001000000010111000011100001100000000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 7) begin
	always @(*) begin
		case(address)
			// PEs: 7, 7 -> 0
			// srcs: (1, 0)(11) -1, (212) -3 --> (412) 3:ND0, NW0, *, PENB
			8'd0 : rdata = 43'b0001101100000000010000000000000000100000000;
			// PEs: 7, 7 -> 0
			// srcs: (2, 1)(89) 2, (290) -2 --> (490) -4:ND1, NW1, *, PENB
			8'd1 : rdata = 43'b0001101100000001010000000010000000100000000;
			// PEs: 7, 7 -> 0
			// srcs: (3, 2)(167) -1, (368) 1 --> (568) -1:ND2, NW2, *, PENB
			8'd2 : rdata = 43'b0001101100000010010000000100000000100000000;
			// PEs: 7, 7 -> 0
			// srcs: (4, 3)(116) -2, (317) 0 --> (517) 0:ND3, NW3, *, PENB
			8'd3 : rdata = 43'b0001101100000011010000000110000000100000000;
			// PEs: 5 -> 
			// srcs: (12, 4)(606) -5 --> (606) -5:PEGB5, pass, 
			8'd4 : rdata = 43'b1100011100001010000000000000000000000000000;
			// PEs: 3, 7 -> 0
			// srcs: (15, 5)(605) 3, (606) -5 --> (607) -2:PEGB3, ALU, +, PENB
			8'd5 : rdata = 43'b0000111100000110001111111110000000100000000;
			// PEs: 0, 7 -> 
			// srcs: (211, 6)(809) 0, (11) -1 --> (817) 0:PEGB0, ND0, *, 
			8'd6 : rdata = 43'b0001111100000000011000000000000000000000000;
			// PEs: 7, 7 -> 
			// srcs: (214, 10)(3) 1, (817) 0 --> (1017) 0:NM0, ALU, *, 
			8'd7 : rdata = 43'b0001110000000000001111111110000000000000000;
			// PEs: 7, 7 -> 7
			// srcs: (217, 15)(212) -3, (1017) 0 --> (1217) -3:NW0, ALU, -, NW0
			8'd8 : rdata = 43'b0001001000000000001111111110001000000000000;
			// PEs: 0, 7 -> 
			// srcs: (288, 7)(809) 0, (89) 2 --> (895) 0:PEGB0, ND1, *, 
			8'd9 : rdata = 43'b0001111100000000011000000010000000000000000;
			// PEs: 7, 7 -> 
			// srcs: (291, 11)(3) 1, (895) 0 --> (1095) 0:NM0, ALU, *, 
			8'd10 : rdata = 43'b0001110000000000001111111110000000000000000;
			// PEs: 7, 7 -> 7
			// srcs: (294, 16)(290) -2, (1095) 0 --> (1295) -2:NW1, ALU, -, NW1
			8'd11 : rdata = 43'b0001001000000001001111111110001010000000000;
			// PEs: 0, 7 -> 
			// srcs: (315, 8)(809) 0, (116) -2 --> (922) 0:PEGB0, ND3, *, 
			8'd12 : rdata = 43'b0001111100000000011000000110000000000000000;
			// PEs: 7, 7 -> 
			// srcs: (318, 12)(3) 1, (922) 0 --> (1122) 0:NM0, ALU, *, 
			8'd13 : rdata = 43'b0001110000000000001111111110000000000000000;
			// PEs: 7, 7 -> 7
			// srcs: (321, 17)(317) 0, (1122) 0 --> (1322) 0:NW3, ALU, -, NW3
			8'd14 : rdata = 43'b0001001000000011001111111110001110000000000;
			// PEs: 0, 7 -> 7
			// srcs: (366, 9)(809) 0, (167) -1 --> (973) 0:PEGB0, ND2, *, NI0
			8'd15 : rdata = 43'b0001111100000000011000000101000000000000000;
			// PEs: 7, 6 -> 6
			// srcs: (367, 13)(3) 1, (971) 0 --> (1171) 0:NM0, PENB, *, PEGB6
			8'd16 : rdata = 43'b0001110000000000110111111100000000011100000;
			// PEs: 7, 7 -> 
			// srcs: (369, 14)(3) 1, (973) 0 --> (1173) 0:NM0, NI0, *, 
			8'd17 : rdata = 43'b0001110000000000101000000000000000000000000;
			// PEs: 7, 7 -> 7
			// srcs: (372, 18)(368) 1, (1173) 0 --> (1373) 1:NW2, ALU, -, NW2
			8'd18 : rdata = 43'b0001001000000010001111111110001100000000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 8) begin
	always @(*) begin
		case(address)
			// PEs: 0 -> 9
			// srcs: (5, 0)(412) 3 --> (412) 3:PUNB, pass, PENB
			8'd0 : rdata = 43'b1100011011111111000000000000000000100000000;
			// PEs: 0 -> 9
			// srcs: (6, 1)(490) -4 --> (490) -4:PUNB, pass, PENB
			8'd1 : rdata = 43'b1100011011111111000000000000000000100000000;
			// PEs: 0 -> 9
			// srcs: (7, 2)(568) -1 --> (568) -1:PUNB, pass, PENB
			8'd2 : rdata = 43'b1100011011111111000000000000000000100000000;
			// PEs: 15 -> 0
			// srcs: (8, 13)(695) 0 --> (695) 0:PENB, pass, PUGB0
			8'd3 : rdata = 43'b1100011011111110000000000000000000000001000;
			// PEs: 11 -> 24
			// srcs: (9, 16)(526) -2 --> (526) -2:PEGB3, pass, PUGB3
			8'd4 : rdata = 43'b1100011100000110000000000000000000000001011;
			// PEs: 10 -> 16
			// srcs: (12, 4)(613) 4 --> (613) 4:PEGB2, pass, PUNB
			8'd5 : rdata = 43'b1100011100000100000000000000000001000000000;
			// PEs: 9 -> 32
			// srcs: (13, 3)(611) -3 --> (611) -3:PEGB1, pass, PUGB4
			8'd6 : rdata = 43'b1100011100000010000000000000000000000001100;
			// PEs: 11 -> 32
			// srcs: (14, 5)(617) -1 --> (617) -1:PEGB3, pass, PUGB4
			8'd7 : rdata = 43'b1100011100000110000000000000000000000001100;
			// PEs: 12 -> 40
			// srcs: (15, 6)(619) -2 --> (619) -2:PEGB4, pass, PUGB5
			8'd8 : rdata = 43'b1100011100001000000000000000000000000001101;
			// PEs: 13 -> 40
			// srcs: (16, 18)(536) 0 --> (536) 0:PEGB5, pass, PUGB5
			8'd9 : rdata = 43'b1100011100001010000000000000000000000001101;
			// PEs: 15 -> 48
			// srcs: (17, 20)(542) 0 --> (542) 0:PENB, pass, PUGB6
			8'd10 : rdata = 43'b1100011011111110000000000000000000000001110;
			// PEs: 9 -> 24
			// srcs: (18, 21)(765) -1 --> (765) -1:PEGB1, pass, PUGB3
			8'd11 : rdata = 43'b1100011100000010000000000000000000000001011;
			// PEs: 14 -> 24
			// srcs: (19, 22)(767) 6 --> (767) 6:PEGB6, pass, PUGB3
			8'd12 : rdata = 43'b1100011100001100000000000000000000000001011;
			// PEs: 24 -> 8
			// srcs: (20, 7)(635) 4 --> (635) 4:PUGB3, pass, NI0
			8'd13 : rdata = 43'b1100011100000111000000000001000000000000000;
			// PEs: 40 -> 9
			// srcs: (21, 8)(439) 0 --> (439) 0:PUGB5, pass, PENB
			8'd14 : rdata = 43'b1100011100001011000000000000000000100000000;
			// PEs: 9 -> 16
			// srcs: (23, 14)(520) 3 --> (520) 3:PEGB1, pass, PUNB
			8'd15 : rdata = 43'b1100011100000010000000000000000001000000000;
			// PEs: 10 -> 32
			// srcs: (24, 15)(523) 6 --> (523) 6:PEGB2, pass, PUGB4
			8'd16 : rdata = 43'b1100011100000100000000000000000000000001100;
			// PEs: 15 -> 24
			// srcs: (26, 24)(772) -2 --> (772) -2:PENB, pass, PUGB3
			8'd17 : rdata = 43'b1100011011111110000000000000000000000001011;
			// PEs: 8 -> 9
			// srcs: (27, 9)(635) 4 --> (635) 4:NI0, pass, PENB
			8'd18 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 56 -> 9
			// srcs: (28, 10)(492) 2 --> (492) 2:PUGB7, pass, PENB
			8'd19 : rdata = 43'b1100011100001111000000000000000000100000000;
			// PEs: 0 -> 9
			// srcs: (29, 11)(495) -1 --> (495) -1:PUNB, pass, PENB
			8'd20 : rdata = 43'b1100011011111111000000000000000000100000000;
			// PEs: 0 -> 9
			// srcs: (30, 12)(498) 4 --> (498) 4:PUNB, pass, PENB
			8'd21 : rdata = 43'b1100011011111111000000000000000000100000000;
			// PEs: 40 -> 9
			// srcs: (31, 19)(734) -2 --> (734) -2:PUGB5, pass, PENB
			8'd22 : rdata = 43'b1100011100001011000000000000000000100000000;
			// PEs: 12 -> 32
			// srcs: (32, 17)(529) -6 --> (529) -6:PEGB4, pass, PUGB4
			8'd23 : rdata = 43'b1100011100001000000000000000000000000001100;
			// PEs: 13 -> 32
			// srcs: (33, 23)(770) 0 --> (770) 0:PEGB5, pass, PUGB4
			8'd24 : rdata = 43'b1100011100001010000000000000000000000001100;
			// PEs: 9 -> 16
			// srcs: (38, 27)(735) 2 --> (735) 2:PEGB1, pass, PUNB
			8'd25 : rdata = 43'b1100011100000010000000000000000001000000000;
			// PEs: 10 -> 16
			// srcs: (46, 30)(694) 0 --> (694) 0:PEGB2, pass, PUNB
			8'd26 : rdata = 43'b1100011100000100000000000000000001000000000;
			// PEs: 32 -> 9
			// srcs: (47, 25)(638) 9 --> (638) 9:PUGB4, pass, PENB
			8'd27 : rdata = 43'b1100011100001001000000000000000000100000000;
			// PEs: 0 -> 9
			// srcs: (48, 26)(685) -4 --> (685) -4:PUNB, pass, PENB
			8'd28 : rdata = 43'b1100011011111111000000000000000000100000000;
			// PEs: 48 -> 9
			// srcs: (69, 28)(634) -2 --> (634) -2:PUGB6, pass, PENB
			8'd29 : rdata = 43'b1100011100001101000000000000000000100000000;
			// PEs: 0 -> 9
			// srcs: (70, 29)(683) -3 --> (683) -3:PUNB, pass, PENB
			8'd30 : rdata = 43'b1100011011111111000000000000000000100000000;
			// PEs: 40 -> 8
			// srcs: (77, 31)(616) -5 --> (616) -5:PUGB5, pass, NI0
			8'd31 : rdata = 43'b1100011100001011000000000001000000000000000;
			// PEs: 9 -> 16
			// srcs: (78, 34)(640) 11 --> (640) 11:PEGB1, pass, PUNB
			8'd32 : rdata = 43'b1100011100000010000000000000000001000000000;
			// PEs: 9 -> 16
			// srcs: (79, 35)(689) -12 --> (689) -12:PEGB1, pass, PUNB
			8'd33 : rdata = 43'b1100011100000010000000000000000001000000000;
			// PEs: 56 -> 9
			// srcs: (82, 32)(627) 5 --> (627) 5:PUGB7, pass, PENB
			8'd34 : rdata = 43'b1100011100001111000000000000000000100000000;
			// PEs: 8 -> 9
			// srcs: (89, 33)(616) -5 --> (616) -5:NI0, pass, PENB
			8'd35 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 9 -> 16
			// srcs: (96, 36)(628) 0 --> (628) 0:PEGB1, pass, PUNB
			8'd36 : rdata = 43'b1100011100000010000000000000000001000000000;
			// PEs: 32 -> 9
			// srcs: (207, 37)(809) 0 --> (809) 0:PUGB4, pass, PENB
			8'd37 : rdata = 43'b1100011100001001000000000000000000100000000;
			// PEs: 32 -> 10
			// srcs: (209, 38)(809) 0 --> (809) 0:PUGB4, pass, PEGB2
			8'd38 : rdata = 43'b1100011100001001000000000000000000010100000;
			// PEs: 32 -> 11
			// srcs: (210, 39)(809) 0 --> (809) 0:PUGB4, pass, PEGB3
			8'd39 : rdata = 43'b1100011100001001000000000000000000010110000;
			// PEs: 32 -> 12
			// srcs: (211, 40)(809) 0 --> (809) 0:PUGB4, pass, PEGB4
			8'd40 : rdata = 43'b1100011100001001000000000000000000011000000;
			// PEs: 32 -> 13
			// srcs: (212, 41)(809) 0 --> (809) 0:PUGB4, pass, PEGB5
			8'd41 : rdata = 43'b1100011100001001000000000000000000011010000;
			// PEs: 32 -> 14
			// srcs: (214, 42)(809) 0 --> (809) 0:PUGB4, pass, PEGB6
			8'd42 : rdata = 43'b1100011100001001000000000000000000011100000;
			// PEs: 32 -> 15
			// srcs: (215, 43)(809) 0 --> (809) 0:PUGB4, pass, PEGB7
			8'd43 : rdata = 43'b1100011100001001000000000000000000011110000;
			// PEs: 32 -> 9
			// srcs: (284, 44)(809) 0 --> (809) 0:PUGB4, pass, PENB
			8'd44 : rdata = 43'b1100011100001001000000000000000000100000000;
			// PEs: 32 -> 10
			// srcs: (286, 45)(809) 0 --> (809) 0:PUGB4, pass, PEGB2
			8'd45 : rdata = 43'b1100011100001001000000000000000000010100000;
			// PEs: 32 -> 11
			// srcs: (287, 46)(809) 0 --> (809) 0:PUGB4, pass, PEGB3
			8'd46 : rdata = 43'b1100011100001001000000000000000000010110000;
			// PEs: 32 -> 12
			// srcs: (289, 47)(809) 0 --> (809) 0:PUGB4, pass, PEGB4
			8'd47 : rdata = 43'b1100011100001001000000000000000000011000000;
			// PEs: 32 -> 13
			// srcs: (290, 48)(809) 0 --> (809) 0:PUGB4, pass, PEGB5
			8'd48 : rdata = 43'b1100011100001001000000000000000000011010000;
			// PEs: 32 -> 14
			// srcs: (292, 49)(809) 0 --> (809) 0:PUGB4, pass, PEGB6
			8'd49 : rdata = 43'b1100011100001001000000000000000000011100000;
			// PEs: 32 -> 15
			// srcs: (293, 50)(809) 0 --> (809) 0:PUGB4, pass, PEGB7
			8'd50 : rdata = 43'b1100011100001001000000000000000000011110000;
			// PEs: 32 -> 9
			// srcs: (313, 51)(809) 0 --> (809) 0:PUGB4, pass, PENB
			8'd51 : rdata = 43'b1100011100001001000000000000000000100000000;
			// PEs: 32 -> 10
			// srcs: (316, 52)(809) 0 --> (809) 0:PUGB4, pass, PEGB2
			8'd52 : rdata = 43'b1100011100001001000000000000000000010100000;
			// PEs: 32 -> 11
			// srcs: (319, 53)(809) 0 --> (809) 0:PUGB4, pass, PEGB3
			8'd53 : rdata = 43'b1100011100001001000000000000000000010110000;
			// PEs: 32 -> 12
			// srcs: (322, 54)(809) 0 --> (809) 0:PUGB4, pass, PEGB4
			8'd54 : rdata = 43'b1100011100001001000000000000000000011000000;
			// PEs: 32 -> 13
			// srcs: (329, 55)(809) 0 --> (809) 0:PUGB4, pass, PEGB5
			8'd55 : rdata = 43'b1100011100001001000000000000000000011010000;
			// PEs: 32 -> 14
			// srcs: (332, 56)(809) 0 --> (809) 0:PUGB4, pass, PEGB6
			8'd56 : rdata = 43'b1100011100001001000000000000000000011100000;
			// PEs: 32 -> 15
			// srcs: (335, 57)(809) 0 --> (809) 0:PUGB4, pass, PEGB7
			8'd57 : rdata = 43'b1100011100001001000000000000000000011110000;
			// PEs: 32 -> 9
			// srcs: (362, 58)(809) 0 --> (809) 0:PUGB4, pass, PENB
			8'd58 : rdata = 43'b1100011100001001000000000000000000100000000;
			// PEs: 32 -> 10
			// srcs: (364, 59)(809) 0 --> (809) 0:PUGB4, pass, PEGB2
			8'd59 : rdata = 43'b1100011100001001000000000000000000010100000;
			// PEs: 32 -> 11
			// srcs: (365, 60)(809) 0 --> (809) 0:PUGB4, pass, PEGB3
			8'd60 : rdata = 43'b1100011100001001000000000000000000010110000;
			// PEs: 32 -> 12
			// srcs: (367, 61)(809) 0 --> (809) 0:PUGB4, pass, PEGB4
			8'd61 : rdata = 43'b1100011100001001000000000000000000011000000;
			// PEs: 32 -> 13
			// srcs: (368, 62)(809) 0 --> (809) 0:PUGB4, pass, PEGB5
			8'd62 : rdata = 43'b1100011100001001000000000000000000011010000;
			// PEs: 32 -> 14
			// srcs: (370, 63)(809) 0 --> (809) 0:PUGB4, pass, PEGB6
			8'd63 : rdata = 43'b1100011100001001000000000000000000011100000;
			// PEs: 32 -> 15
			// srcs: (371, 64)(809) 0 --> (809) 0:PUGB4, pass, PEGB7
			8'd64 : rdata = 43'b1100011100001001000000000000000000011110000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 9) begin
	always @(*) begin
		case(address)
			// PEs: 9, 9 -> 9
			// srcs: (1, 0)(12) 2, (213) -3 --> (413) -6:ND0, NW0, *, NI0
			8'd0 : rdata = 43'b0001101100000000010000000001000000000000000;
			// PEs: 9, 9 -> 9
			// srcs: (2, 1)(90) -3, (291) 1 --> (491) -3:ND1, NW1, *, NI1
			8'd1 : rdata = 43'b0001101100000001010000000011010000000000000;
			// PEs: 9, 9 -> 9
			// srcs: (3, 2)(168) -1, (369) 0 --> (569) 0:ND2, NW2, *, NI2
			8'd2 : rdata = 43'b0001101100000010010000000101100000000000000;
			// PEs: 9, 9 -> 9
			// srcs: (4, 3)(119) -1, (320) -3 --> (520) 3:ND3, NW3, *, NI3
			8'd3 : rdata = 43'b0001101100000011010000000111110000000000000;
			// PEs: 8, 9 -> 8
			// srcs: (8, 4)(412) 3, (413) -6 --> (611) -3:PENB, NI0, +, PEGB0
			8'd4 : rdata = 43'b0000111011111110101000000000000000010000000;
			// PEs: 8, 9 -> 9
			// srcs: (9, 5)(490) -4, (491) -3 --> (686) -7:PENB, NI1, +, NI0
			8'd5 : rdata = 43'b0000111011111110101000000011000000000000000;
			// PEs: 8, 9 -> 8
			// srcs: (10, 6)(568) -1, (569) 0 --> (765) -1:PENB, NI2, +, PEGB0
			8'd6 : rdata = 43'b0000111011111110101000000100000000010000000;
			// PEs: 9 -> 8
			// srcs: (18, 12)(520) 3 --> (520) 3:NI3, pass, PEGB0
			8'd7 : rdata = 43'b1100010100000011000000000000000000010000000;
			// PEs: 8 -> 
			// srcs: (23, 7)(439) 0 --> (439) 0:PENB, pass, 
			8'd8 : rdata = 43'b1100011011111110000000000000000000000000000;
			// PEs: 8, 9 -> 9
			// srcs: (29, 8)(635) 4, (439) 0 --> (636) 4:PENB, ALU, +, NI1
			8'd9 : rdata = 43'b0000111011111110001111111111010000000000000;
			// PEs: 9, 8 -> 9
			// srcs: (30, 9)(686) -7, (492) 2 --> (687) -5:NI0, PENB, +, NI2
			8'd10 : rdata = 43'b0000110100000000110111111101100000000000000;
			// PEs: 11, 8 -> 9
			// srcs: (31, 10)(690) -8, (495) -1 --> (691) -9:PEGB3, PENB, +, NI0
			8'd11 : rdata = 43'b0000111100000110110111111101000000000000000;
			// PEs: 13, 8 -> 10
			// srcs: (32, 11)(692) 5, (498) 4 --> (693) 9:PEGB5, PENB, +, PENB
			8'd12 : rdata = 43'b0000111100001010110111111100000000100000000;
			// PEs: 8, 14 -> 8
			// srcs: (33, 13)(734) -2, (539) 4 --> (735) 2:PENB, PEGB6, +, PEGB0
			8'd13 : rdata = 43'b0000111011111110111000011000000000010000000;
			// PEs: 9 -> 10
			// srcs: (39, 16)(691) -9 --> (691) -9:NI0, pass, PENB
			8'd14 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 9, 8 -> 9
			// srcs: (49, 14)(636) 4, (638) 9 --> (639) 13:NI1, PENB, +, NI0
			8'd15 : rdata = 43'b0000110100000001110111111101000000000000000;
			// PEs: 8, 9 -> 9
			// srcs: (50, 15)(685) -4, (687) -5 --> (688) -9:PENB, NI2, +, NI1
			8'd16 : rdata = 43'b0000111011111110101000000101010000000000000;
			// PEs: 8, 9 -> 8
			// srcs: (72, 17)(634) -2, (639) 13 --> (640) 11:PENB, NI0, +, PEGB0
			8'd17 : rdata = 43'b0000111011111110101000000000000000010000000;
			// PEs: 8, 9 -> 8
			// srcs: (73, 18)(683) -3, (688) -9 --> (689) -12:PENB, NI1, +, PEGB0
			8'd18 : rdata = 43'b0000111011111110101000000010000000010000000;
			// PEs: 8 -> 
			// srcs: (84, 19)(627) 5 --> (627) 5:PENB, pass, 
			8'd19 : rdata = 43'b1100011011111110000000000000000000000000000;
			// PEs: 8, 9 -> 8
			// srcs: (91, 20)(616) -5, (627) 5 --> (628) 0:PENB, ALU, +, PEGB0
			8'd20 : rdata = 43'b0000111011111110001111111110000000010000000;
			// PEs: 8, 9 -> 10
			// srcs: (209, 21)(809) 0, (12) 2 --> (818) 0:PENB, ND0, *, PENB
			8'd21 : rdata = 43'b0001111011111110011000000000000000100000000;
			// PEs: 9, 10 -> 9
			// srcs: (218, 25)(213) -3, (1018) 0 --> (1218) -3:NW0, PEGB2, -, NW0
			8'd22 : rdata = 43'b0001001000000000111000001000001000000000000;
			// PEs: 8, 9 -> 10
			// srcs: (286, 22)(809) 0, (90) -3 --> (896) 0:PENB, ND1, *, PENB
			8'd23 : rdata = 43'b0001111011111110011000000010000000100000000;
			// PEs: 9, 10 -> 9
			// srcs: (295, 26)(291) 1, (1096) 0 --> (1296) 1:NW1, PEGB2, -, NW1
			8'd24 : rdata = 43'b0001001000000001111000001000001010000000000;
			// PEs: 8, 9 -> 10
			// srcs: (315, 23)(809) 0, (119) -1 --> (925) 0:PENB, ND3, *, PENB
			8'd25 : rdata = 43'b0001111011111110011000000110000000100000000;
			// PEs: 9, 10 -> 9
			// srcs: (324, 27)(320) -3, (1125) 0 --> (1325) -3:NW3, PEGB2, -, NW3
			8'd26 : rdata = 43'b0001001000000011111000001000001110000000000;
			// PEs: 8, 9 -> 10
			// srcs: (364, 24)(809) 0, (168) -1 --> (974) 0:PENB, ND2, *, PENB
			8'd27 : rdata = 43'b0001111011111110011000000100000000100000000;
			// PEs: 9, 10 -> 9
			// srcs: (373, 28)(369) 0, (1174) 0 --> (1374) 0:NW2, PEGB2, -, NW2
			8'd28 : rdata = 43'b0001001000000010111000001000001100000000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 10) begin
	always @(*) begin
		case(address)
			// PEs: 10, 10 -> 10
			// srcs: (1, 0)(14) -3, (215) -1 --> (415) 3:ND0, NW0, *, NI0
			8'd0 : rdata = 43'b0001101100000000010000000001000000000000000;
			// PEs: 10, 10 -> 11
			// srcs: (2, 1)(92) 1, (293) -2 --> (493) -2:ND1, NW1, *, PENB
			8'd1 : rdata = 43'b0001101100000001010000000010000000100000000;
			// PEs: 10, 10 -> 14
			// srcs: (3, 2)(170) -2, (371) -3 --> (571) 6:ND2, NW2, *, PEGB6
			8'd2 : rdata = 43'b0001101100000010010000000100000000011100000;
			// PEs: 10, 10 -> 10
			// srcs: (4, 3)(122) -3, (323) -2 --> (523) 6:ND3, NW3, *, NI1
			8'd3 : rdata = 43'b0001101100000011010000000111010000000000000;
			// PEs: 10, 11 -> 8
			// srcs: (7, 4)(415) 3, (416) 1 --> (613) 4:NI0, PEGB3, +, PEGB0
			8'd4 : rdata = 43'b0000110100000000111000001100000000010000000;
			// PEs: 10 -> 8
			// srcs: (18, 5)(523) 6 --> (523) 6:NI1, pass, PEGB0
			8'd5 : rdata = 43'b1100010100000001000000000000000000010000000;
			// PEs: 9 -> 
			// srcs: (34, 6)(693) 9 --> (693) 9:PENB, pass, 
			8'd6 : rdata = 43'b1100011011111110000000000000000000000000000;
			// PEs: 9, 10 -> 8
			// srcs: (41, 7)(691) -9, (693) 9 --> (694) 0:PENB, ALU, +, PEGB0
			8'd7 : rdata = 43'b0000111011111110001111111110000000010000000;
			// PEs: 10, 9 -> 9
			// srcs: (212, 12)(3) 1, (818) 0 --> (1018) 0:NM0, PENB, *, PEGB1
			8'd8 : rdata = 43'b0001110000000000110111111100000000010010000;
			// PEs: 8, 10 -> 11
			// srcs: (214, 8)(809) 0, (14) -3 --> (820) 0:PEGB0, ND0, *, PENB
			8'd9 : rdata = 43'b0001111100000000011000000000000000100000000;
			// PEs: 10, 11 -> 10
			// srcs: (223, 17)(215) -1, (1020) 0 --> (1220) -1:NW0, PEGB3, -, NW0
			8'd10 : rdata = 43'b0001001000000000111000001100001000000000000;
			// PEs: 10, 9 -> 9
			// srcs: (289, 13)(3) 1, (896) 0 --> (1096) 0:NM0, PENB, *, PEGB1
			8'd11 : rdata = 43'b0001110000000000110111111100000000010010000;
			// PEs: 8, 10 -> 11
			// srcs: (291, 9)(809) 0, (92) 1 --> (898) 0:PEGB0, ND1, *, PENB
			8'd12 : rdata = 43'b0001111100000000011000000010000000100000000;
			// PEs: 10, 11 -> 10
			// srcs: (300, 18)(293) -2, (1098) 0 --> (1298) -2:NW1, PEGB3, -, NW1
			8'd13 : rdata = 43'b0001001000000001111000001100001010000000000;
			// PEs: 10, 9 -> 9
			// srcs: (318, 14)(3) 1, (925) 0 --> (1125) 0:NM0, PENB, *, PEGB1
			8'd14 : rdata = 43'b0001110000000000110111111100000000010010000;
			// PEs: 8, 10 -> 
			// srcs: (321, 10)(809) 0, (122) -3 --> (928) 0:PEGB0, ND3, *, 
			8'd15 : rdata = 43'b0001111100000000011000000110000000000000000;
			// PEs: 10, 10 -> 
			// srcs: (324, 15)(3) 1, (928) 0 --> (1128) 0:NM0, ALU, *, 
			8'd16 : rdata = 43'b0001110000000000001111111110000000000000000;
			// PEs: 10, 10 -> 10
			// srcs: (327, 19)(323) -2, (1128) 0 --> (1328) -2:NW3, ALU, -, NW3
			8'd17 : rdata = 43'b0001001000000011001111111110001110000000000;
			// PEs: 10, 9 -> 9
			// srcs: (367, 16)(3) 1, (974) 0 --> (1174) 0:NM0, PENB, *, PEGB1
			8'd18 : rdata = 43'b0001110000000000110111111100000000010010000;
			// PEs: 8, 10 -> 11
			// srcs: (369, 11)(809) 0, (170) -2 --> (976) 0:PEGB0, ND2, *, PENB
			8'd19 : rdata = 43'b0001111100000000011000000100000000100000000;
			// PEs: 10, 11 -> 10
			// srcs: (378, 20)(371) -3, (1176) 0 --> (1376) -3:NW2, PEGB3, -, NW2
			8'd20 : rdata = 43'b0001001000000010111000001100001100000000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 11) begin
	always @(*) begin
		case(address)
			// PEs: 11, 11 -> 10
			// srcs: (1, 0)(15) 1, (216) 1 --> (416) 1:ND0, NW0, *, PEGB2
			8'd0 : rdata = 43'b0001101100000000010000000000000000010100000;
			// PEs: 11, 11 -> 11
			// srcs: (2, 1)(93) -3, (294) 2 --> (494) -6:ND1, NW1, *, NI0
			8'd1 : rdata = 43'b0001101100000001010000000011000000000000000;
			// PEs: 11, 11 -> 14
			// srcs: (3, 2)(171) 1, (372) 0 --> (572) 0:ND2, NW2, *, PEGB6
			8'd2 : rdata = 43'b0001101100000010010000000100000000011100000;
			// PEs: 11, 11 -> 8
			// srcs: (4, 3)(125) -1, (326) 2 --> (526) -2:ND3, NW3, *, PEGB0
			8'd3 : rdata = 43'b0001101100000011010000000110000000010000000;
			// PEs: 10, 11 -> 9
			// srcs: (5, 6)(493) -2, (494) -6 --> (690) -8:PENB, NI0, +, PEGB1
			8'd4 : rdata = 43'b0000111011111110101000000000000000010010000;
			// PEs: 13 -> 
			// srcs: (6, 4)(419) 0 --> (419) 0:PEGB5, pass, 
			8'd5 : rdata = 43'b1100011100001010000000000000000000000000000;
			// PEs: 12, 11 -> 8
			// srcs: (9, 5)(418) -1, (419) 0 --> (617) -1:PEGB4, ALU, +, PEGB0
			8'd6 : rdata = 43'b0000111100001000001111111110000000010000000;
			// PEs: 8, 11 -> 12
			// srcs: (215, 7)(809) 0, (15) 1 --> (821) 0:PEGB0, ND0, *, PENB
			8'd7 : rdata = 43'b0001111100000000011000000000000000100000000;
			// PEs: 11, 10 -> 10
			// srcs: (217, 11)(3) 1, (820) 0 --> (1020) 0:NM0, PENB, *, PEGB2
			8'd8 : rdata = 43'b0001110000000000110111111100000000010100000;
			// PEs: 11, 12 -> 11
			// srcs: (224, 15)(216) 1, (1021) 0 --> (1221) 1:NW0, PEGB4, -, NW0
			8'd9 : rdata = 43'b0001001000000000111000010000001000000000000;
			// PEs: 8, 11 -> 12
			// srcs: (292, 8)(809) 0, (93) -3 --> (899) 0:PEGB0, ND1, *, PENB
			8'd10 : rdata = 43'b0001111100000000011000000010000000100000000;
			// PEs: 11, 10 -> 10
			// srcs: (294, 12)(3) 1, (898) 0 --> (1098) 0:NM0, PENB, *, PEGB2
			8'd11 : rdata = 43'b0001110000000000110111111100000000010100000;
			// PEs: 11, 12 -> 11
			// srcs: (301, 16)(294) 2, (1099) 0 --> (1299) 2:NW1, PEGB4, -, NW1
			8'd12 : rdata = 43'b0001001000000001111000010000001010000000000;
			// PEs: 8, 11 -> 
			// srcs: (324, 9)(809) 0, (125) -1 --> (931) 0:PEGB0, ND3, *, 
			8'd13 : rdata = 43'b0001111100000000011000000110000000000000000;
			// PEs: 11, 11 -> 
			// srcs: (327, 13)(3) 1, (931) 0 --> (1131) 0:NM0, ALU, *, 
			8'd14 : rdata = 43'b0001110000000000001111111110000000000000000;
			// PEs: 11, 11 -> 11
			// srcs: (330, 17)(326) 2, (1131) 0 --> (1331) 2:NW3, ALU, -, NW3
			8'd15 : rdata = 43'b0001001000000011001111111110001110000000000;
			// PEs: 8, 11 -> 12
			// srcs: (370, 10)(809) 0, (171) 1 --> (977) 0:PEGB0, ND2, *, PENB
			8'd16 : rdata = 43'b0001111100000000011000000100000000100000000;
			// PEs: 11, 10 -> 10
			// srcs: (372, 14)(3) 1, (976) 0 --> (1176) 0:NM0, PENB, *, PEGB2
			8'd17 : rdata = 43'b0001110000000000110111111100000000010100000;
			// PEs: 11, 12 -> 11
			// srcs: (379, 18)(372) 0, (1177) 0 --> (1377) 0:NW2, PEGB4, -, NW2
			8'd18 : rdata = 43'b0001001000000010111000010000001100000000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 12) begin
	always @(*) begin
		case(address)
			// PEs: 12, 12 -> 11
			// srcs: (1, 0)(17) -1, (218) 1 --> (418) -1:ND0, NW0, *, PEGB3
			8'd0 : rdata = 43'b0001101100000000010000000000000000010110000;
			// PEs: 12, 12 -> 13
			// srcs: (2, 1)(95) -2, (296) -3 --> (496) 6:ND1, NW1, *, PENB
			8'd1 : rdata = 43'b0001101100000001010000000010000000100000000;
			// PEs: 12, 12 -> 13
			// srcs: (3, 2)(173) -3, (374) 0 --> (574) 0:ND2, NW2, *, PENB
			8'd2 : rdata = 43'b0001101100000010010000000100000000100000000;
			// PEs: 12, 12 -> 12
			// srcs: (4, 3)(128) -3, (329) 2 --> (529) -6:ND3, NW3, *, NI0
			8'd3 : rdata = 43'b0001101100000011010000000111000000000000000;
			// PEs: 15 -> 
			// srcs: (6, 4)(422) 0 --> (422) 0:PEGB7, pass, 
			8'd4 : rdata = 43'b1100011100001110000000000000000000000000000;
			// PEs: 14, 12 -> 8
			// srcs: (9, 5)(421) -2, (422) 0 --> (619) -2:PEGB6, ALU, +, PEGB0
			8'd5 : rdata = 43'b0000111100001100001111111110000000010000000;
			// PEs: 12 -> 8
			// srcs: (27, 6)(529) -6 --> (529) -6:NI0, pass, PEGB0
			8'd6 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 8, 12 -> 13
			// srcs: (216, 7)(809) 0, (17) -1 --> (823) 0:PEGB0, ND0, *, PENB
			8'd7 : rdata = 43'b0001111100000000011000000000000000100000000;
			// PEs: 12, 11 -> 11
			// srcs: (218, 11)(3) 1, (821) 0 --> (1021) 0:NM0, PENB, *, PEGB3
			8'd8 : rdata = 43'b0001110000000000110111111100000000010110000;
			// PEs: 12, 13 -> 12
			// srcs: (225, 15)(218) 1, (1023) 0 --> (1223) 1:NW0, PEGB5, -, NW0
			8'd9 : rdata = 43'b0001001000000000111000010100001000000000000;
			// PEs: 8, 12 -> 13
			// srcs: (294, 8)(809) 0, (95) -2 --> (901) 0:PEGB0, ND1, *, PENB
			8'd10 : rdata = 43'b0001111100000000011000000010000000100000000;
			// PEs: 12, 11 -> 11
			// srcs: (295, 12)(3) 1, (899) 0 --> (1099) 0:NM0, PENB, *, PEGB3
			8'd11 : rdata = 43'b0001110000000000110111111100000000010110000;
			// PEs: 12, 13 -> 12
			// srcs: (303, 16)(296) -3, (1101) 0 --> (1301) -3:NW1, PEGB5, -, NW1
			8'd12 : rdata = 43'b0001001000000001111000010100001010000000000;
			// PEs: 8, 12 -> 
			// srcs: (327, 9)(809) 0, (128) -3 --> (934) 0:PEGB0, ND3, *, 
			8'd13 : rdata = 43'b0001111100000000011000000110000000000000000;
			// PEs: 12, 12 -> 
			// srcs: (330, 13)(3) 1, (934) 0 --> (1134) 0:NM0, ALU, *, 
			8'd14 : rdata = 43'b0001110000000000001111111110000000000000000;
			// PEs: 12, 12 -> 12
			// srcs: (333, 17)(329) 2, (1134) 0 --> (1334) 2:NW3, ALU, -, NW3
			8'd15 : rdata = 43'b0001001000000011001111111110001110000000000;
			// PEs: 8, 12 -> 13
			// srcs: (372, 10)(809) 0, (173) -3 --> (979) 0:PEGB0, ND2, *, PENB
			8'd16 : rdata = 43'b0001111100000000011000000100000000100000000;
			// PEs: 12, 11 -> 11
			// srcs: (373, 14)(3) 1, (977) 0 --> (1177) 0:NM0, PENB, *, PEGB3
			8'd17 : rdata = 43'b0001110000000000110111111100000000010110000;
			// PEs: 12, 13 -> 12
			// srcs: (381, 18)(374) 0, (1179) 0 --> (1379) 0:NW2, PEGB5, -, NW2
			8'd18 : rdata = 43'b0001001000000010111000010100001100000000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 13) begin
	always @(*) begin
		case(address)
			// PEs: 13, 13 -> 11
			// srcs: (1, 0)(18) 0, (219) -3 --> (419) 0:ND0, NW0, *, PEGB3
			8'd0 : rdata = 43'b0001101100000000010000000000000000010110000;
			// PEs: 13, 13 -> 13
			// srcs: (2, 1)(96) -1, (297) 1 --> (497) -1:ND1, NW1, *, NI0
			8'd1 : rdata = 43'b0001101100000001010000000011000000000000000;
			// PEs: 13, 13 -> 13
			// srcs: (3, 2)(174) 0, (375) 0 --> (575) 0:ND2, NW2, *, NI1
			8'd2 : rdata = 43'b0001101100000010010000000101010000000000000;
			// PEs: 13, 13 -> 8
			// srcs: (4, 3)(135) 2, (336) 0 --> (536) 0:ND3, NW3, *, PEGB0
			8'd3 : rdata = 43'b0001101100000011010000000110000000010000000;
			// PEs: 12, 13 -> 9
			// srcs: (5, 4)(496) 6, (497) -1 --> (692) 5:PENB, NI0, +, PEGB1
			8'd4 : rdata = 43'b0000111011111110101000000000000000010010000;
			// PEs: 12, 13 -> 8
			// srcs: (6, 5)(574) 0, (575) 0 --> (770) 0:PENB, NI1, +, PEGB0
			8'd5 : rdata = 43'b0000111011111110101000000010000000010000000;
			// PEs: 8, 13 -> 14
			// srcs: (217, 6)(809) 0, (18) 0 --> (824) 0:PEGB0, ND0, *, PENB
			8'd6 : rdata = 43'b0001111100000000011000000000000000100000000;
			// PEs: 13, 12 -> 12
			// srcs: (219, 10)(3) 1, (823) 0 --> (1023) 0:NM0, PENB, *, PEGB4
			8'd7 : rdata = 43'b0001110000000000110111111100000000011000000;
			// PEs: 13, 14 -> 13
			// srcs: (226, 15)(219) -3, (1024) 0 --> (1224) -3:NW0, PEGB6, -, NW0
			8'd8 : rdata = 43'b0001001000000000111000011000001000000000000;
			// PEs: 8, 13 -> 13
			// srcs: (295, 7)(809) 0, (96) -1 --> (902) 0:PEGB0, ND1, *, NI0
			8'd9 : rdata = 43'b0001111100000000011000000011000000000000000;
			// PEs: 13, 12 -> 12
			// srcs: (297, 11)(3) 1, (901) 0 --> (1101) 0:NM0, PENB, *, PEGB4
			8'd10 : rdata = 43'b0001110000000000110111111100000000011000000;
			// PEs: 13, 13 -> 
			// srcs: (298, 12)(3) 1, (902) 0 --> (1102) 0:NM0, NI0, *, 
			8'd11 : rdata = 43'b0001110000000000101000000000000000000000000;
			// PEs: 13, 13 -> 13
			// srcs: (301, 16)(297) 1, (1102) 0 --> (1302) 1:NW1, ALU, -, NW1
			8'd12 : rdata = 43'b0001001000000001001111111110001010000000000;
			// PEs: 8, 13 -> 
			// srcs: (334, 8)(809) 0, (135) 2 --> (941) 0:PEGB0, ND3, *, 
			8'd13 : rdata = 43'b0001111100000000011000000110000000000000000;
			// PEs: 13, 13 -> 
			// srcs: (337, 13)(3) 1, (941) 0 --> (1141) 0:NM0, ALU, *, 
			8'd14 : rdata = 43'b0001110000000000001111111110000000000000000;
			// PEs: 13, 13 -> 13
			// srcs: (340, 17)(336) 0, (1141) 0 --> (1341) 0:NW3, ALU, -, NW3
			8'd15 : rdata = 43'b0001001000000011001111111110001110000000000;
			// PEs: 8, 13 -> 14
			// srcs: (373, 9)(809) 0, (174) 0 --> (980) 0:PEGB0, ND2, *, PENB
			8'd16 : rdata = 43'b0001111100000000011000000100000000100000000;
			// PEs: 13, 12 -> 12
			// srcs: (375, 14)(3) 1, (979) 0 --> (1179) 0:NM0, PENB, *, PEGB4
			8'd17 : rdata = 43'b0001110000000000110111111100000000011000000;
			// PEs: 13, 14 -> 13
			// srcs: (382, 18)(375) 0, (1180) 0 --> (1380) 0:NW2, PEGB6, -, NW2
			8'd18 : rdata = 43'b0001001000000010111000011000001100000000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 14) begin
	always @(*) begin
		case(address)
			// PEs: 14, 14 -> 12
			// srcs: (1, 0)(20) -1, (221) 2 --> (421) -2:ND0, NW0, *, PEGB4
			8'd0 : rdata = 43'b0001101100000000010000000000000000011000000;
			// PEs: 14, 14 -> 15
			// srcs: (2, 1)(98) 0, (299) -1 --> (499) 0:ND1, NW1, *, PENB
			8'd1 : rdata = 43'b0001101100000001010000000010000000100000000;
			// PEs: 14, 14 -> 15
			// srcs: (3, 2)(176) -2, (377) 1 --> (577) -2:ND2, NW2, *, PENB
			8'd2 : rdata = 43'b0001101100000010010000000100000000100000000;
			// PEs: 14, 14 -> 9
			// srcs: (4, 3)(138) -2, (339) -2 --> (539) 4:ND3, NW3, *, PEGB1
			8'd3 : rdata = 43'b0001101100000011010000000110000000010010000;
			// PEs: 11 -> 
			// srcs: (8, 4)(572) 0 --> (572) 0:PEGB3, pass, 
			8'd4 : rdata = 43'b1100011100000110000000000000000000000000000;
			// PEs: 10, 14 -> 8
			// srcs: (11, 5)(571) 6, (572) 0 --> (767) 6:PEGB2, ALU, +, PEGB0
			8'd5 : rdata = 43'b0000111100000100001111111110000000010000000;
			// PEs: 8, 14 -> 14
			// srcs: (219, 6)(809) 0, (20) -1 --> (826) 0:PEGB0, ND0, *, NI0
			8'd6 : rdata = 43'b0001111100000000011000000001000000000000000;
			// PEs: 14, 13 -> 13
			// srcs: (220, 10)(3) 1, (824) 0 --> (1024) 0:NM0, PENB, *, PEGB5
			8'd7 : rdata = 43'b0001110000000000110111111100000000011010000;
			// PEs: 14, 14 -> 
			// srcs: (222, 11)(3) 1, (826) 0 --> (1026) 0:NM0, NI0, *, 
			8'd8 : rdata = 43'b0001110000000000101000000000000000000000000;
			// PEs: 14, 14 -> 14
			// srcs: (225, 16)(221) 2, (1026) 0 --> (1226) 2:NW0, ALU, -, NW0
			8'd9 : rdata = 43'b0001001000000000001111111110001000000000000;
			// PEs: 8, 14 -> 
			// srcs: (297, 7)(809) 0, (98) 0 --> (904) 0:PEGB0, ND1, *, 
			8'd10 : rdata = 43'b0001111100000000011000000010000000000000000;
			// PEs: 14, 14 -> 
			// srcs: (300, 12)(3) 1, (904) 0 --> (1104) 0:NM0, ALU, *, 
			8'd11 : rdata = 43'b0001110000000000001111111110000000000000000;
			// PEs: 14, 14 -> 14
			// srcs: (303, 17)(299) -1, (1104) 0 --> (1304) -1:NW1, ALU, -, NW1
			8'd12 : rdata = 43'b0001001000000001001111111110001010000000000;
			// PEs: 8, 14 -> 
			// srcs: (337, 8)(809) 0, (138) -2 --> (944) 0:PEGB0, ND3, *, 
			8'd13 : rdata = 43'b0001111100000000011000000110000000000000000;
			// PEs: 14, 14 -> 
			// srcs: (340, 13)(3) 1, (944) 0 --> (1144) 0:NM0, ALU, *, 
			8'd14 : rdata = 43'b0001110000000000001111111110000000000000000;
			// PEs: 14, 14 -> 14
			// srcs: (343, 18)(339) -2, (1144) 0 --> (1344) -2:NW3, ALU, -, NW3
			8'd15 : rdata = 43'b0001001000000011001111111110001110000000000;
			// PEs: 8, 14 -> 14
			// srcs: (375, 9)(809) 0, (176) -2 --> (982) 0:PEGB0, ND2, *, NI0
			8'd16 : rdata = 43'b0001111100000000011000000101000000000000000;
			// PEs: 14, 13 -> 13
			// srcs: (376, 14)(3) 1, (980) 0 --> (1180) 0:NM0, PENB, *, PEGB5
			8'd17 : rdata = 43'b0001110000000000110111111100000000011010000;
			// PEs: 14, 14 -> 
			// srcs: (378, 15)(3) 1, (982) 0 --> (1182) 0:NM0, NI0, *, 
			8'd18 : rdata = 43'b0001110000000000101000000000000000000000000;
			// PEs: 14, 14 -> 14
			// srcs: (381, 19)(377) 1, (1182) 0 --> (1382) 1:NW2, ALU, -, NW2
			8'd19 : rdata = 43'b0001001000000010001111111110001100000000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 15) begin
	always @(*) begin
		case(address)
			// PEs: 15, 15 -> 12
			// srcs: (1, 0)(21) 0, (222) -1 --> (422) 0:ND0, NW0, *, PEGB4
			8'd0 : rdata = 43'b0001101100000000010000000000000000011000000;
			// PEs: 15, 15 -> 15
			// srcs: (2, 1)(99) 1, (300) 0 --> (500) 0:ND1, NW1, *, NI0
			8'd1 : rdata = 43'b0001101100000001010000000011000000000000000;
			// PEs: 15, 15 -> 15
			// srcs: (3, 2)(177) -2, (378) 0 --> (578) 0:ND2, NW2, *, NI1
			8'd2 : rdata = 43'b0001101100000010010000000101010000000000000;
			// PEs: 15, 15 -> 15
			// srcs: (4, 3)(141) -3, (342) 0 --> (542) 0:ND3, NW3, *, NI2
			8'd3 : rdata = 43'b0001101100000011010000000111100000000000000;
			// PEs: 14, 15 -> 8
			// srcs: (5, 4)(499) 0, (500) 0 --> (695) 0:PENB, NI0, +, PENB
			8'd4 : rdata = 43'b0000111011111110101000000000000000100000000;
			// PEs: 14, 15 -> 15
			// srcs: (6, 5)(577) -2, (578) 0 --> (772) -2:PENB, NI1, +, NI0
			8'd5 : rdata = 43'b0000111011111110101000000011000000000000000;
			// PEs: 15 -> 8
			// srcs: (12, 6)(542) 0 --> (542) 0:NI2, pass, PENB
			8'd6 : rdata = 43'b1100010100000010000000000000000000100000000;
			// PEs: 15 -> 8
			// srcs: (24, 7)(772) -2 --> (772) -2:NI0, pass, PENB
			8'd7 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 8, 15 -> 
			// srcs: (220, 8)(809) 0, (21) 0 --> (827) 0:PEGB0, ND0, *, 
			8'd8 : rdata = 43'b0001111100000000011000000000000000000000000;
			// PEs: 15, 15 -> 
			// srcs: (223, 12)(3) 1, (827) 0 --> (1027) 0:NM0, ALU, *, 
			8'd9 : rdata = 43'b0001110000000000001111111110000000000000000;
			// PEs: 15, 15 -> 15
			// srcs: (226, 16)(222) -1, (1027) 0 --> (1227) -1:NW0, ALU, -, NW0
			8'd10 : rdata = 43'b0001001000000000001111111110001000000000000;
			// PEs: 8, 15 -> 
			// srcs: (298, 9)(809) 0, (99) 1 --> (905) 0:PEGB0, ND1, *, 
			8'd11 : rdata = 43'b0001111100000000011000000010000000000000000;
			// PEs: 15, 15 -> 
			// srcs: (301, 13)(3) 1, (905) 0 --> (1105) 0:NM0, ALU, *, 
			8'd12 : rdata = 43'b0001110000000000001111111110000000000000000;
			// PEs: 15, 15 -> 15
			// srcs: (304, 17)(300) 0, (1105) 0 --> (1305) 0:NW1, ALU, -, NW1
			8'd13 : rdata = 43'b0001001000000001001111111110001010000000000;
			// PEs: 8, 15 -> 
			// srcs: (340, 10)(809) 0, (141) -3 --> (947) 0:PEGB0, ND3, *, 
			8'd14 : rdata = 43'b0001111100000000011000000110000000000000000;
			// PEs: 15, 15 -> 
			// srcs: (343, 14)(3) 1, (947) 0 --> (1147) 0:NM0, ALU, *, 
			8'd15 : rdata = 43'b0001110000000000001111111110000000000000000;
			// PEs: 15, 15 -> 15
			// srcs: (346, 18)(342) 0, (1147) 0 --> (1347) 0:NW3, ALU, -, NW3
			8'd16 : rdata = 43'b0001001000000011001111111110001110000000000;
			// PEs: 8, 15 -> 
			// srcs: (376, 11)(809) 0, (177) -2 --> (983) 0:PEGB0, ND2, *, 
			8'd17 : rdata = 43'b0001111100000000011000000100000000000000000;
			// PEs: 15, 15 -> 
			// srcs: (379, 15)(3) 1, (983) 0 --> (1183) 0:NM0, ALU, *, 
			8'd18 : rdata = 43'b0001110000000000001111111110000000000000000;
			// PEs: 15, 15 -> 15
			// srcs: (382, 19)(378) 0, (1183) 0 --> (1383) 0:NW2, ALU, -, NW2
			8'd19 : rdata = 43'b0001001000000010001111111110001100000000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 16) begin
	always @(*) begin
		case(address)
			// PEs: 23 -> 24
			// srcs: (4, 0)(509) 0 --> (509) 0:PENB, pass, PUNB
			8'd0 : rdata = 43'b1100011011111110000000000000000001000000000;
			// PEs: 23 -> 24
			// srcs: (5, 1)(587) 0 --> (587) 0:PENB, pass, PUNB
			8'd1 : rdata = 43'b1100011011111110000000000000000001000000000;
			// PEs: 18 -> 32
			// srcs: (9, 20)(548) 0 --> (548) 0:PEGB2, pass, PUGB4
			8'd2 : rdata = 43'b1100011100000100000000000000000000000001100;
			// PEs: 23 -> 24
			// srcs: (10, 2)(432) 0 --> (432) 0:PENB, pass, PUNB
			8'd3 : rdata = 43'b1100011011111110000000000000000001000000000;
			// PEs: 32 -> 16
			// srcs: (11, 4)(417) -6 --> (417) -6:PUGB4, pass, NI0
			8'd4 : rdata = 43'b1100011100001001000000000001000000000000000;
			// PEs: 17 -> 48
			// srcs: (12, 6)(622) 1 --> (622) 1:PEGB1, pass, PUGB6
			8'd5 : rdata = 43'b1100011100000010000000000000000000000001110;
			// PEs: 18 -> 40
			// srcs: (13, 12)(697) -1 --> (697) -1:PEGB2, pass, PUGB5
			8'd6 : rdata = 43'b1100011100000100000000000000000000000001101;
			// PEs: 8 -> 17
			// srcs: (14, 3)(613) 4 --> (613) 4:PUNB, pass, PENB
			8'd7 : rdata = 43'b1100011011111111000000000000000000100000000;
			// PEs: 18 -> 56
			// srcs: (15, 7)(624) 2 --> (624) 2:PEGB2, pass, PUGB7
			8'd8 : rdata = 43'b1100011100000100000000000000000000000001111;
			// PEs: 19 -> 24
			// srcs: (16, 8)(629) -1 --> (629) -1:PEGB3, pass, PUNB
			8'd9 : rdata = 43'b1100011100000110000000000000000001000000000;
			// PEs: 20 -> 40
			// srcs: (17, 22)(554) 0 --> (554) 0:PEGB4, pass, PUGB5
			8'd10 : rdata = 43'b1100011100001000000000000000000000000001101;
			// PEs: 21 -> 0
			// srcs: (18, 23)(561) 2 --> (561) 2:PEGB5, pass, PUGB0
			8'd11 : rdata = 43'b1100011100001010000000000000000000000001000;
			// PEs: 16 -> 17
			// srcs: (21, 5)(417) -6 --> (417) -6:NI0, pass, PENB
			8'd12 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 32 -> 16
			// srcs: (22, 9)(641) 8 --> (641) 8:PUGB4, pass, NI0
			8'd13 : rdata = 43'b1100011100001001000000000001000000000000000;
			// PEs: 48 -> 17
			// srcs: (23, 10)(445) 4 --> (445) 4:PUGB6, pass, PENB
			8'd14 : rdata = 43'b1100011100001101000000000000000000100000000;
			// PEs: 17 -> 56
			// srcs: (24, 19)(545) -3 --> (545) -3:PEGB1, pass, PUGB7
			8'd15 : rdata = 43'b1100011100000010000000000000000000000001111;
			// PEs: 19 -> 48
			// srcs: (25, 21)(551) 9 --> (551) 9:PEGB3, pass, PUGB6
			8'd16 : rdata = 43'b1100011100000110000000000000000000000001110;
			// PEs: 22 -> 56
			// srcs: (26, 24)(564) -4 --> (564) -4:PEGB6, pass, PUGB7
			8'd17 : rdata = 43'b1100011100001100000000000000000000000001111;
			// PEs: 23 -> 0
			// srcs: (27, 25)(567) 0 --> (567) 0:PENB, pass, PUGB0
			8'd18 : rdata = 43'b1100011011111110000000000000000000000001000;
			// PEs: 22 -> 24
			// srcs: (28, 26)(780) -1 --> (780) -1:PEGB6, pass, PUNB
			8'd19 : rdata = 43'b1100011100001100000000000000000001000000000;
			// PEs: 16 -> 17
			// srcs: (29, 11)(641) 8 --> (641) 8:NI0, pass, PENB
			8'd20 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 24 -> 16
			// srcs: (30, 13)(710) 1 --> (710) 1:PUGB3, pass, NI0
			8'd21 : rdata = 43'b1100011100000111000000000001000000000000000;
			// PEs: 0 -> 17
			// srcs: (31, 14)(514) -4 --> (514) -4:PUGB0, pass, PENB
			8'd22 : rdata = 43'b1100011100000001000000000000000000100000000;
			// PEs: 17 -> 40
			// srcs: (32, 27)(614) -2 --> (614) -2:PEGB1, pass, PUGB5
			8'd23 : rdata = 43'b1100011100000010000000000000000000000001101;
			// PEs: 17 -> 0
			// srcs: (36, 28)(642) 12 --> (642) 12:PEGB1, pass, PUGB0
			8'd24 : rdata = 43'b1100011100000010000000000000000000000001000;
			// PEs: 16 -> 17
			// srcs: (37, 15)(710) 1 --> (710) 1:NI0, pass, PENB
			8'd25 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 24 -> 16
			// srcs: (38, 16)(716) 7 --> (716) 7:PUGB3, pass, NI0
			8'd26 : rdata = 43'b1100011100000111000000000001000000000000000;
			// PEs: 8 -> 17
			// srcs: (39, 17)(520) 3 --> (520) 3:PUNB, pass, PENB
			8'd27 : rdata = 43'b1100011011111111000000000000000000100000000;
			// PEs: 23 -> 56
			// srcs: (40, 32)(706) 1 --> (706) 1:PENB, pass, PUGB7
			8'd28 : rdata = 43'b1100011011111110000000000000000000000001111;
			// PEs: 17 -> 24
			// srcs: (44, 33)(711) -3 --> (711) -3:PEGB1, pass, PUNB
			8'd29 : rdata = 43'b1100011100000010000000000000000001000000000;
			// PEs: 16 -> 17
			// srcs: (45, 18)(716) 7 --> (716) 7:NI0, pass, PENB
			8'd30 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 16
			// srcs: (46, 29)(696) 9 --> (696) 9:PUGB0, pass, NI0
			8'd31 : rdata = 43'b1100011100000001000000000001000000000000000;
			// PEs: 21 -> 24
			// srcs: (47, 38)(779) -1 --> (779) -1:PEGB5, pass, PUNB
			8'd32 : rdata = 43'b1100011100001010000000000000000001000000000;
			// PEs: 40 -> 17
			// srcs: (48, 30)(698) 1 --> (698) 1:PUGB5, pass, PENB
			8'd33 : rdata = 43'b1100011100001011000000000000000000100000000;
			// PEs: 17 -> 40
			// srcs: (52, 34)(717) 10 --> (717) 10:PEGB1, pass, PUGB5
			8'd34 : rdata = 43'b1100011100000010000000000000000000000001101;
			// PEs: 16 -> 17
			// srcs: (55, 31)(696) 9 --> (696) 9:NI0, pass, PENB
			8'd35 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 8 -> 16
			// srcs: (56, 35)(735) 2 --> (735) 2:PUNB, pass, NI0
			8'd36 : rdata = 43'b1100011011111111000000000001000000000000000;
			// PEs: 48 -> 17
			// srcs: (57, 36)(737) 1 --> (737) 1:PUGB6, pass, PENB
			8'd37 : rdata = 43'b1100011100001101000000000000000000100000000;
			// PEs: 16 -> 17
			// srcs: (63, 37)(735) 2 --> (735) 2:NI0, pass, PENB
			8'd38 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 8 -> 17
			// srcs: (64, 39)(694) 0 --> (694) 0:PUNB, pass, PENB
			8'd39 : rdata = 43'b1100011011111111000000000000000000100000000;
			// PEs: 17 -> 48
			// srcs: (70, 40)(738) 3 --> (738) 3:PEGB1, pass, PUGB6
			8'd40 : rdata = 43'b1100011100000010000000000000000000000001110;
			// PEs: 8 -> 16
			// srcs: (80, 41)(640) 11 --> (640) 11:PUNB, pass, NI0
			8'd41 : rdata = 43'b1100011011111111000000000001000000000000000;
			// PEs: 48 -> 17
			// srcs: (83, 42)(651) 10 --> (651) 10:PUGB6, pass, PENB
			8'd42 : rdata = 43'b1100011100001101000000000000000000100000000;
			// PEs: 16 -> 17
			// srcs: (90, 43)(640) 11 --> (640) 11:NI0, pass, PENB
			8'd43 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 8 -> 17
			// srcs: (91, 44)(689) -12 --> (689) -12:PUNB, pass, PENB
			8'd44 : rdata = 43'b1100011011111111000000000000000000100000000;
			// PEs: 8 -> 17
			// srcs: (98, 45)(628) 0 --> (628) 0:PUNB, pass, PENB
			8'd45 : rdata = 43'b1100011011111111000000000000000000100000000;
			// PEs: 17 -> 24
			// srcs: (99, 46)(701) -2 --> (701) -2:PEGB1, pass, PUNB
			8'd46 : rdata = 43'b1100011100000010000000000000000001000000000;
			// PEs: 17 -> 24
			// srcs: (107, 47)(653) 21 --> (653) 21:PEGB1, pass, PUNB
			8'd47 : rdata = 43'b1100011100000010000000000000000001000000000;
			// PEs: 32 -> 17
			// srcs: (217, 48)(809) 0 --> (809) 0:PUGB4, pass, PENB
			8'd48 : rdata = 43'b1100011100001001000000000000000000100000000;
			// PEs: 32 -> 18
			// srcs: (218, 49)(809) 0 --> (809) 0:PUGB4, pass, PEGB2
			8'd49 : rdata = 43'b1100011100001001000000000000000000010100000;
			// PEs: 32 -> 19
			// srcs: (220, 50)(809) 0 --> (809) 0:PUGB4, pass, PEGB3
			8'd50 : rdata = 43'b1100011100001001000000000000000000010110000;
			// PEs: 32 -> 20
			// srcs: (221, 51)(809) 0 --> (809) 0:PUGB4, pass, PEGB4
			8'd51 : rdata = 43'b1100011100001001000000000000000000011000000;
			// PEs: 32 -> 21
			// srcs: (223, 52)(809) 0 --> (809) 0:PUGB4, pass, PEGB5
			8'd52 : rdata = 43'b1100011100001001000000000000000000011010000;
			// PEs: 32 -> 22
			// srcs: (224, 53)(809) 0 --> (809) 0:PUGB4, pass, PEGB6
			8'd53 : rdata = 43'b1100011100001001000000000000000000011100000;
			// PEs: 32 -> 23
			// srcs: (225, 54)(809) 0 --> (809) 0:PUGB4, pass, PEGB7
			8'd54 : rdata = 43'b1100011100001001000000000000000000011110000;
			// PEs: 32 -> 17
			// srcs: (295, 55)(809) 0 --> (809) 0:PUGB4, pass, PENB
			8'd55 : rdata = 43'b1100011100001001000000000000000000100000000;
			// PEs: 32 -> 18
			// srcs: (296, 56)(809) 0 --> (809) 0:PUGB4, pass, PEGB2
			8'd56 : rdata = 43'b1100011100001001000000000000000000010100000;
			// PEs: 32 -> 19
			// srcs: (298, 57)(809) 0 --> (809) 0:PUGB4, pass, PEGB3
			8'd57 : rdata = 43'b1100011100001001000000000000000000010110000;
			// PEs: 32 -> 20
			// srcs: (299, 58)(809) 0 --> (809) 0:PUGB4, pass, PEGB4
			8'd58 : rdata = 43'b1100011100001001000000000000000000011000000;
			// PEs: 32 -> 21
			// srcs: (300, 59)(809) 0 --> (809) 0:PUGB4, pass, PEGB5
			8'd59 : rdata = 43'b1100011100001001000000000000000000011010000;
			// PEs: 32 -> 22
			// srcs: (301, 60)(809) 0 --> (809) 0:PUGB4, pass, PEGB6
			8'd60 : rdata = 43'b1100011100001001000000000000000000011100000;
			// PEs: 32 -> 23
			// srcs: (302, 61)(809) 0 --> (809) 0:PUGB4, pass, PEGB7
			8'd61 : rdata = 43'b1100011100001001000000000000000000011110000;
			// PEs: 32 -> 17
			// srcs: (338, 62)(809) 0 --> (809) 0:PUGB4, pass, PENB
			8'd62 : rdata = 43'b1100011100001001000000000000000000100000000;
			// PEs: 32 -> 18
			// srcs: (341, 63)(809) 0 --> (809) 0:PUGB4, pass, PEGB2
			8'd63 : rdata = 43'b1100011100001001000000000000000000010100000;
			// PEs: 32 -> 19
			// srcs: (344, 64)(809) 0 --> (809) 0:PUGB4, pass, PEGB3
			8'd64 : rdata = 43'b1100011100001001000000000000000000010110000;
			// PEs: 32 -> 20
			// srcs: (347, 65)(809) 0 --> (809) 0:PUGB4, pass, PEGB4
			8'd65 : rdata = 43'b1100011100001001000000000000000000011000000;
			// PEs: 32 -> 21
			// srcs: (354, 66)(809) 0 --> (809) 0:PUGB4, pass, PEGB5
			8'd66 : rdata = 43'b1100011100001001000000000000000000011010000;
			// PEs: 32 -> 22
			// srcs: (357, 67)(809) 0 --> (809) 0:PUGB4, pass, PEGB6
			8'd67 : rdata = 43'b1100011100001001000000000000000000011100000;
			// PEs: 32 -> 23
			// srcs: (360, 68)(809) 0 --> (809) 0:PUGB4, pass, PEGB7
			8'd68 : rdata = 43'b1100011100001001000000000000000000011110000;
			// PEs: 32 -> 17
			// srcs: (373, 69)(809) 0 --> (809) 0:PUGB4, pass, PENB
			8'd69 : rdata = 43'b1100011100001001000000000000000000100000000;
			// PEs: 32 -> 18
			// srcs: (374, 70)(809) 0 --> (809) 0:PUGB4, pass, PEGB2
			8'd70 : rdata = 43'b1100011100001001000000000000000000010100000;
			// PEs: 32 -> 19
			// srcs: (375, 71)(809) 0 --> (809) 0:PUGB4, pass, PEGB3
			8'd71 : rdata = 43'b1100011100001001000000000000000000010110000;
			// PEs: 32 -> 20
			// srcs: (376, 72)(809) 0 --> (809) 0:PUGB4, pass, PEGB4
			8'd72 : rdata = 43'b1100011100001001000000000000000000011000000;
			// PEs: 32 -> 21
			// srcs: (377, 73)(809) 0 --> (809) 0:PUGB4, pass, PEGB5
			8'd73 : rdata = 43'b1100011100001001000000000000000000011010000;
			// PEs: 32 -> 22
			// srcs: (378, 74)(809) 0 --> (809) 0:PUGB4, pass, PEGB6
			8'd74 : rdata = 43'b1100011100001001000000000000000000011100000;
			// PEs: 32 -> 23
			// srcs: (380, 75)(809) 0 --> (809) 0:PUGB4, pass, PEGB7
			8'd75 : rdata = 43'b1100011100001001000000000000000000011110000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 17) begin
	always @(*) begin
		case(address)
			// PEs: 17, 17 -> 17
			// srcs: (1, 0)(23) 1, (224) -1 --> (424) -1:ND0, NW0, *, NI0
			8'd0 : rdata = 43'b0001101100000000010000000001000000000000000;
			// PEs: 17, 17 -> 18
			// srcs: (2, 1)(101) 0, (302) 2 --> (502) 0:ND1, NW1, *, PENB
			8'd1 : rdata = 43'b0001101100000001010000000010000000100000000;
			// PEs: 17, 17 -> 21
			// srcs: (3, 2)(179) 2, (380) 0 --> (580) 0:ND2, NW2, *, PEGB5
			8'd2 : rdata = 43'b0001101100000010010000000100000000011010000;
			// PEs: 17, 17 -> 17
			// srcs: (4, 3)(144) 1, (345) -3 --> (545) -3:ND3, NW3, *, NI1
			8'd3 : rdata = 43'b0001101100000011010000000111010000000000000;
			// PEs: 17, 18 -> 16
			// srcs: (7, 4)(424) -1, (425) 2 --> (622) 1:NI0, PEGB2, +, PEGB0
			8'd4 : rdata = 43'b0000110100000000111000001000000000010000000;
			// PEs: 16 -> 17
			// srcs: (16, 5)(613) 4 --> (613) 4:PENB, pass, NI0
			8'd5 : rdata = 43'b1100011011111110000000000001000000000000000;
			// PEs: 17 -> 16
			// srcs: (19, 13)(545) -3 --> (545) -3:NI1, pass, PEGB0
			8'd6 : rdata = 43'b1100010100000001000000000000000000010000000;
			// PEs: 17, 16 -> 16
			// srcs: (23, 6)(613) 4, (417) -6 --> (614) -2:NI0, PENB, +, PEGB0
			8'd7 : rdata = 43'b0000110100000000110111111100000000010000000;
			// PEs: 16 -> 
			// srcs: (25, 7)(445) 4 --> (445) 4:PENB, pass, 
			8'd8 : rdata = 43'b1100011011111110000000000000000000000000000;
			// PEs: 16, 17 -> 16
			// srcs: (31, 8)(641) 8, (445) 4 --> (642) 12:PENB, ALU, +, PEGB0
			8'd9 : rdata = 43'b0000111011111110001111111110000000010000000;
			// PEs: 16 -> 
			// srcs: (33, 9)(514) -4 --> (514) -4:PENB, pass, 
			8'd10 : rdata = 43'b1100011011111110000000000000000000000000000;
			// PEs: 16, 17 -> 16
			// srcs: (39, 10)(710) 1, (514) -4 --> (711) -3:PENB, ALU, +, PEGB0
			8'd11 : rdata = 43'b0000111011111110001111111110000000010000000;
			// PEs: 16 -> 
			// srcs: (41, 11)(520) 3 --> (520) 3:PENB, pass, 
			8'd12 : rdata = 43'b1100011011111110000000000000000000000000000;
			// PEs: 16, 17 -> 16
			// srcs: (47, 12)(716) 7, (520) 3 --> (717) 10:PENB, ALU, +, PEGB0
			8'd13 : rdata = 43'b0000111011111110001111111110000000010000000;
			// PEs: 16 -> 
			// srcs: (50, 14)(698) 1 --> (698) 1:PENB, pass, 
			8'd14 : rdata = 43'b1100011011111110000000000000000000000000000;
			// PEs: 16, 17 -> 17
			// srcs: (57, 15)(696) 9, (698) 1 --> (699) 10:PENB, ALU, +, NI0
			8'd15 : rdata = 43'b0000111011111110001111111111000000000000000;
			// PEs: 16 -> 
			// srcs: (59, 16)(737) 1 --> (737) 1:PENB, pass, 
			8'd16 : rdata = 43'b1100011011111110000000000000000000000000000;
			// PEs: 16, 17 -> 16
			// srcs: (65, 17)(735) 2, (737) 1 --> (738) 3:PENB, ALU, +, PEGB0
			8'd17 : rdata = 43'b0000111011111110001111111110000000010000000;
			// PEs: 16, 17 -> 17
			// srcs: (67, 18)(694) 0, (699) 10 --> (700) 10:PENB, NI0, +, NI1
			8'd18 : rdata = 43'b0000111011111110101000000001010000000000000;
			// PEs: 16 -> 
			// srcs: (85, 19)(651) 10 --> (651) 10:PENB, pass, 
			8'd19 : rdata = 43'b1100011011111110000000000000000000000000000;
			// PEs: 16, 17 -> 17
			// srcs: (92, 20)(640) 11, (651) 10 --> (652) 21:PENB, ALU, +, NI0
			8'd20 : rdata = 43'b0000111011111110001111111111000000000000000;
			// PEs: 16, 17 -> 16
			// srcs: (93, 21)(689) -12, (700) 10 --> (701) -2:PENB, NI1, +, PEGB0
			8'd21 : rdata = 43'b0000111011111110101000000010000000010000000;
			// PEs: 16, 17 -> 16
			// srcs: (102, 22)(628) 0, (652) 21 --> (653) 21:PENB, NI0, +, PEGB0
			8'd22 : rdata = 43'b0000111011111110101000000000000000010000000;
			// PEs: 16, 17 -> 18
			// srcs: (219, 23)(809) 0, (23) 1 --> (829) 0:PENB, ND0, *, PENB
			8'd23 : rdata = 43'b0001111011111110011000000000000000100000000;
			// PEs: 17, 18 -> 17
			// srcs: (228, 27)(224) -1, (1029) 0 --> (1229) -1:NW0, PEGB2, -, NW0
			8'd24 : rdata = 43'b0001001000000000111000001000001000000000000;
			// PEs: 16, 17 -> 18
			// srcs: (297, 24)(809) 0, (101) 0 --> (907) 0:PENB, ND1, *, PENB
			8'd25 : rdata = 43'b0001111011111110011000000010000000100000000;
			// PEs: 17, 18 -> 17
			// srcs: (306, 28)(302) 2, (1107) 0 --> (1307) 2:NW1, PEGB2, -, NW1
			8'd26 : rdata = 43'b0001001000000001111000001000001010000000000;
			// PEs: 16, 17 -> 18
			// srcs: (340, 25)(809) 0, (144) 1 --> (950) 0:PENB, ND3, *, PENB
			8'd27 : rdata = 43'b0001111011111110011000000110000000100000000;
			// PEs: 17, 18 -> 17
			// srcs: (349, 29)(345) -3, (1150) 0 --> (1350) -3:NW3, PEGB2, -, NW3
			8'd28 : rdata = 43'b0001001000000011111000001000001110000000000;
			// PEs: 16, 17 -> 18
			// srcs: (375, 26)(809) 0, (179) 2 --> (985) 0:PENB, ND2, *, PENB
			8'd29 : rdata = 43'b0001111011111110011000000100000000100000000;
			// PEs: 17, 18 -> 17
			// srcs: (384, 30)(380) 0, (1185) 0 --> (1385) 0:NW2, PEGB2, -, NW2
			8'd30 : rdata = 43'b0001001000000010111000001000001100000000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 18) begin
	always @(*) begin
		case(address)
			// PEs: 18, 18 -> 17
			// srcs: (1, 0)(24) -2, (225) -1 --> (425) 2:ND0, NW0, *, PEGB1
			8'd0 : rdata = 43'b0001101100000000010000000000000000010010000;
			// PEs: 18, 18 -> 18
			// srcs: (2, 1)(102) 1, (303) -1 --> (503) -1:ND1, NW1, *, NI0
			8'd1 : rdata = 43'b0001101100000001010000000011000000000000000;
			// PEs: 18, 18 -> 21
			// srcs: (3, 2)(180) -1, (381) 2 --> (581) -2:ND2, NW2, *, PEGB5
			8'd2 : rdata = 43'b0001101100000010010000000100000000011010000;
			// PEs: 18, 18 -> 16
			// srcs: (4, 3)(147) 0, (348) 0 --> (548) 0:ND3, NW3, *, PEGB0
			8'd3 : rdata = 43'b0001101100000011010000000110000000010000000;
			// PEs: 17, 18 -> 16
			// srcs: (5, 6)(502) 0, (503) -1 --> (697) -1:PENB, NI0, +, PEGB0
			8'd4 : rdata = 43'b0000111011111110101000000000000000010000000;
			// PEs: 20 -> 
			// srcs: (6, 4)(428) 0 --> (428) 0:PEGB4, pass, 
			8'd5 : rdata = 43'b1100011100001000000000000000000000000000000;
			// PEs: 19, 18 -> 16
			// srcs: (9, 5)(427) 2, (428) 0 --> (624) 2:PEGB3, ALU, +, PEGB0
			8'd6 : rdata = 43'b0000111100000110001111111110000000010000000;
			// PEs: 18, 17 -> 17
			// srcs: (222, 11)(3) 1, (829) 0 --> (1029) 0:NM0, PENB, *, PEGB1
			8'd7 : rdata = 43'b0001110000000000110111111100000000010010000;
			// PEs: 16, 18 -> 19
			// srcs: (223, 7)(809) 0, (24) -2 --> (830) 0:PEGB0, ND0, *, PENB
			8'd8 : rdata = 43'b0001111100000000011000000000000000100000000;
			// PEs: 18, 19 -> 18
			// srcs: (232, 16)(225) -1, (1030) 0 --> (1230) -1:NW0, PEGB3, -, NW0
			8'd9 : rdata = 43'b0001001000000000111000001100001000000000000;
			// PEs: 18, 17 -> 17
			// srcs: (300, 12)(3) 1, (907) 0 --> (1107) 0:NM0, PENB, *, PEGB1
			8'd10 : rdata = 43'b0001110000000000110111111100000000010010000;
			// PEs: 16, 18 -> 19
			// srcs: (301, 8)(809) 0, (102) 1 --> (908) 0:PEGB0, ND1, *, PENB
			8'd11 : rdata = 43'b0001111100000000011000000010000000100000000;
			// PEs: 18, 19 -> 18
			// srcs: (310, 17)(303) -1, (1108) 0 --> (1308) -1:NW1, PEGB3, -, NW1
			8'd12 : rdata = 43'b0001001000000001111000001100001010000000000;
			// PEs: 18, 17 -> 17
			// srcs: (343, 13)(3) 1, (950) 0 --> (1150) 0:NM0, PENB, *, PEGB1
			8'd13 : rdata = 43'b0001110000000000110111111100000000010010000;
			// PEs: 16, 18 -> 
			// srcs: (346, 9)(809) 0, (147) 0 --> (953) 0:PEGB0, ND3, *, 
			8'd14 : rdata = 43'b0001111100000000011000000110000000000000000;
			// PEs: 18, 18 -> 
			// srcs: (349, 14)(3) 1, (953) 0 --> (1153) 0:NM0, ALU, *, 
			8'd15 : rdata = 43'b0001110000000000001111111110000000000000000;
			// PEs: 18, 18 -> 18
			// srcs: (352, 18)(348) 0, (1153) 0 --> (1353) 0:NW3, ALU, -, NW3
			8'd16 : rdata = 43'b0001001000000011001111111110001110000000000;
			// PEs: 18, 17 -> 17
			// srcs: (378, 15)(3) 1, (985) 0 --> (1185) 0:NM0, PENB, *, PEGB1
			8'd17 : rdata = 43'b0001110000000000110111111100000000010010000;
			// PEs: 16, 18 -> 19
			// srcs: (379, 10)(809) 0, (180) -1 --> (986) 0:PEGB0, ND2, *, PENB
			8'd18 : rdata = 43'b0001111100000000011000000100000000100000000;
			// PEs: 18, 19 -> 18
			// srcs: (388, 19)(381) 2, (1186) 0 --> (1386) 2:NW2, PEGB3, -, NW2
			8'd19 : rdata = 43'b0001001000000010111000001100001100000000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 19) begin
	always @(*) begin
		case(address)
			// PEs: 19, 19 -> 18
			// srcs: (1, 0)(26) -2, (227) -1 --> (427) 2:ND0, NW0, *, PEGB2
			8'd0 : rdata = 43'b0001101100000000010000000000000000010100000;
			// PEs: 19, 19 -> 20
			// srcs: (2, 1)(104) 1, (305) -1 --> (505) -1:ND1, NW1, *, PENB
			8'd1 : rdata = 43'b0001101100000001010000000010000000100000000;
			// PEs: 19, 19 -> 20
			// srcs: (3, 2)(181) 1, (382) 1 --> (582) 1:ND2, NW2, *, PENB
			8'd2 : rdata = 43'b0001101100000010010000000100000000100000000;
			// PEs: 19, 19 -> 19
			// srcs: (4, 3)(150) -3, (351) -3 --> (551) 9:ND3, NW3, *, NI0
			8'd3 : rdata = 43'b0001101100000011010000000111000000000000000;
			// PEs: 22 -> 
			// srcs: (6, 4)(431) 2 --> (431) 2:PEGB6, pass, 
			8'd4 : rdata = 43'b1100011100001100000000000000000000000000000;
			// PEs: 21, 19 -> 16
			// srcs: (9, 5)(430) -3, (431) 2 --> (629) -1:PEGB5, ALU, +, PEGB0
			8'd5 : rdata = 43'b0000111100001010001111111110000000010000000;
			// PEs: 19 -> 16
			// srcs: (19, 6)(551) 9 --> (551) 9:NI0, pass, PEGB0
			8'd6 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 16, 19 -> 20
			// srcs: (225, 7)(809) 0, (26) -2 --> (832) 0:PEGB0, ND0, *, PENB
			8'd7 : rdata = 43'b0001111100000000011000000000000000100000000;
			// PEs: 19, 18 -> 18
			// srcs: (226, 11)(3) 1, (830) 0 --> (1030) 0:NM0, PENB, *, PEGB2
			8'd8 : rdata = 43'b0001110000000000110111111100000000010100000;
			// PEs: 19, 20 -> 19
			// srcs: (234, 15)(227) -1, (1032) 0 --> (1232) -1:NW0, PEGB4, -, NW0
			8'd9 : rdata = 43'b0001001000000000111000010000001000000000000;
			// PEs: 16, 19 -> 20
			// srcs: (303, 8)(809) 0, (104) 1 --> (910) 0:PEGB0, ND1, *, PENB
			8'd10 : rdata = 43'b0001111100000000011000000010000000100000000;
			// PEs: 19, 18 -> 18
			// srcs: (304, 12)(3) 1, (908) 0 --> (1108) 0:NM0, PENB, *, PEGB2
			8'd11 : rdata = 43'b0001110000000000110111111100000000010100000;
			// PEs: 19, 20 -> 19
			// srcs: (312, 16)(305) -1, (1110) 0 --> (1310) -1:NW1, PEGB4, -, NW1
			8'd12 : rdata = 43'b0001001000000001111000010000001010000000000;
			// PEs: 16, 19 -> 
			// srcs: (349, 9)(809) 0, (150) -3 --> (956) 0:PEGB0, ND3, *, 
			8'd13 : rdata = 43'b0001111100000000011000000110000000000000000;
			// PEs: 19, 19 -> 
			// srcs: (352, 13)(3) 1, (956) 0 --> (1156) 0:NM0, ALU, *, 
			8'd14 : rdata = 43'b0001110000000000001111111110000000000000000;
			// PEs: 19, 19 -> 19
			// srcs: (355, 17)(351) -3, (1156) 0 --> (1356) -3:NW3, ALU, -, NW3
			8'd15 : rdata = 43'b0001001000000011001111111110001110000000000;
			// PEs: 16, 19 -> 20
			// srcs: (380, 10)(809) 0, (181) 1 --> (987) 0:PEGB0, ND2, *, PENB
			8'd16 : rdata = 43'b0001111100000000011000000100000000100000000;
			// PEs: 19, 18 -> 18
			// srcs: (382, 14)(3) 1, (986) 0 --> (1186) 0:NM0, PENB, *, PEGB2
			8'd17 : rdata = 43'b0001110000000000110111111100000000010100000;
			// PEs: 19, 20 -> 19
			// srcs: (389, 18)(382) 1, (1187) 0 --> (1387) 1:NW2, PEGB4, -, NW2
			8'd18 : rdata = 43'b0001001000000010111000010000001100000000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 20) begin
	always @(*) begin
		case(address)
			// PEs: 20, 20 -> 18
			// srcs: (1, 0)(27) 0, (228) 0 --> (428) 0:ND0, NW0, *, PEGB2
			8'd0 : rdata = 43'b0001101100000000010000000000000000010100000;
			// PEs: 20, 20 -> 20
			// srcs: (2, 1)(105) 1, (306) 2 --> (506) 2:ND1, NW1, *, NI0
			8'd1 : rdata = 43'b0001101100000001010000000011000000000000000;
			// PEs: 20, 20 -> 20
			// srcs: (3, 2)(182) 0, (383) -2 --> (583) 0:ND2, NW2, *, NI1
			8'd2 : rdata = 43'b0001101100000010010000000101010000000000000;
			// PEs: 20, 20 -> 16
			// srcs: (4, 3)(153) 0, (354) 1 --> (554) 0:ND3, NW3, *, PEGB0
			8'd3 : rdata = 43'b0001101100000011010000000110000000010000000;
			// PEs: 19, 20 -> 23
			// srcs: (5, 4)(505) -1, (506) 2 --> (704) 1:PENB, NI0, +, PEGB7
			8'd4 : rdata = 43'b0000111011111110101000000000000000011110000;
			// PEs: 19, 20 -> 21
			// srcs: (6, 5)(582) 1, (583) 0 --> (778) 1:PENB, NI1, +, PENB
			8'd5 : rdata = 43'b0000111011111110101000000010000000100000000;
			// PEs: 16, 20 -> 20
			// srcs: (226, 6)(809) 0, (27) 0 --> (833) 0:PEGB0, ND0, *, NI0
			8'd6 : rdata = 43'b0001111100000000011000000001000000000000000;
			// PEs: 20, 19 -> 19
			// srcs: (228, 10)(3) 1, (832) 0 --> (1032) 0:NM0, PENB, *, PEGB3
			8'd7 : rdata = 43'b0001110000000000110111111100000000010110000;
			// PEs: 20, 20 -> 
			// srcs: (229, 11)(3) 1, (833) 0 --> (1033) 0:NM0, NI0, *, 
			8'd8 : rdata = 43'b0001110000000000101000000000000000000000000;
			// PEs: 20, 20 -> 20
			// srcs: (232, 15)(228) 0, (1033) 0 --> (1233) 0:NW0, ALU, -, NW0
			8'd9 : rdata = 43'b0001001000000000001111111110001000000000000;
			// PEs: 16, 20 -> 21
			// srcs: (304, 7)(809) 0, (105) 1 --> (911) 0:PEGB0, ND1, *, PENB
			8'd10 : rdata = 43'b0001111100000000011000000010000000100000000;
			// PEs: 20, 19 -> 19
			// srcs: (306, 12)(3) 1, (910) 0 --> (1110) 0:NM0, PENB, *, PEGB3
			8'd11 : rdata = 43'b0001110000000000110111111100000000010110000;
			// PEs: 20, 21 -> 20
			// srcs: (313, 16)(306) 2, (1111) 0 --> (1311) 2:NW1, PEGB5, -, NW1
			8'd12 : rdata = 43'b0001001000000001111000010100001010000000000;
			// PEs: 16, 20 -> 
			// srcs: (352, 8)(809) 0, (153) 0 --> (959) 0:PEGB0, ND3, *, 
			8'd13 : rdata = 43'b0001111100000000011000000110000000000000000;
			// PEs: 20, 20 -> 
			// srcs: (355, 13)(3) 1, (959) 0 --> (1159) 0:NM0, ALU, *, 
			8'd14 : rdata = 43'b0001110000000000001111111110000000000000000;
			// PEs: 20, 20 -> 20
			// srcs: (358, 17)(354) 1, (1159) 0 --> (1359) 1:NW3, ALU, -, NW3
			8'd15 : rdata = 43'b0001001000000011001111111110001110000000000;
			// PEs: 16, 20 -> 21
			// srcs: (381, 9)(809) 0, (182) 0 --> (988) 0:PEGB0, ND2, *, PENB
			8'd16 : rdata = 43'b0001111100000000011000000100000000100000000;
			// PEs: 20, 19 -> 19
			// srcs: (383, 14)(3) 1, (987) 0 --> (1187) 0:NM0, PENB, *, PEGB3
			8'd17 : rdata = 43'b0001110000000000110111111100000000010110000;
			// PEs: 20, 21 -> 20
			// srcs: (390, 18)(383) -2, (1188) 0 --> (1388) -2:NW2, PEGB5, -, NW2
			8'd18 : rdata = 43'b0001001000000010111000010100001100000000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 21) begin
	always @(*) begin
		case(address)
			// PEs: 21, 21 -> 19
			// srcs: (1, 0)(29) -3, (230) 1 --> (430) -3:ND0, NW0, *, PEGB3
			8'd0 : rdata = 43'b0001101100000000010000000000000000010110000;
			// PEs: 21, 21 -> 22
			// srcs: (2, 1)(106) -2, (307) -3 --> (507) 6:ND1, NW1, *, PENB
			8'd1 : rdata = 43'b0001101100000001010000000010000000100000000;
			// PEs: 21, 21 -> 22
			// srcs: (3, 2)(183) 1, (384) -1 --> (584) -1:ND2, NW2, *, PENB
			8'd2 : rdata = 43'b0001101100000010010000000100000000100000000;
			// PEs: 21, 21 -> 16
			// srcs: (4, 3)(160) 2, (361) 1 --> (561) 2:ND3, NW3, *, PEGB0
			8'd3 : rdata = 43'b0001101100000011010000000110000000010000000;
			// PEs: 18 -> 
			// srcs: (8, 4)(581) -2 --> (581) -2:PEGB2, pass, 
			8'd4 : rdata = 43'b1100011100000100000000000000000000000000000;
			// PEs: 17, 21 -> 
			// srcs: (11, 5)(580) 0, (581) -2 --> (777) -2:PEGB1, ALU, +, 
			8'd5 : rdata = 43'b0000111100000010001111111110000000000000000;
			// PEs: 21, 20 -> 16
			// srcs: (14, 6)(777) -2, (778) 1 --> (779) -1:ALU, PENB, +, PEGB0
			8'd6 : rdata = 43'b0000100111111111110111111100000000010000000;
			// PEs: 16, 21 -> 22
			// srcs: (228, 7)(809) 0, (29) -3 --> (835) 0:PEGB0, ND0, *, PENB
			8'd7 : rdata = 43'b0001111100000000011000000000000000100000000;
			// PEs: 21, 22 -> 21
			// srcs: (237, 15)(230) 1, (1035) 0 --> (1235) 1:NW0, PEGB6, -, NW0
			8'd8 : rdata = 43'b0001001000000000111000011000001000000000000;
			// PEs: 16, 21 -> 21
			// srcs: (305, 8)(809) 0, (106) -2 --> (912) 0:PEGB0, ND1, *, NI0
			8'd9 : rdata = 43'b0001111100000000011000000011000000000000000;
			// PEs: 21, 20 -> 20
			// srcs: (307, 11)(3) 1, (911) 0 --> (1111) 0:NM0, PENB, *, PEGB4
			8'd10 : rdata = 43'b0001110000000000110111111100000000011000000;
			// PEs: 21, 21 -> 
			// srcs: (308, 12)(3) 1, (912) 0 --> (1112) 0:NM0, NI0, *, 
			8'd11 : rdata = 43'b0001110000000000101000000000000000000000000;
			// PEs: 21, 21 -> 21
			// srcs: (311, 16)(307) -3, (1112) 0 --> (1312) -3:NW1, ALU, -, NW1
			8'd12 : rdata = 43'b0001001000000001001111111110001010000000000;
			// PEs: 16, 21 -> 
			// srcs: (359, 9)(809) 0, (160) 2 --> (966) 0:PEGB0, ND3, *, 
			8'd13 : rdata = 43'b0001111100000000011000000110000000000000000;
			// PEs: 21, 21 -> 
			// srcs: (362, 13)(3) 1, (966) 0 --> (1166) 0:NM0, ALU, *, 
			8'd14 : rdata = 43'b0001110000000000001111111110000000000000000;
			// PEs: 21, 21 -> 21
			// srcs: (365, 17)(361) 1, (1166) 0 --> (1366) 1:NW3, ALU, -, NW3
			8'd15 : rdata = 43'b0001001000000011001111111110001110000000000;
			// PEs: 16, 21 -> 22
			// srcs: (382, 10)(809) 0, (183) 1 --> (989) 0:PEGB0, ND2, *, PENB
			8'd16 : rdata = 43'b0001111100000000011000000100000000100000000;
			// PEs: 21, 20 -> 20
			// srcs: (384, 14)(3) 1, (988) 0 --> (1188) 0:NM0, PENB, *, PEGB4
			8'd17 : rdata = 43'b0001110000000000110111111100000000011000000;
			// PEs: 21, 22 -> 21
			// srcs: (391, 18)(384) -1, (1189) 0 --> (1389) -1:NW2, PEGB6, -, NW2
			8'd18 : rdata = 43'b0001001000000010111000011000001100000000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 22) begin
	always @(*) begin
		case(address)
			// PEs: 22, 22 -> 19
			// srcs: (1, 0)(30) 2, (231) 1 --> (431) 2:ND0, NW0, *, PEGB3
			8'd0 : rdata = 43'b0001101100000000010000000000000000010110000;
			// PEs: 22, 22 -> 22
			// srcs: (2, 1)(107) 2, (308) -3 --> (508) -6:ND1, NW1, *, NI0
			8'd1 : rdata = 43'b0001101100000001010000000011000000000000000;
			// PEs: 22, 22 -> 22
			// srcs: (3, 2)(184) 1, (385) 0 --> (585) 0:ND2, NW2, *, NI1
			8'd2 : rdata = 43'b0001101100000010010000000101010000000000000;
			// PEs: 22, 22 -> 16
			// srcs: (4, 3)(163) 2, (364) -2 --> (564) -4:ND3, NW3, *, PEGB0
			8'd3 : rdata = 43'b0001101100000011010000000110000000010000000;
			// PEs: 21, 22 -> 23
			// srcs: (5, 5)(507) 6, (508) -6 --> (705) 0:PENB, NI0, +, PENB
			8'd4 : rdata = 43'b0000111011111110101000000000000000100000000;
			// PEs: 21, 22 -> 16
			// srcs: (6, 4)(584) -1, (585) 0 --> (780) -1:PENB, NI1, +, PEGB0
			8'd5 : rdata = 43'b0000111011111110101000000010000000010000000;
			// PEs: 16, 22 -> 22
			// srcs: (229, 6)(809) 0, (30) 2 --> (836) 0:PEGB0, ND0, *, NI0
			8'd6 : rdata = 43'b0001111100000000011000000001000000000000000;
			// PEs: 22, 21 -> 21
			// srcs: (231, 10)(3) 1, (835) 0 --> (1035) 0:NM0, PENB, *, PEGB5
			8'd7 : rdata = 43'b0001110000000000110111111100000000011010000;
			// PEs: 22, 22 -> 
			// srcs: (232, 11)(3) 1, (836) 0 --> (1036) 0:NM0, NI0, *, 
			8'd8 : rdata = 43'b0001110000000000101000000000000000000000000;
			// PEs: 22, 22 -> 22
			// srcs: (235, 16)(231) 1, (1036) 0 --> (1236) 1:NW0, ALU, -, NW0
			8'd9 : rdata = 43'b0001001000000000001111111110001000000000000;
			// PEs: 16, 22 -> 
			// srcs: (306, 7)(809) 0, (107) 2 --> (913) 0:PEGB0, ND1, *, 
			8'd10 : rdata = 43'b0001111100000000011000000010000000000000000;
			// PEs: 22, 22 -> 
			// srcs: (309, 12)(3) 1, (913) 0 --> (1113) 0:NM0, ALU, *, 
			8'd11 : rdata = 43'b0001110000000000001111111110000000000000000;
			// PEs: 22, 22 -> 22
			// srcs: (312, 17)(308) -3, (1113) 0 --> (1313) -3:NW1, ALU, -, NW1
			8'd12 : rdata = 43'b0001001000000001001111111110001010000000000;
			// PEs: 16, 22 -> 
			// srcs: (362, 8)(809) 0, (163) 2 --> (969) 0:PEGB0, ND3, *, 
			8'd13 : rdata = 43'b0001111100000000011000000110000000000000000;
			// PEs: 22, 22 -> 
			// srcs: (365, 13)(3) 1, (969) 0 --> (1169) 0:NM0, ALU, *, 
			8'd14 : rdata = 43'b0001110000000000001111111110000000000000000;
			// PEs: 22, 22 -> 22
			// srcs: (368, 18)(364) -2, (1169) 0 --> (1369) -2:NW3, ALU, -, NW3
			8'd15 : rdata = 43'b0001001000000011001111111110001110000000000;
			// PEs: 16, 22 -> 22
			// srcs: (383, 9)(809) 0, (184) 1 --> (990) 0:PEGB0, ND2, *, NI0
			8'd16 : rdata = 43'b0001111100000000011000000101000000000000000;
			// PEs: 22, 21 -> 21
			// srcs: (385, 14)(3) 1, (989) 0 --> (1189) 0:NM0, PENB, *, PEGB5
			8'd17 : rdata = 43'b0001110000000000110111111100000000011010000;
			// PEs: 22, 22 -> 
			// srcs: (386, 15)(3) 1, (990) 0 --> (1190) 0:NM0, NI0, *, 
			8'd18 : rdata = 43'b0001110000000000101000000000000000000000000;
			// PEs: 22, 22 -> 22
			// srcs: (389, 19)(385) 0, (1190) 0 --> (1390) 0:NW2, ALU, -, NW2
			8'd19 : rdata = 43'b0001001000000010001111111110001100000000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 23) begin
	always @(*) begin
		case(address)
			// PEs: 23, 23 -> 23
			// srcs: (1, 0)(31) 0, (232) 1 --> (432) 0:ND0, NW0, *, NI0
			8'd0 : rdata = 43'b0001101100000000010000000001000000000000000;
			// PEs: 23, 23 -> 16
			// srcs: (2, 1)(108) 1, (309) 0 --> (509) 0:ND1, NW1, *, PENB
			8'd1 : rdata = 43'b0001101100000001010000000010000000100000000;
			// PEs: 23, 23 -> 16
			// srcs: (3, 2)(186) 0, (387) -2 --> (587) 0:ND2, NW2, *, PENB
			8'd2 : rdata = 43'b0001101100000010010000000100000000100000000;
			// PEs: 23, 23 -> 23
			// srcs: (4, 3)(166) 1, (367) 0 --> (567) 0:ND3, NW3, *, NI1
			8'd3 : rdata = 43'b0001101100000011010000000111010000000000000;
			// PEs: 23 -> 16
			// srcs: (8, 4)(432) 0 --> (432) 0:NI0, pass, PENB
			8'd4 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 20, 22 -> 23
			// srcs: (11, 5)(704) 1, (705) 0 --> (706) 1:PEGB4, PENB, +, NI0
			8'd5 : rdata = 43'b0000111100001000110111111101000000000000000;
			// PEs: 23 -> 16
			// srcs: (21, 6)(567) 0 --> (567) 0:NI1, pass, PENB
			8'd6 : rdata = 43'b1100010100000001000000000000000000100000000;
			// PEs: 23 -> 16
			// srcs: (35, 7)(706) 1 --> (706) 1:NI0, pass, PENB
			8'd7 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 16, 23 -> 
			// srcs: (230, 8)(809) 0, (31) 0 --> (837) 0:PEGB0, ND0, *, 
			8'd8 : rdata = 43'b0001111100000000011000000000000000000000000;
			// PEs: 23, 23 -> 
			// srcs: (233, 12)(3) 1, (837) 0 --> (1037) 0:NM0, ALU, *, 
			8'd9 : rdata = 43'b0001110000000000001111111110000000000000000;
			// PEs: 23, 23 -> 23
			// srcs: (236, 16)(232) 1, (1037) 0 --> (1237) 1:NW0, ALU, -, NW0
			8'd10 : rdata = 43'b0001001000000000001111111110001000000000000;
			// PEs: 16, 23 -> 
			// srcs: (307, 9)(809) 0, (108) 1 --> (914) 0:PEGB0, ND1, *, 
			8'd11 : rdata = 43'b0001111100000000011000000010000000000000000;
			// PEs: 23, 23 -> 
			// srcs: (310, 13)(3) 1, (914) 0 --> (1114) 0:NM0, ALU, *, 
			8'd12 : rdata = 43'b0001110000000000001111111110000000000000000;
			// PEs: 23, 23 -> 23
			// srcs: (313, 17)(309) 0, (1114) 0 --> (1314) 0:NW1, ALU, -, NW1
			8'd13 : rdata = 43'b0001001000000001001111111110001010000000000;
			// PEs: 16, 23 -> 
			// srcs: (365, 10)(809) 0, (166) 1 --> (972) 0:PEGB0, ND3, *, 
			8'd14 : rdata = 43'b0001111100000000011000000110000000000000000;
			// PEs: 23, 23 -> 
			// srcs: (368, 14)(3) 1, (972) 0 --> (1172) 0:NM0, ALU, *, 
			8'd15 : rdata = 43'b0001110000000000001111111110000000000000000;
			// PEs: 23, 23 -> 23
			// srcs: (371, 18)(367) 0, (1172) 0 --> (1372) 0:NW3, ALU, -, NW3
			8'd16 : rdata = 43'b0001001000000011001111111110001110000000000;
			// PEs: 16, 23 -> 
			// srcs: (385, 11)(809) 0, (186) 0 --> (992) 0:PEGB0, ND2, *, 
			8'd17 : rdata = 43'b0001111100000000011000000100000000000000000;
			// PEs: 23, 23 -> 
			// srcs: (388, 15)(3) 1, (992) 0 --> (1192) 0:NM0, ALU, *, 
			8'd18 : rdata = 43'b0001110000000000001111111110000000000000000;
			// PEs: 23, 23 -> 23
			// srcs: (391, 19)(387) -2, (1192) 0 --> (1392) -2:NW2, ALU, -, NW2
			8'd19 : rdata = 43'b0001001000000010001111111110001100000000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 24) begin
	always @(*) begin
		case(address)
			// PEs: 16 -> 28
			// srcs: (6, 0)(509) 0 --> (509) 0:PUNB, pass, PEGB4
			8'd0 : rdata = 43'b1100011011111111000000000000000000011000000;
			// PEs: 16 -> 25
			// srcs: (7, 1)(587) 0 --> (587) 0:PUNB, pass, PENB
			8'd1 : rdata = 43'b1100011011111111000000000000000000100000000;
			// PEs: 27 -> 16
			// srcs: (10, 8)(710) 1 --> (710) 1:PEGB3, pass, PUGB2
			8'd2 : rdata = 43'b1100011100000110000000000000000000000001010;
			// PEs: 31 -> 16
			// srcs: (11, 10)(716) 7 --> (716) 7:PENB, pass, PUGB2
			8'd3 : rdata = 43'b1100011011111110000000000000000000000001010;
			// PEs: 25 -> 0
			// srcs: (14, 4)(632) 2 --> (632) 2:PEGB1, pass, PUGB0
			8'd4 : rdata = 43'b1100011100000010000000000000000000000001000;
			// PEs: 26 -> 8
			// srcs: (15, 5)(635) 4 --> (635) 4:PEGB2, pass, PUGB1
			8'd5 : rdata = 43'b1100011100000100000000000000000000000001001;
			// PEs: 27 -> 32
			// srcs: (16, 6)(637) 9 --> (637) 9:PEGB3, pass, PUNB
			8'd6 : rdata = 43'b1100011100000110000000000000000001000000000;
			// PEs: 16 -> 25
			// srcs: (17, 2)(432) 0 --> (432) 0:PUNB, pass, PENB
			8'd7 : rdata = 43'b1100011011111111000000000000000000100000000;
			// PEs: 16 -> 25
			// srcs: (18, 3)(629) -1 --> (629) -1:PUNB, pass, PENB
			8'd8 : rdata = 43'b1100011011111111000000000000000000100000000;
			// PEs: 28 -> 56
			// srcs: (19, 7)(707) -4 --> (707) -4:PEGB4, pass, PUGB7
			8'd9 : rdata = 43'b1100011100001000000000000000000000000001111;
			// PEs: 0 -> 25
			// srcs: (20, 9)(517) 0 --> (517) 0:PUGB0, pass, PENB
			8'd10 : rdata = 43'b1100011100000001000000000000000000100000000;
			// PEs: 32 -> 24
			// srcs: (21, 11)(721) 8 --> (721) 8:PUGB4, pass, NI0
			8'd11 : rdata = 43'b1100011100001001000000000001000000000000000;
			// PEs: 8 -> 25
			// srcs: (22, 12)(526) -2 --> (526) -2:PUGB1, pass, PENB
			8'd12 : rdata = 43'b1100011100000011000000000000000000100000000;
			// PEs: 27 -> 32
			// srcs: (30, 16)(576) 1 --> (576) 1:PEGB3, pass, PUNB
			8'd13 : rdata = 43'b1100011100000110000000000000000001000000000;
			// PEs: 29 -> 32
			// srcs: (31, 19)(789) -4 --> (789) -4:PEGB5, pass, PUNB
			8'd14 : rdata = 43'b1100011100001010000000000000000001000000000;
			// PEs: 31 -> 32
			// srcs: (32, 20)(791) 3 --> (791) 3:PENB, pass, PUNB
			8'd15 : rdata = 43'b1100011011111110000000000000000001000000000;
			// PEs: 24 -> 25
			// srcs: (34, 13)(721) 8 --> (721) 8:NI0, pass, PENB
			8'd16 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 8 -> 25
			// srcs: (35, 14)(765) -1 --> (765) -1:PUGB1, pass, PENB
			8'd17 : rdata = 43'b1100011100000011000000000000000000100000000;
			// PEs: 8 -> 25
			// srcs: (36, 15)(767) 6 --> (767) 6:PUGB1, pass, PENB
			8'd18 : rdata = 43'b1100011100000011000000000000000000100000000;
			// PEs: 25 -> 48
			// srcs: (37, 21)(631) -3 --> (631) -3:PEGB1, pass, PUGB6
			8'd19 : rdata = 43'b1100011100000010000000000000000000000001110;
			// PEs: 25 -> 32
			// srcs: (41, 23)(722) 6 --> (722) 6:PEGB1, pass, PUNB
			8'd20 : rdata = 43'b1100011100000010000000000000000001000000000;
			// PEs: 8 -> 25
			// srcs: (47, 17)(772) -2 --> (772) -2:PUGB1, pass, PENB
			8'd21 : rdata = 43'b1100011100000011000000000000000000100000000;
			// PEs: 16 -> 25
			// srcs: (48, 18)(780) -1 --> (780) -1:PUNB, pass, PENB
			8'd22 : rdata = 43'b1100011011111111000000000000000000100000000;
			// PEs: 16 -> 28
			// srcs: (49, 22)(711) -3 --> (711) -3:PUNB, pass, PEGB4
			8'd23 : rdata = 43'b1100011011111111000000000000000000011000000;
			// PEs: 25 -> 32
			// srcs: (54, 27)(773) -2 --> (773) -2:PEGB1, pass, PUNB
			8'd24 : rdata = 43'b1100011100000010000000000000000001000000000;
			// PEs: 26 -> 32
			// srcs: (55, 31)(769) 8 --> (769) 8:PEGB2, pass, PUNB
			8'd25 : rdata = 43'b1100011100000100000000000000000001000000000;
			// PEs: 56 -> 24
			// srcs: (60, 24)(741) -2 --> (741) -2:PUGB7, pass, NI0
			8'd26 : rdata = 43'b1100011100001111000000000001000000000000000;
			// PEs: 28 -> 56
			// srcs: (61, 29)(714) 8 --> (714) 8:PEGB4, pass, PUGB7
			8'd27 : rdata = 43'b1100011100001000000000000000000000000001111;
			// PEs: 32 -> 25
			// srcs: (78, 25)(743) 9 --> (743) 9:PUGB4, pass, PENB
			8'd28 : rdata = 43'b1100011100001001000000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (85, 26)(741) -2 --> (741) -2:NI0, pass, PENB
			8'd29 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 16 -> 25
			// srcs: (86, 28)(779) -1 --> (779) -1:PUNB, pass, PENB
			8'd30 : rdata = 43'b1100011011111111000000000000000000100000000;
			// PEs: 25 -> 56
			// srcs: (92, 30)(744) 7 --> (744) 7:PEGB1, pass, PUGB7
			8'd31 : rdata = 43'b1100011100000010000000000000000000000001111;
			// PEs: 29 -> 32
			// srcs: (101, 32)(788) -13 --> (788) -13:PEGB5, pass, PUNB
			8'd32 : rdata = 43'b1100011100001010000000000000000001000000000;
			// PEs: 56 -> 24
			// srcs: (117, 33)(677) 16 --> (677) 16:PUGB7, pass, NI0
			8'd33 : rdata = 43'b1100011100001111000000000001000000000000000;
			// PEs: 16 -> 25
			// srcs: (118, 34)(701) -2 --> (701) -2:PUNB, pass, PENB
			8'd34 : rdata = 43'b1100011011111111000000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (124, 35)(677) 16 --> (677) 16:NI0, pass, PENB
			8'd35 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 16 -> 25
			// srcs: (125, 36)(653) 21 --> (653) 21:PUNB, pass, PENB
			8'd36 : rdata = 43'b1100011011111111000000000000000000100000000;
			// PEs: 25 -> 0
			// srcs: (141, 37)(703) 35 --> (703) 35:PEGB1, pass, PUGB0
			8'd37 : rdata = 43'b1100011100000010000000000000000000000001000;
			// PEs: 32 -> 25
			// srcs: (226, 38)(809) 0 --> (809) 0:PUGB4, pass, PENB
			8'd38 : rdata = 43'b1100011100001001000000000000000000100000000;
			// PEs: 32 -> 26
			// srcs: (227, 39)(809) 0 --> (809) 0:PUGB4, pass, PEGB2
			8'd39 : rdata = 43'b1100011100001001000000000000000000010100000;
			// PEs: 32 -> 27
			// srcs: (228, 40)(809) 0 --> (809) 0:PUGB4, pass, PEGB3
			8'd40 : rdata = 43'b1100011100001001000000000000000000010110000;
			// PEs: 32 -> 28
			// srcs: (230, 41)(809) 0 --> (809) 0:PUGB4, pass, PEGB4
			8'd41 : rdata = 43'b1100011100001001000000000000000000011000000;
			// PEs: 32 -> 29
			// srcs: (231, 42)(809) 0 --> (809) 0:PUGB4, pass, PEGB5
			8'd42 : rdata = 43'b1100011100001001000000000000000000011010000;
			// PEs: 32 -> 30
			// srcs: (233, 43)(809) 0 --> (809) 0:PUGB4, pass, PEGB6
			8'd43 : rdata = 43'b1100011100001001000000000000000000011100000;
			// PEs: 32 -> 31
			// srcs: (234, 44)(809) 0 --> (809) 0:PUGB4, pass, PEGB7
			8'd44 : rdata = 43'b1100011100001001000000000000000000011110000;
			// PEs: 32 -> 25
			// srcs: (303, 45)(809) 0 --> (809) 0:PUGB4, pass, PENB
			8'd45 : rdata = 43'b1100011100001001000000000000000000100000000;
			// PEs: 32 -> 26
			// srcs: (305, 46)(809) 0 --> (809) 0:PUGB4, pass, PEGB2
			8'd46 : rdata = 43'b1100011100001001000000000000000000010100000;
			// PEs: 32 -> 27
			// srcs: (306, 47)(809) 0 --> (809) 0:PUGB4, pass, PEGB3
			8'd47 : rdata = 43'b1100011100001001000000000000000000010110000;
			// PEs: 32 -> 28
			// srcs: (308, 48)(809) 0 --> (809) 0:PUGB4, pass, PEGB4
			8'd48 : rdata = 43'b1100011100001001000000000000000000011000000;
			// PEs: 32 -> 29
			// srcs: (309, 49)(809) 0 --> (809) 0:PUGB4, pass, PEGB5
			8'd49 : rdata = 43'b1100011100001001000000000000000000011010000;
			// PEs: 32 -> 30
			// srcs: (311, 50)(809) 0 --> (809) 0:PUGB4, pass, PEGB6
			8'd50 : rdata = 43'b1100011100001001000000000000000000011100000;
			// PEs: 32 -> 31
			// srcs: (312, 51)(809) 0 --> (809) 0:PUGB4, pass, PEGB7
			8'd51 : rdata = 43'b1100011100001001000000000000000000011110000;
			// PEs: 32 -> 25
			// srcs: (363, 52)(809) 0 --> (809) 0:PUGB4, pass, PENB
			8'd52 : rdata = 43'b1100011100001001000000000000000000100000000;
			// PEs: 32 -> 26
			// srcs: (366, 53)(809) 0 --> (809) 0:PUGB4, pass, PEGB2
			8'd53 : rdata = 43'b1100011100001001000000000000000000010100000;
			// PEs: 32 -> 27
			// srcs: (369, 54)(809) 0 --> (809) 0:PUGB4, pass, PEGB3
			8'd54 : rdata = 43'b1100011100001001000000000000000000010110000;
			// PEs: 32 -> 28
			// srcs: (372, 55)(809) 0 --> (809) 0:PUGB4, pass, PEGB4
			8'd55 : rdata = 43'b1100011100001001000000000000000000011000000;
			// PEs: 32 -> 29
			// srcs: (379, 56)(809) 0 --> (809) 0:PUGB4, pass, PEGB5
			8'd56 : rdata = 43'b1100011100001001000000000000000000011010000;
			// PEs: 32 -> 25
			// srcs: (381, 57)(809) 0 --> (809) 0:PUGB4, pass, PENB
			8'd57 : rdata = 43'b1100011100001001000000000000000000100000000;
			// PEs: 32 -> 30
			// srcs: (382, 58)(809) 0 --> (809) 0:PUGB4, pass, PEGB6
			8'd58 : rdata = 43'b1100011100001001000000000000000000011100000;
			// PEs: 32 -> 26
			// srcs: (383, 59)(809) 0 --> (809) 0:PUGB4, pass, PEGB2
			8'd59 : rdata = 43'b1100011100001001000000000000000000010100000;
			// PEs: 32 -> 27
			// srcs: (384, 60)(809) 0 --> (809) 0:PUGB4, pass, PEGB3
			8'd60 : rdata = 43'b1100011100001001000000000000000000010110000;
			// PEs: 32 -> 31
			// srcs: (385, 61)(809) 0 --> (809) 0:PUGB4, pass, PEGB7
			8'd61 : rdata = 43'b1100011100001001000000000000000000011110000;
			// PEs: 32 -> 28
			// srcs: (386, 62)(809) 0 --> (809) 0:PUGB4, pass, PEGB4
			8'd62 : rdata = 43'b1100011100001001000000000000000000011000000;
			// PEs: 32 -> 29
			// srcs: (387, 63)(809) 0 --> (809) 0:PUGB4, pass, PEGB5
			8'd63 : rdata = 43'b1100011100001001000000000000000000011010000;
			// PEs: 32 -> 30
			// srcs: (389, 64)(809) 0 --> (809) 0:PUGB4, pass, PEGB6
			8'd64 : rdata = 43'b1100011100001001000000000000000000011100000;
			// PEs: 32 -> 31
			// srcs: (390, 65)(809) 0 --> (809) 0:PUGB4, pass, PEGB7
			8'd65 : rdata = 43'b1100011100001001000000000000000000011110000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 25) begin
	always @(*) begin
		case(address)
			// PEs: 25, 25 -> 25
			// srcs: (1, 0)(32) -1, (233) 2 --> (433) -2:ND0, NW0, *, NI0
			8'd0 : rdata = 43'b0001101100000000010000000001000000000000000;
			// PEs: 25, 25 -> 28
			// srcs: (2, 1)(109) 2, (310) -2 --> (510) -4:ND1, NW1, *, PEGB4
			8'd1 : rdata = 43'b0001101100000001010000000010000000011000000;
			// PEs: 25, 25 -> 25
			// srcs: (3, 2)(187) 2, (388) 0 --> (588) 0:ND2, NW2, *, NI1
			8'd2 : rdata = 43'b0001101100000010010000000101010000000000000;
			// PEs: 25, 25 -> 25
			// srcs: (4, 3)(169) -1, (370) -3 --> (570) 3:ND3, NW3, *, NI2
			8'd3 : rdata = 43'b0001101100000011010000000111100000000000000;
			// PEs: 27 -> 
			// srcs: (6, 4)(435) 2 --> (435) 2:PEGB3, pass, 
			8'd4 : rdata = 43'b1100011100000110000000000000000000000000000;
			// PEs: 26, 25 -> 24
			// srcs: (9, 5)(434) 0, (435) 2 --> (632) 2:PEGB2, ALU, +, PEGB0
			8'd5 : rdata = 43'b0000111100000100001111111110000000010000000;
			// PEs: 24, 25 -> 26
			// srcs: (10, 6)(587) 0, (588) 0 --> (783) 0:PENB, NI1, +, PENB
			8'd6 : rdata = 43'b0000111011111110101000000010000000100000000;
			// PEs: 24, 25 -> 
			// srcs: (19, 7)(432) 0, (433) -2 --> (630) -2:PENB, NI0, +, 
			8'd7 : rdata = 43'b0000111011111110101000000000000000000000000;
			// PEs: 24, 25 -> 24
			// srcs: (29, 8)(629) -1, (630) -2 --> (631) -3:PENB, ALU, +, PEGB0
			8'd8 : rdata = 43'b0000111011111110001111111110000000010000000;
			// PEs: 29, 24 -> 28
			// srcs: (30, 9)(712) 11, (517) 0 --> (713) 11:PEGB5, PENB, +, PEGB4
			8'd9 : rdata = 43'b0000111100001010110111111100000000011000000;
			// PEs: 24 -> 
			// srcs: (31, 10)(526) -2 --> (526) -2:PENB, pass, 
			8'd10 : rdata = 43'b1100011011111110000000000000000000000000000;
			// PEs: 24, 25 -> 24
			// srcs: (36, 11)(721) 8, (526) -2 --> (722) 6:PENB, ALU, +, PEGB0
			8'd11 : rdata = 43'b0000111011111110001111111110000000010000000;
			// PEs: 24, 25 -> 25
			// srcs: (37, 12)(765) -1, (570) 3 --> (766) 2:PENB, NI2, +, NI0
			8'd12 : rdata = 43'b0000111011111110101000000101000000000000000;
			// PEs: 24, 26 -> 26
			// srcs: (38, 13)(767) 6, (573) 0 --> (768) 6:PENB, PEGB2, +, PENB
			8'd13 : rdata = 43'b0000111011111110111000001000000000100000000;
			// PEs: 25 -> 26
			// srcs: (45, 18)(766) 2 --> (766) 2:NI0, pass, PENB
			8'd14 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 24, 28 -> 24
			// srcs: (49, 14)(772) -2, (579) 0 --> (773) -2:PENB, PEGB4, +, PEGB0
			8'd15 : rdata = 43'b0000111011111110111000010000000000010000000;
			// PEs: 24, 29 -> 25
			// srcs: (57, 15)(780) -1, (586) -2 --> (781) -3:PENB, PEGB5, +, NI0
			8'd16 : rdata = 43'b0000111011111110111000010101000000000000000;
			// PEs: 24 -> 
			// srcs: (80, 16)(743) 9 --> (743) 9:PENB, pass, 
			8'd17 : rdata = 43'b1100011011111110000000000000000000000000000;
			// PEs: 24, 25 -> 24
			// srcs: (87, 17)(741) -2, (743) 9 --> (744) 7:PENB, ALU, +, PEGB0
			8'd18 : rdata = 43'b0000111011111110001111111110000000010000000;
			// PEs: 24, 25 -> 29
			// srcs: (88, 19)(779) -1, (781) -3 --> (782) -4:PENB, NI0, +, PEGB5
			8'd19 : rdata = 43'b0000111011111110101000000000000000011010000;
			// PEs: 24 -> 
			// srcs: (120, 20)(701) -2 --> (701) -2:PENB, pass, 
			8'd20 : rdata = 43'b1100011011111110000000000000000000000000000;
			// PEs: 24, 25 -> 
			// srcs: (126, 21)(677) 16, (701) -2 --> (702) 14:PENB, ALU, +, 
			8'd21 : rdata = 43'b0000111011111110001111111110000000000000000;
			// PEs: 24, 25 -> 24
			// srcs: (136, 22)(653) 21, (702) 14 --> (703) 35:PENB, ALU, +, PEGB0
			8'd22 : rdata = 43'b0000111011111110001111111110000000010000000;
			// PEs: 24, 25 -> 26
			// srcs: (228, 23)(809) 0, (32) -1 --> (838) 0:PENB, ND0, *, PENB
			8'd23 : rdata = 43'b0001111011111110011000000000000000100000000;
			// PEs: 25, 26 -> 25
			// srcs: (237, 27)(233) 2, (1038) 0 --> (1238) 2:NW0, PEGB2, -, NW0
			8'd24 : rdata = 43'b0001001000000000111000001000001000000000000;
			// PEs: 24, 25 -> 26
			// srcs: (305, 24)(809) 0, (109) 2 --> (915) 0:PENB, ND1, *, PENB
			8'd25 : rdata = 43'b0001111011111110011000000010000000100000000;
			// PEs: 25, 26 -> 25
			// srcs: (314, 28)(310) -2, (1115) 0 --> (1315) -2:NW1, PEGB2, -, NW1
			8'd26 : rdata = 43'b0001001000000001111000001000001010000000000;
			// PEs: 24, 25 -> 26
			// srcs: (365, 25)(809) 0, (169) -1 --> (975) 0:PENB, ND3, *, PENB
			8'd27 : rdata = 43'b0001111011111110011000000110000000100000000;
			// PEs: 25, 26 -> 25
			// srcs: (374, 29)(370) -3, (1175) 0 --> (1375) -3:NW3, PEGB2, -, NW3
			8'd28 : rdata = 43'b0001001000000011111000001000001110000000000;
			// PEs: 24, 25 -> 26
			// srcs: (383, 26)(809) 0, (187) 2 --> (993) 0:PENB, ND2, *, PENB
			8'd29 : rdata = 43'b0001111011111110011000000100000000100000000;
			// PEs: 25, 26 -> 25
			// srcs: (392, 30)(388) 0, (1193) 0 --> (1393) 0:NW2, PEGB2, -, NW2
			8'd30 : rdata = 43'b0001001000000010111000001000001100000000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 26) begin
	always @(*) begin
		case(address)
			// PEs: 26, 26 -> 25
			// srcs: (1, 0)(33) 0, (234) 0 --> (434) 0:ND0, NW0, *, PEGB1
			8'd0 : rdata = 43'b0001101100000000010000000000000000010010000;
			// PEs: 26, 26 -> 27
			// srcs: (2, 1)(111) 1, (312) -3 --> (512) -3:ND1, NW1, *, PENB
			8'd1 : rdata = 43'b0001101100000001010000000010000000100000000;
			// PEs: 26, 26 -> 30
			// srcs: (3, 2)(189) -1, (390) -3 --> (590) 3:ND2, NW2, *, PEGB6
			8'd2 : rdata = 43'b0001101100000010010000000100000000011100000;
			// PEs: 26, 26 -> 25
			// srcs: (4, 3)(172) 1, (373) 0 --> (573) 0:ND3, NW3, *, PEGB1
			8'd3 : rdata = 43'b0001101100000011010000000110000000010010000;
			// PEs: 29 -> 
			// srcs: (6, 4)(438) 0 --> (438) 0:PEGB5, pass, 
			8'd4 : rdata = 43'b1100011100001010000000000000000000000000000;
			// PEs: 28, 26 -> 24
			// srcs: (9, 5)(437) 4, (438) 0 --> (635) 4:PEGB4, ALU, +, PEGB0
			8'd5 : rdata = 43'b0000111100001000001111111110000000010000000;
			// PEs: 25, 30 -> 30
			// srcs: (16, 6)(783) 0, (589) 0 --> (784) 0:PENB, PEGB6, +, PEGB6
			8'd6 : rdata = 43'b0000111011111110111000011000000000011100000;
			// PEs: 25 -> 
			// srcs: (40, 7)(768) 6 --> (768) 6:PENB, pass, 
			8'd7 : rdata = 43'b1100011011111110000000000000000000000000000;
			// PEs: 25, 26 -> 24
			// srcs: (47, 8)(766) 2, (768) 6 --> (769) 8:PENB, ALU, +, PEGB0
			8'd8 : rdata = 43'b0000111011111110001111111110000000010000000;
			// PEs: 26, 25 -> 25
			// srcs: (231, 13)(3) 1, (838) 0 --> (1038) 0:NM0, PENB, *, PEGB1
			8'd9 : rdata = 43'b0001110000000000110111111100000000010010000;
			// PEs: 24, 26 -> 27
			// srcs: (232, 9)(809) 0, (33) 0 --> (839) 0:PEGB0, ND0, *, PENB
			8'd10 : rdata = 43'b0001111100000000011000000000000000100000000;
			// PEs: 26, 27 -> 26
			// srcs: (241, 18)(234) 0, (1039) 0 --> (1239) 0:NW0, PEGB3, -, NW0
			8'd11 : rdata = 43'b0001001000000000111000001100001000000000000;
			// PEs: 26, 25 -> 25
			// srcs: (308, 14)(3) 1, (915) 0 --> (1115) 0:NM0, PENB, *, PEGB1
			8'd12 : rdata = 43'b0001110000000000110111111100000000010010000;
			// PEs: 24, 26 -> 27
			// srcs: (310, 10)(809) 0, (111) 1 --> (917) 0:PEGB0, ND1, *, PENB
			8'd13 : rdata = 43'b0001111100000000011000000010000000100000000;
			// PEs: 26, 27 -> 26
			// srcs: (319, 19)(312) -3, (1117) 0 --> (1317) -3:NW1, PEGB3, -, NW1
			8'd14 : rdata = 43'b0001001000000001111000001100001010000000000;
			// PEs: 26, 25 -> 25
			// srcs: (368, 15)(3) 1, (975) 0 --> (1175) 0:NM0, PENB, *, PEGB1
			8'd15 : rdata = 43'b0001110000000000110111111100000000010010000;
			// PEs: 24, 26 -> 
			// srcs: (371, 11)(809) 0, (172) 1 --> (978) 0:PEGB0, ND3, *, 
			8'd16 : rdata = 43'b0001111100000000011000000110000000000000000;
			// PEs: 26, 26 -> 
			// srcs: (374, 16)(3) 1, (978) 0 --> (1178) 0:NM0, ALU, *, 
			8'd17 : rdata = 43'b0001110000000000001111111110000000000000000;
			// PEs: 26, 26 -> 26
			// srcs: (377, 20)(373) 0, (1178) 0 --> (1378) 0:NW3, ALU, -, NW3
			8'd18 : rdata = 43'b0001001000000011001111111110001110000000000;
			// PEs: 26, 25 -> 25
			// srcs: (386, 17)(3) 1, (993) 0 --> (1193) 0:NM0, PENB, *, PEGB1
			8'd19 : rdata = 43'b0001110000000000110111111100000000010010000;
			// PEs: 24, 26 -> 27
			// srcs: (388, 12)(809) 0, (189) -1 --> (995) 0:PEGB0, ND2, *, PENB
			8'd20 : rdata = 43'b0001111100000000011000000100000000100000000;
			// PEs: 26, 27 -> 26
			// srcs: (397, 21)(390) -3, (1195) 0 --> (1395) -3:NW2, PEGB3, -, NW2
			8'd21 : rdata = 43'b0001001000000010111000001100001100000000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 27) begin
	always @(*) begin
		case(address)
			// PEs: 27, 27 -> 25
			// srcs: (1, 0)(34) 2, (235) 1 --> (435) 2:ND0, NW0, *, PEGB1
			8'd0 : rdata = 43'b0001101100000000010000000000000000010010000;
			// PEs: 27, 27 -> 27
			// srcs: (2, 1)(112) 2, (313) 2 --> (513) 4:ND1, NW1, *, NI0
			8'd1 : rdata = 43'b0001101100000001010000000011000000000000000;
			// PEs: 27, 27 -> 30
			// srcs: (3, 2)(190) -3, (391) 2 --> (591) -6:ND2, NW2, *, PEGB6
			8'd2 : rdata = 43'b0001101100000010010000000100000000011100000;
			// PEs: 27, 27 -> 27
			// srcs: (4, 3)(175) -1, (376) -1 --> (576) 1:ND3, NW3, *, NI1
			8'd3 : rdata = 43'b0001101100000011010000000111010000000000000;
			// PEs: 26, 27 -> 24
			// srcs: (5, 6)(512) -3, (513) 4 --> (710) 1:PENB, NI0, +, PEGB0
			8'd4 : rdata = 43'b0000111011111110101000000000000000010000000;
			// PEs: 31 -> 
			// srcs: (6, 4)(441) 0 --> (441) 0:PEGB7, pass, 
			8'd5 : rdata = 43'b1100011100001110000000000000000000000000000;
			// PEs: 30, 27 -> 24
			// srcs: (9, 5)(440) 9, (441) 0 --> (637) 9:PEGB6, ALU, +, PEGB0
			8'd6 : rdata = 43'b0000111100001100001111111110000000010000000;
			// PEs: 27 -> 24
			// srcs: (25, 7)(576) 1 --> (576) 1:NI1, pass, PEGB0
			8'd7 : rdata = 43'b1100010100000001000000000000000000010000000;
			// PEs: 24, 27 -> 28
			// srcs: (233, 8)(809) 0, (34) 2 --> (840) 0:PEGB0, ND0, *, PENB
			8'd8 : rdata = 43'b0001111100000000011000000000000000100000000;
			// PEs: 27, 26 -> 26
			// srcs: (235, 12)(3) 1, (839) 0 --> (1039) 0:NM0, PENB, *, PEGB2
			8'd9 : rdata = 43'b0001110000000000110111111100000000010100000;
			// PEs: 27, 28 -> 27
			// srcs: (242, 17)(235) 1, (1040) 0 --> (1240) 1:NW0, PEGB4, -, NW0
			8'd10 : rdata = 43'b0001001000000000111000010000001000000000000;
			// PEs: 24, 27 -> 27
			// srcs: (311, 9)(809) 0, (112) 2 --> (918) 0:PEGB0, ND1, *, NI0
			8'd11 : rdata = 43'b0001111100000000011000000011000000000000000;
			// PEs: 27, 26 -> 26
			// srcs: (313, 13)(3) 1, (917) 0 --> (1117) 0:NM0, PENB, *, PEGB2
			8'd12 : rdata = 43'b0001110000000000110111111100000000010100000;
			// PEs: 27, 27 -> 
			// srcs: (314, 14)(3) 1, (918) 0 --> (1118) 0:NM0, NI0, *, 
			8'd13 : rdata = 43'b0001110000000000101000000000000000000000000;
			// PEs: 27, 27 -> 27
			// srcs: (317, 18)(313) 2, (1118) 0 --> (1318) 2:NW1, ALU, -, NW1
			8'd14 : rdata = 43'b0001001000000001001111111110001010000000000;
			// PEs: 24, 27 -> 
			// srcs: (374, 10)(809) 0, (175) -1 --> (981) 0:PEGB0, ND3, *, 
			8'd15 : rdata = 43'b0001111100000000011000000110000000000000000;
			// PEs: 27, 27 -> 
			// srcs: (377, 15)(3) 1, (981) 0 --> (1181) 0:NM0, ALU, *, 
			8'd16 : rdata = 43'b0001110000000000001111111110000000000000000;
			// PEs: 27, 27 -> 27
			// srcs: (380, 19)(376) -1, (1181) 0 --> (1381) -1:NW3, ALU, -, NW3
			8'd17 : rdata = 43'b0001001000000011001111111110001110000000000;
			// PEs: 24, 27 -> 28
			// srcs: (389, 11)(809) 0, (190) -3 --> (996) 0:PEGB0, ND2, *, PENB
			8'd18 : rdata = 43'b0001111100000000011000000100000000100000000;
			// PEs: 27, 26 -> 26
			// srcs: (391, 16)(3) 1, (995) 0 --> (1195) 0:NM0, PENB, *, PEGB2
			8'd19 : rdata = 43'b0001110000000000110111111100000000010100000;
			// PEs: 27, 28 -> 27
			// srcs: (398, 20)(391) 2, (1196) 0 --> (1396) 2:NW2, PEGB4, -, NW2
			8'd20 : rdata = 43'b0001001000000010111000010000001100000000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 28) begin
	always @(*) begin
		case(address)
			// PEs: 28, 28 -> 26
			// srcs: (1, 0)(36) -2, (237) -2 --> (437) 4:ND0, NW0, *, PEGB2
			8'd0 : rdata = 43'b0001101100000000010000000000000000010100000;
			// PEs: 28, 28 -> 29
			// srcs: (2, 1)(114) -3, (315) -3 --> (515) 9:ND1, NW1, *, PENB
			8'd1 : rdata = 43'b0001101100000001010000000010000000100000000;
			// PEs: 28, 28 -> 29
			// srcs: (3, 2)(192) 1, (393) -2 --> (593) -2:ND2, NW2, *, PENB
			8'd2 : rdata = 43'b0001101100000010010000000100000000100000000;
			// PEs: 28, 28 -> 25
			// srcs: (4, 3)(178) 0, (379) 1 --> (579) 0:ND3, NW3, *, PEGB1
			8'd3 : rdata = 43'b0001101100000011010000000110000000010010000;
			// PEs: 24 -> 
			// srcs: (11, 4)(509) 0 --> (509) 0:PEGB0, pass, 
			8'd4 : rdata = 43'b1100011100000000000000000000000000000000000;
			// PEs: 28, 25 -> 24
			// srcs: (14, 5)(509) 0, (510) -4 --> (707) -4:ALU, PEGB1, +, PEGB0
			8'd5 : rdata = 43'b0000100111111111111000000100000000010000000;
			// PEs: 24 -> 
			// srcs: (54, 6)(711) -3 --> (711) -3:PEGB0, pass, 
			8'd6 : rdata = 43'b1100011100000000000000000000000000000000000;
			// PEs: 28, 25 -> 24
			// srcs: (56, 7)(711) -3, (713) 11 --> (714) 8:ALU, PEGB1, +, PEGB0
			8'd7 : rdata = 43'b0000100111111111111000000100000000010000000;
			// PEs: 24, 28 -> 28
			// srcs: (235, 8)(809) 0, (36) -2 --> (842) 0:PEGB0, ND0, *, NI0
			8'd8 : rdata = 43'b0001111100000000011000000001000000000000000;
			// PEs: 28, 27 -> 27
			// srcs: (236, 12)(3) 1, (840) 0 --> (1040) 0:NM0, PENB, *, PEGB3
			8'd9 : rdata = 43'b0001110000000000110111111100000000010110000;
			// PEs: 28, 28 -> 
			// srcs: (238, 13)(3) 1, (842) 0 --> (1042) 0:NM0, NI0, *, 
			8'd10 : rdata = 43'b0001110000000000101000000000000000000000000;
			// PEs: 28, 28 -> 28
			// srcs: (241, 16)(237) -2, (1042) 0 --> (1242) -2:NW0, ALU, -, NW0
			8'd11 : rdata = 43'b0001001000000000001111111110001000000000000;
			// PEs: 24, 28 -> 29
			// srcs: (313, 9)(809) 0, (114) -3 --> (920) 0:PEGB0, ND1, *, PENB
			8'd12 : rdata = 43'b0001111100000000011000000010000000100000000;
			// PEs: 28, 29 -> 28
			// srcs: (322, 17)(315) -3, (1120) 0 --> (1320) -3:NW1, PEGB5, -, NW1
			8'd13 : rdata = 43'b0001001000000001111000010100001010000000000;
			// PEs: 24, 28 -> 
			// srcs: (377, 10)(809) 0, (178) 0 --> (984) 0:PEGB0, ND3, *, 
			8'd14 : rdata = 43'b0001111100000000011000000110000000000000000;
			// PEs: 28, 28 -> 
			// srcs: (380, 14)(3) 1, (984) 0 --> (1184) 0:NM0, ALU, *, 
			8'd15 : rdata = 43'b0001110000000000001111111110000000000000000;
			// PEs: 28, 28 -> 28
			// srcs: (383, 18)(379) 1, (1184) 0 --> (1384) 1:NW3, ALU, -, NW3
			8'd16 : rdata = 43'b0001001000000011001111111110001110000000000;
			// PEs: 24, 28 -> 29
			// srcs: (391, 11)(809) 0, (192) 1 --> (998) 0:PEGB0, ND2, *, PENB
			8'd17 : rdata = 43'b0001111100000000011000000100000000100000000;
			// PEs: 28, 27 -> 27
			// srcs: (392, 15)(3) 1, (996) 0 --> (1196) 0:NM0, PENB, *, PEGB3
			8'd18 : rdata = 43'b0001110000000000110111111100000000010110000;
			// PEs: 28, 29 -> 28
			// srcs: (400, 19)(393) -2, (1198) 0 --> (1398) -2:NW2, PEGB5, -, NW2
			8'd19 : rdata = 43'b0001001000000010111000010100001100000000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 29) begin
	always @(*) begin
		case(address)
			// PEs: 29, 29 -> 26
			// srcs: (1, 0)(37) 0, (238) 0 --> (438) 0:ND0, NW0, *, PEGB2
			8'd0 : rdata = 43'b0001101100000000010000000000000000010100000;
			// PEs: 29, 29 -> 29
			// srcs: (2, 1)(115) -1, (316) -2 --> (516) 2:ND1, NW1, *, NI0
			8'd1 : rdata = 43'b0001101100000001010000000011000000000000000;
			// PEs: 29, 29 -> 29
			// srcs: (3, 2)(193) 2, (394) -1 --> (594) -2:ND2, NW2, *, NI1
			8'd2 : rdata = 43'b0001101100000010010000000101010000000000000;
			// PEs: 29, 29 -> 29
			// srcs: (4, 3)(185) 1, (386) -2 --> (586) -2:ND3, NW3, *, NI2
			8'd3 : rdata = 43'b0001101100000011010000000111100000000000000;
			// PEs: 28, 29 -> 25
			// srcs: (5, 4)(515) 9, (516) 2 --> (712) 11:PENB, NI0, +, PEGB1
			8'd4 : rdata = 43'b0000111011111110101000000000000000010010000;
			// PEs: 28, 29 -> 24
			// srcs: (6, 5)(593) -2, (594) -2 --> (789) -4:PENB, NI1, +, PEGB0
			8'd5 : rdata = 43'b0000111011111110101000000010000000010000000;
			// PEs: 29 -> 25
			// srcs: (52, 6)(586) -2 --> (586) -2:NI2, pass, PEGB1
			8'd6 : rdata = 43'b1100010100000010000000000000000000010010000;
			// PEs: 25 -> 
			// srcs: (93, 7)(782) -4 --> (782) -4:PEGB1, pass, 
			8'd7 : rdata = 43'b1100011100000010000000000000000000000000000;
			// PEs: 29, 30 -> 24
			// srcs: (96, 8)(782) -4, (787) -9 --> (788) -13:ALU, PEGB6, +, PEGB0
			8'd8 : rdata = 43'b0000100111111111111000011000000000010000000;
			// PEs: 24, 29 -> 30
			// srcs: (236, 9)(809) 0, (37) 0 --> (843) 0:PEGB0, ND0, *, PENB
			8'd9 : rdata = 43'b0001111100000000011000000000000000100000000;
			// PEs: 29, 30 -> 29
			// srcs: (245, 16)(238) 0, (1043) 0 --> (1243) 0:NW0, PEGB6, -, NW0
			8'd10 : rdata = 43'b0001001000000000111000011000001000000000000;
			// PEs: 24, 29 -> 30
			// srcs: (314, 10)(809) 0, (115) -1 --> (921) 0:PEGB0, ND1, *, PENB
			8'd11 : rdata = 43'b0001111100000000011000000010000000100000000;
			// PEs: 29, 28 -> 28
			// srcs: (316, 13)(3) 1, (920) 0 --> (1120) 0:NM0, PENB, *, PEGB4
			8'd12 : rdata = 43'b0001110000000000110111111100000000011000000;
			// PEs: 29, 30 -> 29
			// srcs: (323, 17)(316) -2, (1121) 0 --> (1321) -2:NW1, PEGB6, -, NW1
			8'd13 : rdata = 43'b0001001000000001111000011000001010000000000;
			// PEs: 24, 29 -> 
			// srcs: (384, 11)(809) 0, (185) 1 --> (991) 0:PEGB0, ND3, *, 
			8'd14 : rdata = 43'b0001111100000000011000000110000000000000000;
			// PEs: 29, 29 -> 
			// srcs: (387, 14)(3) 1, (991) 0 --> (1191) 0:NM0, ALU, *, 
			8'd15 : rdata = 43'b0001110000000000001111111110000000000000000;
			// PEs: 29, 29 -> 29
			// srcs: (390, 18)(386) -2, (1191) 0 --> (1391) -2:NW3, ALU, -, NW3
			8'd16 : rdata = 43'b0001001000000011001111111110001110000000000;
			// PEs: 24, 29 -> 30
			// srcs: (392, 12)(809) 0, (193) 2 --> (999) 0:PEGB0, ND2, *, PENB
			8'd17 : rdata = 43'b0001111100000000011000000100000000100000000;
			// PEs: 29, 28 -> 28
			// srcs: (394, 15)(3) 1, (998) 0 --> (1198) 0:NM0, PENB, *, PEGB4
			8'd18 : rdata = 43'b0001110000000000110111111100000000011000000;
			// PEs: 29, 30 -> 29
			// srcs: (401, 19)(394) -1, (1199) 0 --> (1399) -1:NW2, PEGB6, -, NW2
			8'd19 : rdata = 43'b0001001000000010111000011000001100000000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 30) begin
	always @(*) begin
		case(address)
			// PEs: 30, 30 -> 27
			// srcs: (1, 0)(39) -3, (240) -3 --> (440) 9:ND0, NW0, *, PEGB3
			8'd0 : rdata = 43'b0001101100000000010000000000000000010110000;
			// PEs: 30, 30 -> 31
			// srcs: (2, 1)(117) -2, (318) -3 --> (518) 6:ND1, NW1, *, PENB
			8'd1 : rdata = 43'b0001101100000001010000000010000000100000000;
			// PEs: 30, 30 -> 31
			// srcs: (3, 2)(195) -3, (396) -1 --> (596) 3:ND2, NW2, *, PENB
			8'd2 : rdata = 43'b0001101100000010010000000100000000100000000;
			// PEs: 30, 30 -> 26
			// srcs: (4, 3)(188) 0, (389) 2 --> (589) 0:ND3, NW3, *, PEGB2
			8'd3 : rdata = 43'b0001101100000011010000000110000000010100000;
			// PEs: 27 -> 
			// srcs: (8, 4)(591) -6 --> (591) -6:PEGB3, pass, 
			8'd4 : rdata = 43'b1100011100000110000000000000000000000000000;
			// PEs: 26, 30 -> 31
			// srcs: (11, 5)(590) 3, (591) -6 --> (785) -3:PEGB2, ALU, +, PENB
			8'd5 : rdata = 43'b0000111100000100001111111110000000100000000;
			// PEs: 26 -> 
			// srcs: (21, 6)(784) 0 --> (784) 0:PEGB2, pass, 
			8'd6 : rdata = 43'b1100011100000100000000000000000000000000000;
			// PEs: 30, 31 -> 29
			// srcs: (24, 7)(784) 0, (786) -9 --> (787) -9:ALU, PEGB7, +, PEGB5
			8'd7 : rdata = 43'b0000100111111111111000011100000000011010000;
			// PEs: 24, 30 -> 31
			// srcs: (238, 8)(809) 0, (39) -3 --> (845) 0:PEGB0, ND0, *, PENB
			8'd8 : rdata = 43'b0001111100000000011000000000000000100000000;
			// PEs: 30, 29 -> 29
			// srcs: (239, 12)(3) 1, (843) 0 --> (1043) 0:NM0, PENB, *, PEGB5
			8'd9 : rdata = 43'b0001110000000000110111111100000000011010000;
			// PEs: 30, 31 -> 30
			// srcs: (247, 17)(240) -3, (1045) 0 --> (1245) -3:NW0, PEGB7, -, NW0
			8'd10 : rdata = 43'b0001001000000000111000011100001000000000000;
			// PEs: 24, 30 -> 31
			// srcs: (316, 9)(809) 0, (117) -2 --> (923) 0:PEGB0, ND1, *, PENB
			8'd11 : rdata = 43'b0001111100000000011000000010000000100000000;
			// PEs: 30, 29 -> 29
			// srcs: (317, 13)(3) 1, (921) 0 --> (1121) 0:NM0, PENB, *, PEGB5
			8'd12 : rdata = 43'b0001110000000000110111111100000000011010000;
			// PEs: 30, 31 -> 30
			// srcs: (325, 18)(318) -3, (1123) 0 --> (1323) -3:NW1, PEGB7, -, NW1
			8'd13 : rdata = 43'b0001001000000001111000011100001010000000000;
			// PEs: 24, 30 -> 
			// srcs: (387, 10)(809) 0, (188) 0 --> (994) 0:PEGB0, ND3, *, 
			8'd14 : rdata = 43'b0001111100000000011000000110000000000000000;
			// PEs: 30, 30 -> 
			// srcs: (390, 14)(3) 1, (994) 0 --> (1194) 0:NM0, ALU, *, 
			8'd15 : rdata = 43'b0001110000000000001111111110000000000000000;
			// PEs: 30, 30 -> 30
			// srcs: (393, 19)(389) 2, (1194) 0 --> (1394) 2:NW3, ALU, -, NW3
			8'd16 : rdata = 43'b0001001000000011001111111110001110000000000;
			// PEs: 24, 30 -> 30
			// srcs: (394, 11)(809) 0, (195) -3 --> (1001) 0:PEGB0, ND2, *, NI0
			8'd17 : rdata = 43'b0001111100000000011000000101000000000000000;
			// PEs: 30, 29 -> 29
			// srcs: (395, 15)(3) 1, (999) 0 --> (1199) 0:NM0, PENB, *, PEGB5
			8'd18 : rdata = 43'b0001110000000000110111111100000000011010000;
			// PEs: 30, 30 -> 
			// srcs: (397, 16)(3) 1, (1001) 0 --> (1201) 0:NM0, NI0, *, 
			8'd19 : rdata = 43'b0001110000000000101000000000000000000000000;
			// PEs: 30, 30 -> 30
			// srcs: (400, 20)(396) -1, (1201) 0 --> (1401) -1:NW2, ALU, -, NW2
			8'd20 : rdata = 43'b0001001000000010001111111110001100000000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 31) begin
	always @(*) begin
		case(address)
			// PEs: 31, 31 -> 27
			// srcs: (1, 0)(40) 2, (241) 0 --> (441) 0:ND0, NW0, *, PEGB3
			8'd0 : rdata = 43'b0001101100000000010000000000000000010110000;
			// PEs: 31, 31 -> 31
			// srcs: (2, 1)(118) -1, (319) -1 --> (519) 1:ND1, NW1, *, NI0
			8'd1 : rdata = 43'b0001101100000001010000000011000000000000000;
			// PEs: 31, 31 -> 31
			// srcs: (3, 2)(196) 1, (397) 0 --> (597) 0:ND2, NW2, *, NI1
			8'd2 : rdata = 43'b0001101100000010010000000101010000000000000;
			// PEs: 31, 31 -> 31
			// srcs: (4, 3)(191) 2, (392) -3 --> (592) -6:ND3, NW3, *, NI2
			8'd3 : rdata = 43'b0001101100000011010000000111100000000000000;
			// PEs: 30, 31 -> 24
			// srcs: (5, 4)(518) 6, (519) 1 --> (716) 7:PENB, NI0, +, PENB
			8'd4 : rdata = 43'b0000111011111110101000000000000000100000000;
			// PEs: 30, 31 -> 24
			// srcs: (6, 5)(596) 3, (597) 0 --> (791) 3:PENB, NI1, +, PENB
			8'd5 : rdata = 43'b0000111011111110101000000010000000100000000;
			// PEs: 30, 31 -> 30
			// srcs: (14, 6)(785) -3, (592) -6 --> (786) -9:PENB, NI2, +, PEGB6
			8'd6 : rdata = 43'b0000111011111110101000000100000000011100000;
			// PEs: 24, 31 -> 31
			// srcs: (239, 7)(809) 0, (40) 2 --> (846) 0:PEGB0, ND0, *, NI0
			8'd7 : rdata = 43'b0001111100000000011000000001000000000000000;
			// PEs: 31, 30 -> 30
			// srcs: (241, 11)(3) 1, (845) 0 --> (1045) 0:NM0, PENB, *, PEGB6
			8'd8 : rdata = 43'b0001110000000000110111111100000000011100000;
			// PEs: 31, 31 -> 
			// srcs: (242, 12)(3) 1, (846) 0 --> (1046) 0:NM0, NI0, *, 
			8'd9 : rdata = 43'b0001110000000000101000000000000000000000000;
			// PEs: 31, 31 -> 31
			// srcs: (245, 17)(241) 0, (1046) 0 --> (1246) 0:NW0, ALU, -, NW0
			8'd10 : rdata = 43'b0001001000000000001111111110001000000000000;
			// PEs: 24, 31 -> 31
			// srcs: (317, 8)(809) 0, (118) -1 --> (924) 0:PEGB0, ND1, *, NI0
			8'd11 : rdata = 43'b0001111100000000011000000011000000000000000;
			// PEs: 31, 30 -> 30
			// srcs: (319, 13)(3) 1, (923) 0 --> (1123) 0:NM0, PENB, *, PEGB6
			8'd12 : rdata = 43'b0001110000000000110111111100000000011100000;
			// PEs: 31, 31 -> 
			// srcs: (320, 14)(3) 1, (924) 0 --> (1124) 0:NM0, NI0, *, 
			8'd13 : rdata = 43'b0001110000000000101000000000000000000000000;
			// PEs: 31, 31 -> 31
			// srcs: (323, 18)(319) -1, (1124) 0 --> (1324) -1:NW1, ALU, -, NW1
			8'd14 : rdata = 43'b0001001000000001001111111110001010000000000;
			// PEs: 24, 31 -> 
			// srcs: (390, 9)(809) 0, (191) 2 --> (997) 0:PEGB0, ND3, *, 
			8'd15 : rdata = 43'b0001111100000000011000000110000000000000000;
			// PEs: 31, 31 -> 31
			// srcs: (393, 15)(3) 1, (997) 0 --> (1197) 0:NM0, ALU, *, NI0
			8'd16 : rdata = 43'b0001110000000000001111111111000000000000000;
			// PEs: 24, 31 -> 31
			// srcs: (395, 10)(809) 0, (196) 1 --> (1002) 0:PEGB0, ND2, *, NI1
			8'd17 : rdata = 43'b0001111100000000011000000101010000000000000;
			// PEs: 31, 31 -> 31
			// srcs: (396, 19)(392) -3, (1197) 0 --> (1397) -3:NW3, NI0, -, NW3
			8'd18 : rdata = 43'b0001001000000011101000000000001110000000000;
			// PEs: 31, 31 -> 
			// srcs: (398, 16)(3) 1, (1002) 0 --> (1202) 0:NM0, NI1, *, 
			8'd19 : rdata = 43'b0001110000000000101000000010000000000000000;
			// PEs: 31, 31 -> 31
			// srcs: (401, 20)(397) 0, (1202) 0 --> (1402) 0:NW2, ALU, -, NW2
			8'd20 : rdata = 43'b0001001000000010001111111110001100000000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 32) begin
	always @(*) begin
		case(address)
			// PEs: 39 -> 40
			// srcs: (3, 0)(452) -4 --> (452) -4:PENB, pass, PUNB
			8'd0 : rdata = 43'b1100011011111110000000000000000001000000000;
			// PEs: 39 -> 40
			// srcs: (4, 1)(530) 1 --> (530) 1:PENB, pass, PUNB
			8'd1 : rdata = 43'b1100011011111110000000000000000001000000000;
			// PEs: 39 -> 16
			// srcs: (5, 4)(417) -6 --> (417) -6:PENB, pass, PUGB2
			8'd2 : rdata = 43'b1100011011111110000000000000000000000001010;
			// PEs: 37 -> 48
			// srcs: (8, 2)(411) 6 --> (411) 6:PEGB5, pass, PUGB6
			8'd3 : rdata = 43'b1100011100001010000000000000000000000001110;
			// PEs: 38 -> 40
			// srcs: (9, 13)(646) -5 --> (646) -5:PEGB6, pass, PUNB
			8'd4 : rdata = 43'b1100011100001100000000000000000001000000000;
			// PEs: 36 -> 24
			// srcs: (10, 15)(721) 8 --> (721) 8:PEGB4, pass, PUGB3
			8'd5 : rdata = 43'b1100011100001000000000000000000000000001011;
			// PEs: 39 -> 48
			// srcs: (11, 12)(643) 4 --> (643) 4:PENB, pass, PUGB6
			8'd6 : rdata = 43'b1100011011111110000000000000000000000001110;
			// PEs: 38 -> 16
			// srcs: (14, 11)(641) 8 --> (641) 8:PEGB6, pass, PUGB2
			8'd7 : rdata = 43'b1100011100001100000000000000000000000001010;
			// PEs: 8 -> 33
			// srcs: (18, 3)(611) -3 --> (611) -3:PUGB1, pass, PENB
			8'd8 : rdata = 43'b1100011100000011000000000000000000100000000;
			// PEs: 8 -> 32
			// srcs: (19, 5)(617) -1 --> (617) -1:PUGB1, pass, NI0
			8'd9 : rdata = 43'b1100011100000011000000000001000000000000000;
			// PEs: 40 -> 33
			// srcs: (20, 6)(420) 3 --> (420) 3:PUGB5, pass, PENB
			8'd10 : rdata = 43'b1100011100001011000000000000000000100000000;
			// PEs: 32 -> 33
			// srcs: (26, 7)(617) -1 --> (617) -1:NI0, pass, PENB
			8'd11 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 24 -> 32
			// srcs: (27, 8)(637) 9 --> (637) 9:PUNB, pass, NI0
			8'd12 : rdata = 43'b1100011011111111000000000001000000000000000;
			// PEs: 40 -> 33
			// srcs: (28, 9)(442) 0 --> (442) 0:PUGB5, pass, PENB
			8'd13 : rdata = 43'b1100011100001011000000000000000000100000000;
			// PEs: 33 -> 40
			// srcs: (29, 25)(612) -3 --> (612) -3:PEGB1, pass, PUNB
			8'd14 : rdata = 43'b1100011100000010000000000000000001000000000;
			// PEs: 33 -> 40
			// srcs: (33, 26)(618) 2 --> (618) 2:PEGB1, pass, PUNB
			8'd15 : rdata = 43'b1100011100000010000000000000000001000000000;
			// PEs: 32 -> 33
			// srcs: (34, 10)(637) 9 --> (637) 9:NI0, pass, PENB
			8'd16 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 8 -> 33
			// srcs: (41, 14)(523) 6 --> (523) 6:PUGB1, pass, PENB
			8'd17 : rdata = 43'b1100011100000011000000000000000000100000000;
			// PEs: 33 -> 8
			// srcs: (42, 27)(638) 9 --> (638) 9:PEGB1, pass, PUGB1
			8'd18 : rdata = 43'b1100011100000010000000000000000000000001001;
			// PEs: 33 -> 40
			// srcs: (48, 28)(719) 5 --> (719) 5:PEGB1, pass, PUNB
			8'd19 : rdata = 43'b1100011100000010000000000000000001000000000;
			// PEs: 8 -> 33
			// srcs: (58, 16)(529) -6 --> (529) -6:PUGB1, pass, PENB
			8'd20 : rdata = 43'b1100011100000011000000000000000000100000000;
			// PEs: 48 -> 32
			// srcs: (59, 17)(742) 9 --> (742) 9:PUGB6, pass, NI0
			8'd21 : rdata = 43'b1100011100001101000000000001000000000000000;
			// PEs: 16 -> 33
			// srcs: (60, 18)(548) 0 --> (548) 0:PUGB2, pass, PENB
			8'd22 : rdata = 43'b1100011100000101000000000000000000100000000;
			// PEs: 32 -> 33
			// srcs: (66, 19)(742) 9 --> (742) 9:NI0, pass, PENB
			8'd23 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 8 -> 32
			// srcs: (67, 20)(770) 0 --> (770) 0:PUGB1, pass, NI0
			8'd24 : rdata = 43'b1100011100000011000000000001000000000000000;
			// PEs: 24 -> 33
			// srcs: (68, 21)(576) 1 --> (576) 1:PUNB, pass, PENB
			8'd25 : rdata = 43'b1100011011111111000000000000000000100000000;
			// PEs: 33 -> 24
			// srcs: (73, 30)(743) 9 --> (743) 9:PEGB1, pass, PUGB3
			8'd26 : rdata = 43'b1100011100000010000000000000000000000001011;
			// PEs: 32 -> 33
			// srcs: (74, 22)(770) 0 --> (770) 0:NI0, pass, PENB
			8'd27 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 24 -> 33
			// srcs: (75, 23)(789) -4 --> (789) -4:PUNB, pass, PENB
			8'd28 : rdata = 43'b1100011011111111000000000000000000100000000;
			// PEs: 24 -> 33
			// srcs: (76, 24)(791) 3 --> (791) 3:PUNB, pass, PENB
			8'd29 : rdata = 43'b1100011011111111000000000000000000100000000;
			// PEs: 24 -> 35
			// srcs: (77, 29)(722) 6 --> (722) 6:PUNB, pass, PEGB3
			8'd30 : rdata = 43'b1100011011111111000000000000000000010110000;
			// PEs: 24 -> 33
			// srcs: (78, 31)(773) -2 --> (773) -2:PUNB, pass, PENB
			8'd31 : rdata = 43'b1100011011111111000000000000000000100000000;
			// PEs: 24 -> 33
			// srcs: (79, 33)(769) 8 --> (769) 8:PUNB, pass, PENB
			8'd32 : rdata = 43'b1100011011111111000000000000000000100000000;
			// PEs: 35 -> 40
			// srcs: (89, 32)(725) 3 --> (725) 3:PEGB3, pass, PUNB
			8'd33 : rdata = 43'b1100011100000110000000000000000001000000000;
			// PEs: 33 -> 0
			// srcs: (101, 34)(775) 7 --> (775) 7:PEGB1, pass, PUGB0
			8'd34 : rdata = 43'b1100011100000010000000000000000000000001000;
			// PEs: 24 -> 33
			// srcs: (103, 35)(788) -13 --> (788) -13:PUNB, pass, PENB
			8'd35 : rdata = 43'b1100011011111111000000000000000000100000000;
			// PEs: 33 -> 48
			// srcs: (117, 36)(800) -20 --> (800) -20:PEGB1, pass, PUGB6
			8'd36 : rdata = 43'b1100011100000010000000000000000000000001110;
			// PEs: 0 -> 37
			// srcs: (170, 37)(803) 92 --> (803) 92:PUGB0, pass, PEGB5
			8'd37 : rdata = 43'b1100011100000001000000000000000000011010000;
			// PEs: 38 -> 0
			// srcs: (191, 38)(809) 0 --> (809) 0:PEGB6, pass, PUGB0
			8'd38 : rdata = 43'b1100011100001100000000000000000000000001000;
			// PEs: 38 -> 0
			// srcs: (195, 39)(809) 0 --> (809) 0:PEGB6, pass, PUGB0
			8'd39 : rdata = 43'b1100011100001100000000000000000000000001000;
			// PEs: 38 -> 0
			// srcs: (196, 40)(809) 0 --> (809) 0:PEGB6, pass, PUGB0
			8'd40 : rdata = 43'b1100011100001100000000000000000000000001000;
			// PEs: 38 -> 0
			// srcs: (197, 41)(809) 0 --> (809) 0:PEGB6, pass, PUGB0
			8'd41 : rdata = 43'b1100011100001100000000000000000000000001000;
			// PEs: 38 -> 0
			// srcs: (198, 42)(809) 0 --> (809) 0:PEGB6, pass, PUGB0
			8'd42 : rdata = 43'b1100011100001100000000000000000000000001000;
			// PEs: 38 -> 0
			// srcs: (199, 43)(809) 0 --> (809) 0:PEGB6, pass, PUGB0
			8'd43 : rdata = 43'b1100011100001100000000000000000000000001000;
			// PEs: 38 -> 0
			// srcs: (201, 44)(809) 0 --> (809) 0:PEGB6, pass, PUGB0
			8'd44 : rdata = 43'b1100011100001100000000000000000000000001000;
			// PEs: 38 -> 8
			// srcs: (202, 45)(809) 0 --> (809) 0:PEGB6, pass, PUGB1
			8'd45 : rdata = 43'b1100011100001100000000000000000000000001001;
			// PEs: 38 -> 8
			// srcs: (204, 46)(809) 0 --> (809) 0:PEGB6, pass, PUGB1
			8'd46 : rdata = 43'b1100011100001100000000000000000000000001001;
			// PEs: 38 -> 8
			// srcs: (205, 47)(809) 0 --> (809) 0:PEGB6, pass, PUGB1
			8'd47 : rdata = 43'b1100011100001100000000000000000000000001001;
			// PEs: 38 -> 8
			// srcs: (206, 48)(809) 0 --> (809) 0:PEGB6, pass, PUGB1
			8'd48 : rdata = 43'b1100011100001100000000000000000000000001001;
			// PEs: 38 -> 8
			// srcs: (207, 49)(809) 0 --> (809) 0:PEGB6, pass, PUGB1
			8'd49 : rdata = 43'b1100011100001100000000000000000000000001001;
			// PEs: 38 -> 40
			// srcs: (208, 50)(809) 0 --> (809) 0:PEGB6, pass, PUNB
			8'd50 : rdata = 43'b1100011100001100000000000000000001000000000;
			// PEs: 38 -> 8
			// srcs: (209, 51)(809) 0 --> (809) 0:PEGB6, pass, PUGB1
			8'd51 : rdata = 43'b1100011100001100000000000000000000000001001;
			// PEs: 38 -> 8
			// srcs: (210, 52)(809) 0 --> (809) 0:PEGB6, pass, PUGB1
			8'd52 : rdata = 43'b1100011100001100000000000000000000000001001;
			// PEs: 38 -> 40
			// srcs: (211, 53)(809) 0 --> (809) 0:PEGB6, pass, PUNB
			8'd53 : rdata = 43'b1100011100001100000000000000000001000000000;
			// PEs: 38 -> 16
			// srcs: (212, 54)(809) 0 --> (809) 0:PEGB6, pass, PUGB2
			8'd54 : rdata = 43'b1100011100001100000000000000000000000001010;
			// PEs: 38 -> 16
			// srcs: (213, 55)(809) 0 --> (809) 0:PEGB6, pass, PUGB2
			8'd55 : rdata = 43'b1100011100001100000000000000000000000001010;
			// PEs: 38 -> 40
			// srcs: (214, 56)(809) 0 --> (809) 0:PEGB6, pass, PUNB
			8'd56 : rdata = 43'b1100011100001100000000000000000001000000000;
			// PEs: 38 -> 16
			// srcs: (215, 57)(809) 0 --> (809) 0:PEGB6, pass, PUGB2
			8'd57 : rdata = 43'b1100011100001100000000000000000000000001010;
			// PEs: 38 -> 16
			// srcs: (216, 58)(809) 0 --> (809) 0:PEGB6, pass, PUGB2
			8'd58 : rdata = 43'b1100011100001100000000000000000000000001010;
			// PEs: 38 -> 40
			// srcs: (217, 59)(809) 0 --> (809) 0:PEGB6, pass, PUNB
			8'd59 : rdata = 43'b1100011100001100000000000000000001000000000;
			// PEs: 38 -> 16
			// srcs: (218, 60)(809) 0 --> (809) 0:PEGB6, pass, PUGB2
			8'd60 : rdata = 43'b1100011100001100000000000000000000000001010;
			// PEs: 38 -> 16
			// srcs: (219, 61)(809) 0 --> (809) 0:PEGB6, pass, PUGB2
			8'd61 : rdata = 43'b1100011100001100000000000000000000000001010;
			// PEs: 38 -> 16
			// srcs: (220, 62)(809) 0 --> (809) 0:PEGB6, pass, PUGB2
			8'd62 : rdata = 43'b1100011100001100000000000000000000000001010;
			// PEs: 38 -> 24
			// srcs: (221, 63)(809) 0 --> (809) 0:PEGB6, pass, PUGB3
			8'd63 : rdata = 43'b1100011100001100000000000000000000000001011;
			// PEs: 38 -> 24
			// srcs: (222, 64)(809) 0 --> (809) 0:PEGB6, pass, PUGB3
			8'd64 : rdata = 43'b1100011100001100000000000000000000000001011;
			// PEs: 38 -> 24
			// srcs: (223, 65)(809) 0 --> (809) 0:PEGB6, pass, PUGB3
			8'd65 : rdata = 43'b1100011100001100000000000000000000000001011;
			// PEs: 38 -> 40
			// srcs: (224, 66)(809) 0 --> (809) 0:PEGB6, pass, PUNB
			8'd66 : rdata = 43'b1100011100001100000000000000000001000000000;
			// PEs: 38 -> 24
			// srcs: (225, 67)(809) 0 --> (809) 0:PEGB6, pass, PUGB3
			8'd67 : rdata = 43'b1100011100001100000000000000000000000001011;
			// PEs: 38 -> 24
			// srcs: (226, 68)(809) 0 --> (809) 0:PEGB6, pass, PUGB3
			8'd68 : rdata = 43'b1100011100001100000000000000000000000001011;
			// PEs: 38 -> 40
			// srcs: (227, 69)(809) 0 --> (809) 0:PEGB6, pass, PUNB
			8'd69 : rdata = 43'b1100011100001100000000000000000001000000000;
			// PEs: 38 -> 24
			// srcs: (228, 70)(809) 0 --> (809) 0:PEGB6, pass, PUGB3
			8'd70 : rdata = 43'b1100011100001100000000000000000000000001011;
			// PEs: 38 -> 24
			// srcs: (229, 71)(809) 0 --> (809) 0:PEGB6, pass, PUGB3
			8'd71 : rdata = 43'b1100011100001100000000000000000000000001011;
			// PEs: 38 -> 40
			// srcs: (230, 72)(809) 0 --> (809) 0:PEGB6, pass, PUNB
			8'd72 : rdata = 43'b1100011100001100000000000000000001000000000;
			// PEs: 38 -> 48
			// srcs: (233, 73)(809) 0 --> (809) 0:PEGB6, pass, PUGB6
			8'd73 : rdata = 43'b1100011100001100000000000000000000000001110;
			// PEs: 38 -> 48
			// srcs: (236, 74)(809) 0 --> (809) 0:PEGB6, pass, PUGB6
			8'd74 : rdata = 43'b1100011100001100000000000000000000000001110;
			// PEs: 38 -> 48
			// srcs: (239, 75)(809) 0 --> (809) 0:PEGB6, pass, PUGB6
			8'd75 : rdata = 43'b1100011100001100000000000000000000000001110;
			// PEs: 38 -> 40
			// srcs: (241, 76)(809) 0 --> (809) 0:PEGB6, pass, PUNB
			8'd76 : rdata = 43'b1100011100001100000000000000000001000000000;
			// PEs: 38 -> 48
			// srcs: (242, 77)(809) 0 --> (809) 0:PEGB6, pass, PUGB6
			8'd77 : rdata = 43'b1100011100001100000000000000000000000001110;
			// PEs: 38 -> 40
			// srcs: (243, 78)(809) 0 --> (809) 0:PEGB6, pass, PUNB
			8'd78 : rdata = 43'b1100011100001100000000000000000001000000000;
			// PEs: 38 -> 40
			// srcs: (244, 79)(809) 0 --> (809) 0:PEGB6, pass, PUNB
			8'd79 : rdata = 43'b1100011100001100000000000000000001000000000;
			// PEs: 38 -> 40
			// srcs: (245, 80)(809) 0 --> (809) 0:PEGB6, pass, PUNB
			8'd80 : rdata = 43'b1100011100001100000000000000000001000000000;
			// PEs: 38 -> 40
			// srcs: (246, 81)(809) 0 --> (809) 0:PEGB6, pass, PUNB
			8'd81 : rdata = 43'b1100011100001100000000000000000001000000000;
			// PEs: 38 -> 40
			// srcs: (247, 82)(809) 0 --> (809) 0:PEGB6, pass, PUNB
			8'd82 : rdata = 43'b1100011100001100000000000000000001000000000;
			// PEs: 38 -> 40
			// srcs: (248, 83)(809) 0 --> (809) 0:PEGB6, pass, PUNB
			8'd83 : rdata = 43'b1100011100001100000000000000000001000000000;
			// PEs: 38 -> 48
			// srcs: (249, 84)(809) 0 --> (809) 0:PEGB6, pass, PUGB6
			8'd84 : rdata = 43'b1100011100001100000000000000000000000001110;
			// PEs: 38 -> 48
			// srcs: (250, 85)(809) 0 --> (809) 0:PEGB6, pass, PUGB6
			8'd85 : rdata = 43'b1100011100001100000000000000000000000001110;
			// PEs: 38 -> 48
			// srcs: (251, 86)(809) 0 --> (809) 0:PEGB6, pass, PUGB6
			8'd86 : rdata = 43'b1100011100001100000000000000000000000001110;
			// PEs: 38 -> 48
			// srcs: (252, 87)(809) 0 --> (809) 0:PEGB6, pass, PUGB6
			8'd87 : rdata = 43'b1100011100001100000000000000000000000001110;
			// PEs: 38 -> 48
			// srcs: (253, 88)(809) 0 --> (809) 0:PEGB6, pass, PUGB6
			8'd88 : rdata = 43'b1100011100001100000000000000000000000001110;
			// PEs: 38 -> 48
			// srcs: (254, 89)(809) 0 --> (809) 0:PEGB6, pass, PUGB6
			8'd89 : rdata = 43'b1100011100001100000000000000000000000001110;
			// PEs: 38 -> 48
			// srcs: (255, 90)(809) 0 --> (809) 0:PEGB6, pass, PUGB6
			8'd90 : rdata = 43'b1100011100001100000000000000000000000001110;
			// PEs: 38 -> 48
			// srcs: (256, 91)(809) 0 --> (809) 0:PEGB6, pass, PUGB6
			8'd91 : rdata = 43'b1100011100001100000000000000000000000001110;
			// PEs: 38 -> 48
			// srcs: (257, 92)(809) 0 --> (809) 0:PEGB6, pass, PUGB6
			8'd92 : rdata = 43'b1100011100001100000000000000000000000001110;
			// PEs: 38 -> 56
			// srcs: (258, 93)(809) 0 --> (809) 0:PEGB6, pass, PUGB7
			8'd93 : rdata = 43'b1100011100001100000000000000000000000001111;
			// PEs: 38 -> 48
			// srcs: (259, 94)(809) 0 --> (809) 0:PEGB6, pass, PUGB6
			8'd94 : rdata = 43'b1100011100001100000000000000000000000001110;
			// PEs: 38 -> 56
			// srcs: (260, 95)(809) 0 --> (809) 0:PEGB6, pass, PUGB7
			8'd95 : rdata = 43'b1100011100001100000000000000000000000001111;
			// PEs: 38 -> 56
			// srcs: (261, 96)(809) 0 --> (809) 0:PEGB6, pass, PUGB7
			8'd96 : rdata = 43'b1100011100001100000000000000000000000001111;
			// PEs: 38 -> 56
			// srcs: (262, 97)(809) 0 --> (809) 0:PEGB6, pass, PUGB7
			8'd97 : rdata = 43'b1100011100001100000000000000000000000001111;
			// PEs: 38 -> 56
			// srcs: (263, 98)(809) 0 --> (809) 0:PEGB6, pass, PUGB7
			8'd98 : rdata = 43'b1100011100001100000000000000000000000001111;
			// PEs: 38 -> 56
			// srcs: (264, 99)(809) 0 --> (809) 0:PEGB6, pass, PUGB7
			8'd99 : rdata = 43'b1100011100001100000000000000000000000001111;
			// PEs: 38 -> 56
			// srcs: (265, 100)(809) 0 --> (809) 0:PEGB6, pass, PUGB7
			8'd100 : rdata = 43'b1100011100001100000000000000000000000001111;
			// PEs: 38 -> 56
			// srcs: (266, 101)(809) 0 --> (809) 0:PEGB6, pass, PUGB7
			8'd101 : rdata = 43'b1100011100001100000000000000000000000001111;
			// PEs: 38 -> 56
			// srcs: (267, 102)(809) 0 --> (809) 0:PEGB6, pass, PUGB7
			8'd102 : rdata = 43'b1100011100001100000000000000000000000001111;
			// PEs: 38 -> 56
			// srcs: (268, 103)(809) 0 --> (809) 0:PEGB6, pass, PUGB7
			8'd103 : rdata = 43'b1100011100001100000000000000000000000001111;
			// PEs: 38 -> 56
			// srcs: (269, 104)(809) 0 --> (809) 0:PEGB6, pass, PUGB7
			8'd104 : rdata = 43'b1100011100001100000000000000000000000001111;
			// PEs: 38 -> 0
			// srcs: (270, 105)(809) 0 --> (809) 0:PEGB6, pass, PUGB0
			8'd105 : rdata = 43'b1100011100001100000000000000000000000001000;
			// PEs: 38 -> 0
			// srcs: (271, 106)(809) 0 --> (809) 0:PEGB6, pass, PUGB0
			8'd106 : rdata = 43'b1100011100001100000000000000000000000001000;
			// PEs: 38 -> 0
			// srcs: (272, 107)(809) 0 --> (809) 0:PEGB6, pass, PUGB0
			8'd107 : rdata = 43'b1100011100001100000000000000000000000001000;
			// PEs: 38 -> 0
			// srcs: (273, 108)(809) 0 --> (809) 0:PEGB6, pass, PUGB0
			8'd108 : rdata = 43'b1100011100001100000000000000000000000001000;
			// PEs: 38 -> 56
			// srcs: (274, 109)(809) 0 --> (809) 0:PEGB6, pass, PUGB7
			8'd109 : rdata = 43'b1100011100001100000000000000000000000001111;
			// PEs: 38 -> 0
			// srcs: (275, 110)(809) 0 --> (809) 0:PEGB6, pass, PUGB0
			8'd110 : rdata = 43'b1100011100001100000000000000000000000001000;
			// PEs: 38 -> 0
			// srcs: (276, 111)(809) 0 --> (809) 0:PEGB6, pass, PUGB0
			8'd111 : rdata = 43'b1100011100001100000000000000000000000001000;
			// PEs: 38 -> 56
			// srcs: (277, 112)(809) 0 --> (809) 0:PEGB6, pass, PUGB7
			8'd112 : rdata = 43'b1100011100001100000000000000000000000001111;
			// PEs: 38 -> 0
			// srcs: (278, 113)(809) 0 --> (809) 0:PEGB6, pass, PUGB0
			8'd113 : rdata = 43'b1100011100001100000000000000000000000001000;
			// PEs: 38 -> 8
			// srcs: (279, 114)(809) 0 --> (809) 0:PEGB6, pass, PUGB1
			8'd114 : rdata = 43'b1100011100001100000000000000000000000001001;
			// PEs: 38 -> 56
			// srcs: (280, 115)(809) 0 --> (809) 0:PEGB6, pass, PUGB7
			8'd115 : rdata = 43'b1100011100001100000000000000000000000001111;
			// PEs: 38 -> 8
			// srcs: (281, 116)(809) 0 --> (809) 0:PEGB6, pass, PUGB1
			8'd116 : rdata = 43'b1100011100001100000000000000000000000001001;
			// PEs: 38 -> 8
			// srcs: (282, 117)(809) 0 --> (809) 0:PEGB6, pass, PUGB1
			8'd117 : rdata = 43'b1100011100001100000000000000000000000001001;
			// PEs: 38 -> 0
			// srcs: (283, 118)(809) 0 --> (809) 0:PEGB6, pass, PUGB0
			8'd118 : rdata = 43'b1100011100001100000000000000000000000001000;
			// PEs: 38 -> 8
			// srcs: (284, 119)(809) 0 --> (809) 0:PEGB6, pass, PUGB1
			8'd119 : rdata = 43'b1100011100001100000000000000000000000001001;
			// PEs: 38 -> 8
			// srcs: (285, 120)(809) 0 --> (809) 0:PEGB6, pass, PUGB1
			8'd120 : rdata = 43'b1100011100001100000000000000000000000001001;
			// PEs: 38 -> 0
			// srcs: (286, 121)(809) 0 --> (809) 0:PEGB6, pass, PUGB0
			8'd121 : rdata = 43'b1100011100001100000000000000000000000001000;
			// PEs: 38 -> 8
			// srcs: (287, 122)(809) 0 --> (809) 0:PEGB6, pass, PUGB1
			8'd122 : rdata = 43'b1100011100001100000000000000000000000001001;
			// PEs: 38 -> 8
			// srcs: (288, 123)(809) 0 --> (809) 0:PEGB6, pass, PUGB1
			8'd123 : rdata = 43'b1100011100001100000000000000000000000001001;
			// PEs: 38 -> 0
			// srcs: (289, 124)(809) 0 --> (809) 0:PEGB6, pass, PUGB0
			8'd124 : rdata = 43'b1100011100001100000000000000000000000001000;
			// PEs: 38 -> 16
			// srcs: (290, 125)(809) 0 --> (809) 0:PEGB6, pass, PUGB2
			8'd125 : rdata = 43'b1100011100001100000000000000000000000001010;
			// PEs: 38 -> 16
			// srcs: (291, 126)(809) 0 --> (809) 0:PEGB6, pass, PUGB2
			8'd126 : rdata = 43'b1100011100001100000000000000000000000001010;
			// PEs: 38 -> 0
			// srcs: (292, 127)(809) 0 --> (809) 0:PEGB6, pass, PUGB0
			8'd127 : rdata = 43'b1100011100001100000000000000000000000001000;
			// PEs: 38 -> 16
			// srcs: (293, 128)(809) 0 --> (809) 0:PEGB6, pass, PUGB2
			8'd128 : rdata = 43'b1100011100001100000000000000000000000001010;
			// PEs: 38 -> 16
			// srcs: (294, 129)(809) 0 --> (809) 0:PEGB6, pass, PUGB2
			8'd129 : rdata = 43'b1100011100001100000000000000000000000001010;
			// PEs: 38 -> 16
			// srcs: (295, 130)(809) 0 --> (809) 0:PEGB6, pass, PUGB2
			8'd130 : rdata = 43'b1100011100001100000000000000000000000001010;
			// PEs: 38 -> 16
			// srcs: (296, 131)(809) 0 --> (809) 0:PEGB6, pass, PUGB2
			8'd131 : rdata = 43'b1100011100001100000000000000000000000001010;
			// PEs: 38 -> 16
			// srcs: (297, 132)(809) 0 --> (809) 0:PEGB6, pass, PUGB2
			8'd132 : rdata = 43'b1100011100001100000000000000000000000001010;
			// PEs: 38 -> 24
			// srcs: (298, 133)(809) 0 --> (809) 0:PEGB6, pass, PUGB3
			8'd133 : rdata = 43'b1100011100001100000000000000000000000001011;
			// PEs: 38 -> 0
			// srcs: (299, 134)(809) 0 --> (809) 0:PEGB6, pass, PUGB0
			8'd134 : rdata = 43'b1100011100001100000000000000000000000001000;
			// PEs: 38 -> 24
			// srcs: (300, 135)(809) 0 --> (809) 0:PEGB6, pass, PUGB3
			8'd135 : rdata = 43'b1100011100001100000000000000000000000001011;
			// PEs: 38 -> 24
			// srcs: (301, 136)(809) 0 --> (809) 0:PEGB6, pass, PUGB3
			8'd136 : rdata = 43'b1100011100001100000000000000000000000001011;
			// PEs: 38 -> 0
			// srcs: (302, 137)(809) 0 --> (809) 0:PEGB6, pass, PUGB0
			8'd137 : rdata = 43'b1100011100001100000000000000000000000001000;
			// PEs: 38 -> 24
			// srcs: (303, 138)(809) 0 --> (809) 0:PEGB6, pass, PUGB3
			8'd138 : rdata = 43'b1100011100001100000000000000000000000001011;
			// PEs: 38 -> 24
			// srcs: (304, 139)(809) 0 --> (809) 0:PEGB6, pass, PUGB3
			8'd139 : rdata = 43'b1100011100001100000000000000000000000001011;
			// PEs: 38 -> 0
			// srcs: (305, 140)(809) 0 --> (809) 0:PEGB6, pass, PUGB0
			8'd140 : rdata = 43'b1100011100001100000000000000000000000001000;
			// PEs: 38 -> 24
			// srcs: (306, 141)(809) 0 --> (809) 0:PEGB6, pass, PUGB3
			8'd141 : rdata = 43'b1100011100001100000000000000000000000001011;
			// PEs: 38 -> 24
			// srcs: (307, 142)(809) 0 --> (809) 0:PEGB6, pass, PUGB3
			8'd142 : rdata = 43'b1100011100001100000000000000000000000001011;
			// PEs: 38 -> 8
			// srcs: (308, 143)(809) 0 --> (809) 0:PEGB6, pass, PUGB1
			8'd143 : rdata = 43'b1100011100001100000000000000000000000001001;
			// PEs: 38 -> 8
			// srcs: (311, 144)(809) 0 --> (809) 0:PEGB6, pass, PUGB1
			8'd144 : rdata = 43'b1100011100001100000000000000000000000001001;
			// PEs: 38 -> 8
			// srcs: (314, 145)(809) 0 --> (809) 0:PEGB6, pass, PUGB1
			8'd145 : rdata = 43'b1100011100001100000000000000000000000001001;
			// PEs: 38 -> 8
			// srcs: (317, 146)(809) 0 --> (809) 0:PEGB6, pass, PUGB1
			8'd146 : rdata = 43'b1100011100001100000000000000000000000001001;
			// PEs: 38 -> 40
			// srcs: (319, 147)(809) 0 --> (809) 0:PEGB6, pass, PUNB
			8'd147 : rdata = 43'b1100011100001100000000000000000001000000000;
			// PEs: 38 -> 40
			// srcs: (320, 148)(809) 0 --> (809) 0:PEGB6, pass, PUNB
			8'd148 : rdata = 43'b1100011100001100000000000000000001000000000;
			// PEs: 38 -> 40
			// srcs: (321, 149)(809) 0 --> (809) 0:PEGB6, pass, PUNB
			8'd149 : rdata = 43'b1100011100001100000000000000000001000000000;
			// PEs: 38 -> 40
			// srcs: (322, 150)(809) 0 --> (809) 0:PEGB6, pass, PUNB
			8'd150 : rdata = 43'b1100011100001100000000000000000001000000000;
			// PEs: 38 -> 40
			// srcs: (323, 151)(809) 0 --> (809) 0:PEGB6, pass, PUNB
			8'd151 : rdata = 43'b1100011100001100000000000000000001000000000;
			// PEs: 38 -> 8
			// srcs: (324, 152)(809) 0 --> (809) 0:PEGB6, pass, PUGB1
			8'd152 : rdata = 43'b1100011100001100000000000000000000000001001;
			// PEs: 38 -> 40
			// srcs: (325, 153)(809) 0 --> (809) 0:PEGB6, pass, PUNB
			8'd153 : rdata = 43'b1100011100001100000000000000000001000000000;
			// PEs: 38 -> 40
			// srcs: (326, 154)(809) 0 --> (809) 0:PEGB6, pass, PUNB
			8'd154 : rdata = 43'b1100011100001100000000000000000001000000000;
			// PEs: 38 -> 8
			// srcs: (327, 155)(809) 0 --> (809) 0:PEGB6, pass, PUGB1
			8'd155 : rdata = 43'b1100011100001100000000000000000000000001001;
			// PEs: 38 -> 48
			// srcs: (328, 156)(809) 0 --> (809) 0:PEGB6, pass, PUGB6
			8'd156 : rdata = 43'b1100011100001100000000000000000000000001110;
			// PEs: 38 -> 48
			// srcs: (329, 157)(809) 0 --> (809) 0:PEGB6, pass, PUGB6
			8'd157 : rdata = 43'b1100011100001100000000000000000000000001110;
			// PEs: 38 -> 8
			// srcs: (330, 158)(809) 0 --> (809) 0:PEGB6, pass, PUGB1
			8'd158 : rdata = 43'b1100011100001100000000000000000000000001001;
			// PEs: 38 -> 48
			// srcs: (331, 159)(809) 0 --> (809) 0:PEGB6, pass, PUGB6
			8'd159 : rdata = 43'b1100011100001100000000000000000000000001110;
			// PEs: 38 -> 48
			// srcs: (332, 160)(809) 0 --> (809) 0:PEGB6, pass, PUGB6
			8'd160 : rdata = 43'b1100011100001100000000000000000000000001110;
			// PEs: 38 -> 16
			// srcs: (333, 161)(809) 0 --> (809) 0:PEGB6, pass, PUGB2
			8'd161 : rdata = 43'b1100011100001100000000000000000000000001010;
			// PEs: 38 -> 48
			// srcs: (334, 162)(809) 0 --> (809) 0:PEGB6, pass, PUGB6
			8'd162 : rdata = 43'b1100011100001100000000000000000000000001110;
			// PEs: 38 -> 48
			// srcs: (335, 163)(809) 0 --> (809) 0:PEGB6, pass, PUGB6
			8'd163 : rdata = 43'b1100011100001100000000000000000000000001110;
			// PEs: 38 -> 16
			// srcs: (336, 164)(809) 0 --> (809) 0:PEGB6, pass, PUGB2
			8'd164 : rdata = 43'b1100011100001100000000000000000000000001010;
			// PEs: 38 -> 48
			// srcs: (337, 165)(809) 0 --> (809) 0:PEGB6, pass, PUGB6
			8'd165 : rdata = 43'b1100011100001100000000000000000000000001110;
			// PEs: 38 -> 56
			// srcs: (338, 166)(809) 0 --> (809) 0:PEGB6, pass, PUGB7
			8'd166 : rdata = 43'b1100011100001100000000000000000000000001111;
			// PEs: 38 -> 16
			// srcs: (339, 167)(809) 0 --> (809) 0:PEGB6, pass, PUGB2
			8'd167 : rdata = 43'b1100011100001100000000000000000000000001010;
			// PEs: 38 -> 56
			// srcs: (340, 168)(809) 0 --> (809) 0:PEGB6, pass, PUGB7
			8'd168 : rdata = 43'b1100011100001100000000000000000000000001111;
			// PEs: 38 -> 56
			// srcs: (341, 169)(809) 0 --> (809) 0:PEGB6, pass, PUGB7
			8'd169 : rdata = 43'b1100011100001100000000000000000000000001111;
			// PEs: 38 -> 16
			// srcs: (342, 170)(809) 0 --> (809) 0:PEGB6, pass, PUGB2
			8'd170 : rdata = 43'b1100011100001100000000000000000000000001010;
			// PEs: 38 -> 56
			// srcs: (343, 171)(809) 0 --> (809) 0:PEGB6, pass, PUGB7
			8'd171 : rdata = 43'b1100011100001100000000000000000000000001111;
			// PEs: 38 -> 56
			// srcs: (344, 172)(809) 0 --> (809) 0:PEGB6, pass, PUGB7
			8'd172 : rdata = 43'b1100011100001100000000000000000000000001111;
			// PEs: 38 -> 56
			// srcs: (345, 173)(809) 0 --> (809) 0:PEGB6, pass, PUGB7
			8'd173 : rdata = 43'b1100011100001100000000000000000000000001111;
			// PEs: 38 -> 56
			// srcs: (346, 174)(809) 0 --> (809) 0:PEGB6, pass, PUGB7
			8'd174 : rdata = 43'b1100011100001100000000000000000000000001111;
			// PEs: 38 -> 0
			// srcs: (347, 175)(809) 0 --> (809) 0:PEGB6, pass, PUGB0
			8'd175 : rdata = 43'b1100011100001100000000000000000000000001000;
			// PEs: 38 -> 0
			// srcs: (348, 176)(809) 0 --> (809) 0:PEGB6, pass, PUGB0
			8'd176 : rdata = 43'b1100011100001100000000000000000000000001000;
			// PEs: 38 -> 16
			// srcs: (349, 177)(809) 0 --> (809) 0:PEGB6, pass, PUGB2
			8'd177 : rdata = 43'b1100011100001100000000000000000000000001010;
			// PEs: 38 -> 0
			// srcs: (350, 178)(809) 0 --> (809) 0:PEGB6, pass, PUGB0
			8'd178 : rdata = 43'b1100011100001100000000000000000000000001000;
			// PEs: 38 -> 0
			// srcs: (351, 179)(809) 0 --> (809) 0:PEGB6, pass, PUGB0
			8'd179 : rdata = 43'b1100011100001100000000000000000000000001000;
			// PEs: 38 -> 16
			// srcs: (352, 180)(809) 0 --> (809) 0:PEGB6, pass, PUGB2
			8'd180 : rdata = 43'b1100011100001100000000000000000000000001010;
			// PEs: 38 -> 0
			// srcs: (353, 181)(809) 0 --> (809) 0:PEGB6, pass, PUGB0
			8'd181 : rdata = 43'b1100011100001100000000000000000000000001000;
			// PEs: 38 -> 0
			// srcs: (354, 182)(809) 0 --> (809) 0:PEGB6, pass, PUGB0
			8'd182 : rdata = 43'b1100011100001100000000000000000000000001000;
			// PEs: 38 -> 16
			// srcs: (355, 183)(809) 0 --> (809) 0:PEGB6, pass, PUGB2
			8'd183 : rdata = 43'b1100011100001100000000000000000000000001010;
			// PEs: 38 -> 0
			// srcs: (356, 184)(809) 0 --> (809) 0:PEGB6, pass, PUGB0
			8'd184 : rdata = 43'b1100011100001100000000000000000000000001000;
			// PEs: 38 -> 8
			// srcs: (357, 185)(809) 0 --> (809) 0:PEGB6, pass, PUGB1
			8'd185 : rdata = 43'b1100011100001100000000000000000000000001001;
			// PEs: 38 -> 24
			// srcs: (358, 186)(809) 0 --> (809) 0:PEGB6, pass, PUGB3
			8'd186 : rdata = 43'b1100011100001100000000000000000000000001011;
			// PEs: 38 -> 8
			// srcs: (359, 187)(809) 0 --> (809) 0:PEGB6, pass, PUGB1
			8'd187 : rdata = 43'b1100011100001100000000000000000000000001001;
			// PEs: 38 -> 8
			// srcs: (360, 188)(809) 0 --> (809) 0:PEGB6, pass, PUGB1
			8'd188 : rdata = 43'b1100011100001100000000000000000000000001001;
			// PEs: 38 -> 24
			// srcs: (361, 189)(809) 0 --> (809) 0:PEGB6, pass, PUGB3
			8'd189 : rdata = 43'b1100011100001100000000000000000000000001011;
			// PEs: 38 -> 8
			// srcs: (362, 190)(809) 0 --> (809) 0:PEGB6, pass, PUGB1
			8'd190 : rdata = 43'b1100011100001100000000000000000000000001001;
			// PEs: 38 -> 8
			// srcs: (363, 191)(809) 0 --> (809) 0:PEGB6, pass, PUGB1
			8'd191 : rdata = 43'b1100011100001100000000000000000000000001001;
			// PEs: 38 -> 24
			// srcs: (364, 192)(809) 0 --> (809) 0:PEGB6, pass, PUGB3
			8'd192 : rdata = 43'b1100011100001100000000000000000000000001011;
			// PEs: 38 -> 8
			// srcs: (365, 193)(809) 0 --> (809) 0:PEGB6, pass, PUGB1
			8'd193 : rdata = 43'b1100011100001100000000000000000000000001001;
			// PEs: 38 -> 8
			// srcs: (366, 194)(809) 0 --> (809) 0:PEGB6, pass, PUGB1
			8'd194 : rdata = 43'b1100011100001100000000000000000000000001001;
			// PEs: 38 -> 24
			// srcs: (367, 195)(809) 0 --> (809) 0:PEGB6, pass, PUGB3
			8'd195 : rdata = 43'b1100011100001100000000000000000000000001011;
			// PEs: 38 -> 16
			// srcs: (368, 196)(809) 0 --> (809) 0:PEGB6, pass, PUGB2
			8'd196 : rdata = 43'b1100011100001100000000000000000000000001010;
			// PEs: 38 -> 16
			// srcs: (369, 197)(809) 0 --> (809) 0:PEGB6, pass, PUGB2
			8'd197 : rdata = 43'b1100011100001100000000000000000000000001010;
			// PEs: 38 -> 16
			// srcs: (370, 198)(809) 0 --> (809) 0:PEGB6, pass, PUGB2
			8'd198 : rdata = 43'b1100011100001100000000000000000000000001010;
			// PEs: 38 -> 16
			// srcs: (371, 199)(809) 0 --> (809) 0:PEGB6, pass, PUGB2
			8'd199 : rdata = 43'b1100011100001100000000000000000000000001010;
			// PEs: 38 -> 16
			// srcs: (372, 200)(809) 0 --> (809) 0:PEGB6, pass, PUGB2
			8'd200 : rdata = 43'b1100011100001100000000000000000000000001010;
			// PEs: 38 -> 16
			// srcs: (373, 201)(809) 0 --> (809) 0:PEGB6, pass, PUGB2
			8'd201 : rdata = 43'b1100011100001100000000000000000000000001010;
			// PEs: 38 -> 24
			// srcs: (374, 202)(809) 0 --> (809) 0:PEGB6, pass, PUGB3
			8'd202 : rdata = 43'b1100011100001100000000000000000000000001011;
			// PEs: 38 -> 16
			// srcs: (375, 203)(809) 0 --> (809) 0:PEGB6, pass, PUGB2
			8'd203 : rdata = 43'b1100011100001100000000000000000000000001010;
			// PEs: 38 -> 24
			// srcs: (376, 204)(809) 0 --> (809) 0:PEGB6, pass, PUGB3
			8'd204 : rdata = 43'b1100011100001100000000000000000000000001011;
			// PEs: 38 -> 24
			// srcs: (377, 205)(809) 0 --> (809) 0:PEGB6, pass, PUGB3
			8'd205 : rdata = 43'b1100011100001100000000000000000000000001011;
			// PEs: 38 -> 24
			// srcs: (378, 206)(809) 0 --> (809) 0:PEGB6, pass, PUGB3
			8'd206 : rdata = 43'b1100011100001100000000000000000000000001011;
			// PEs: 38 -> 24
			// srcs: (379, 207)(809) 0 --> (809) 0:PEGB6, pass, PUGB3
			8'd207 : rdata = 43'b1100011100001100000000000000000000000001011;
			// PEs: 38 -> 24
			// srcs: (380, 208)(809) 0 --> (809) 0:PEGB6, pass, PUGB3
			8'd208 : rdata = 43'b1100011100001100000000000000000000000001011;
			// PEs: 38 -> 24
			// srcs: (381, 209)(809) 0 --> (809) 0:PEGB6, pass, PUGB3
			8'd209 : rdata = 43'b1100011100001100000000000000000000000001011;
			// PEs: 38 -> 24
			// srcs: (382, 210)(809) 0 --> (809) 0:PEGB6, pass, PUGB3
			8'd210 : rdata = 43'b1100011100001100000000000000000000000001011;
			// PEs: 38 -> 24
			// srcs: (384, 211)(809) 0 --> (809) 0:PEGB6, pass, PUGB3
			8'd211 : rdata = 43'b1100011100001100000000000000000000000001011;
			// PEs: 38 -> 24
			// srcs: (385, 212)(809) 0 --> (809) 0:PEGB6, pass, PUGB3
			8'd212 : rdata = 43'b1100011100001100000000000000000000000001011;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 33) begin
	always @(*) begin
		case(address)
			// PEs: 33, 33 -> 38
			// srcs: (1, 0)(42) -2, (243) -3 --> (443) 6:ND0, NW0, *, PEGB6
			8'd0 : rdata = 43'b0001101100000000010000000000000000011100000;
			// PEs: 33, 33 -> 34
			// srcs: (2, 1)(120) 1, (321) -1 --> (521) -1:ND1, NW1, *, PENB
			8'd1 : rdata = 43'b0001101100000001010000000010000000100000000;
			// PEs: 33, 33 -> 34
			// srcs: (3, 2)(198) 1, (399) 2 --> (599) 2:ND2, NW2, *, PENB
			8'd2 : rdata = 43'b0001101100000010010000000100000000100000000;
			// PEs: 33, 33 -> 33
			// srcs: (4, 3)(194) 0, (395) 0 --> (595) 0:ND3, NW3, *, NI0
			8'd3 : rdata = 43'b0001101100000011010000000111000000000000000;
			// PEs: 32, 38 -> 32
			// srcs: (21, 4)(611) -3, (414) 0 --> (612) -3:PENB, PEGB6, +, PEGB0
			8'd4 : rdata = 43'b0000111011111110111000011000000000010000000;
			// PEs: 32 -> 
			// srcs: (22, 5)(420) 3 --> (420) 3:PENB, pass, 
			8'd5 : rdata = 43'b1100011011111110000000000000000000000000000;
			// PEs: 32, 33 -> 32
			// srcs: (28, 6)(617) -1, (420) 3 --> (618) 2:PENB, ALU, +, PEGB0
			8'd6 : rdata = 43'b0000111011111110001111111110000000010000000;
			// PEs: 32 -> 
			// srcs: (30, 7)(442) 0 --> (442) 0:PENB, pass, 
			8'd7 : rdata = 43'b1100011011111110000000000000000000000000000;
			// PEs: 32, 33 -> 32
			// srcs: (36, 8)(637) 9, (442) 0 --> (638) 9:PENB, ALU, +, PEGB0
			8'd8 : rdata = 43'b0000111011111110001111111110000000010000000;
			// PEs: 34, 32 -> 32
			// srcs: (43, 9)(718) -1, (523) 6 --> (719) 5:PEGB2, PENB, +, PEGB0
			8'd9 : rdata = 43'b0000111100000100110111111100000000010000000;
			// PEs: 38, 32 -> 35
			// srcs: (60, 10)(723) 3, (529) -6 --> (724) -3:PEGB6, PENB, +, PEGB3
			8'd10 : rdata = 43'b0000111100001100110111111100000000010110000;
			// PEs: 32 -> 
			// srcs: (62, 11)(548) 0 --> (548) 0:PENB, pass, 
			8'd11 : rdata = 43'b1100011011111110000000000000000000000000000;
			// PEs: 32, 33 -> 32
			// srcs: (68, 12)(742) 9, (548) 0 --> (743) 9:PENB, ALU, +, PEGB0
			8'd12 : rdata = 43'b0000111011111110001111111110000000010000000;
			// PEs: 32 -> 
			// srcs: (70, 13)(576) 1 --> (576) 1:PENB, pass, 
			8'd13 : rdata = 43'b1100011011111110000000000000000000000000000;
			// PEs: 32, 33 -> 33
			// srcs: (76, 14)(770) 0, (576) 1 --> (771) 1:PENB, ALU, +, NI1
			8'd14 : rdata = 43'b0000111011111110001111111111010000000000000;
			// PEs: 32, 33 -> 33
			// srcs: (77, 15)(789) -4, (595) 0 --> (790) -4:PENB, NI0, +, NI2
			8'd15 : rdata = 43'b0000111011111110101000000001100000000000000;
			// PEs: 32, 34 -> 34
			// srcs: (85, 16)(791) 3, (598) -6 --> (792) -3:PENB, PEGB2, +, PENB
			8'd16 : rdata = 43'b0000111011111110111000001000000000100000000;
			// PEs: 33, 32 -> 33
			// srcs: (86, 17)(771) 1, (773) -2 --> (774) -1:NI1, PENB, +, NI0
			8'd17 : rdata = 43'b0000110100000001110111111101000000000000000;
			// PEs: 33 -> 34
			// srcs: (92, 18)(790) -4 --> (790) -4:NI2, pass, PENB
			8'd18 : rdata = 43'b1100010100000010000000000000000000100000000;
			// PEs: 32, 33 -> 32
			// srcs: (96, 19)(769) 8, (774) -1 --> (775) 7:PENB, NI0, +, PEGB0
			8'd19 : rdata = 43'b0000111011111110101000000000000000010000000;
			// PEs: 32, 37 -> 32
			// srcs: (112, 20)(788) -13, (799) -7 --> (800) -20:PENB, PEGB5, +, PEGB0
			8'd20 : rdata = 43'b0000111011111110111000010100000000010000000;
			// PEs: 38, 33 -> 34
			// srcs: (231, 21)(809) 0, (42) -2 --> (848) 0:PEGB6, ND0, *, PENB
			8'd21 : rdata = 43'b0001111100001100011000000000000000100000000;
			// PEs: 33, 34 -> 33
			// srcs: (240, 26)(243) -3, (1048) 0 --> (1248) -3:NW0, PEGB2, -, NW0
			8'd22 : rdata = 43'b0001001000000000111000001000001000000000000;
			// PEs: 38, 33 -> 34
			// srcs: (309, 22)(809) 0, (120) 1 --> (926) 0:PEGB6, ND1, *, PENB
			8'd23 : rdata = 43'b0001111100001100011000000010000000100000000;
			// PEs: 33, 34 -> 33
			// srcs: (318, 27)(321) -1, (1126) 0 --> (1326) -1:NW1, PEGB2, -, NW1
			8'd24 : rdata = 43'b0001001000000001111000001000001010000000000;
			// PEs: 38, 33 -> 
			// srcs: (383, 23)(809) 0, (194) 0 --> (1000) 0:PEGB6, ND3, *, 
			8'd25 : rdata = 43'b0001111100001100011000000110000000000000000;
			// PEs: 33, 33 -> 33
			// srcs: (386, 25)(3) 1, (1000) 0 --> (1200) 0:NM0, ALU, *, NI0
			8'd26 : rdata = 43'b0001110000000000001111111111000000000000000;
			// PEs: 38, 33 -> 34
			// srcs: (387, 24)(809) 0, (198) 1 --> (1004) 0:PEGB6, ND2, *, PENB
			8'd27 : rdata = 43'b0001111100001100011000000100000000100000000;
			// PEs: 33, 33 -> 33
			// srcs: (389, 28)(395) 0, (1200) 0 --> (1400) 0:NW3, NI0, -, NW3
			8'd28 : rdata = 43'b0001001000000011101000000000001110000000000;
			// PEs: 33, 34 -> 33
			// srcs: (396, 29)(399) 2, (1204) 0 --> (1404) 2:NW2, PEGB2, -, NW2
			8'd29 : rdata = 43'b0001001000000010111000001000001100000000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 34) begin
	always @(*) begin
		case(address)
			// PEs: 34, 34 -> 38
			// srcs: (1, 0)(43) 1, (244) 2 --> (444) 2:ND0, NW0, *, PEGB6
			8'd0 : rdata = 43'b0001101100000000010000000000000000011100000;
			// PEs: 34, 34 -> 34
			// srcs: (2, 1)(121) 0, (322) -3 --> (522) 0:ND1, NW1, *, NI0
			8'd1 : rdata = 43'b0001101100000001010000000011000000000000000;
			// PEs: 34, 34 -> 34
			// srcs: (3, 2)(199) 0, (400) -2 --> (600) 0:ND2, NW2, *, NI1
			8'd2 : rdata = 43'b0001101100000010010000000101010000000000000;
			// PEs: 34, 34 -> 34
			// srcs: (4, 3)(197) -3, (398) 2 --> (598) -6:ND3, NW3, *, NI2
			8'd3 : rdata = 43'b0001101100000011010000000111100000000000000;
			// PEs: 33, 34 -> 33
			// srcs: (5, 4)(521) -1, (522) 0 --> (718) -1:PENB, NI0, +, PEGB1
			8'd4 : rdata = 43'b0000111011111110101000000000000000010010000;
			// PEs: 33, 34 -> 35
			// srcs: (6, 5)(599) 2, (600) 0 --> (794) 2:PENB, NI1, +, PENB
			8'd5 : rdata = 43'b0000111011111110101000000010000000100000000;
			// PEs: 34 -> 33
			// srcs: (80, 6)(598) -6 --> (598) -6:NI2, pass, PEGB1
			8'd6 : rdata = 43'b1100010100000010000000000000000000010010000;
			// PEs: 33 -> 
			// srcs: (87, 7)(792) -3 --> (792) -3:PENB, pass, 
			8'd7 : rdata = 43'b1100011011111110000000000000000000000000000;
			// PEs: 33, 34 -> 37
			// srcs: (94, 8)(790) -4, (792) -3 --> (793) -7:PENB, ALU, +, PEGB5
			8'd8 : rdata = 43'b0000111011111110001111111110000000011010000;
			// PEs: 38, 34 -> 35
			// srcs: (232, 9)(809) 0, (43) 1 --> (849) 0:PEGB6, ND0, *, PENB
			8'd9 : rdata = 43'b0001111100001100011000000000000000100000000;
			// PEs: 34, 33 -> 33
			// srcs: (234, 13)(3) 1, (848) 0 --> (1048) 0:NM0, PENB, *, PEGB1
			8'd10 : rdata = 43'b0001110000000000110111111100000000010010000;
			// PEs: 34, 35 -> 34
			// srcs: (241, 17)(244) 2, (1049) 0 --> (1249) 2:NW0, PEGB3, -, NW0
			8'd11 : rdata = 43'b0001001000000000111000001100001000000000000;
			// PEs: 38, 34 -> 35
			// srcs: (310, 10)(809) 0, (121) 0 --> (927) 0:PEGB6, ND1, *, PENB
			8'd12 : rdata = 43'b0001111100001100011000000010000000100000000;
			// PEs: 34, 33 -> 33
			// srcs: (312, 14)(3) 1, (926) 0 --> (1126) 0:NM0, PENB, *, PEGB1
			8'd13 : rdata = 43'b0001110000000000110111111100000000010010000;
			// PEs: 34, 35 -> 34
			// srcs: (319, 18)(322) -3, (1127) 0 --> (1327) -3:NW1, PEGB3, -, NW1
			8'd14 : rdata = 43'b0001001000000001111000001100001010000000000;
			// PEs: 38, 34 -> 34
			// srcs: (386, 11)(809) 0, (197) -3 --> (1003) 0:PEGB6, ND3, *, NI0
			8'd15 : rdata = 43'b0001111100001100011000000111000000000000000;
			// PEs: 38, 34 -> 35
			// srcs: (388, 12)(809) 0, (199) 0 --> (1005) 0:PEGB6, ND2, *, PENB
			8'd16 : rdata = 43'b0001111100001100011000000100000000100000000;
			// PEs: 34, 34 -> 34
			// srcs: (389, 15)(3) 1, (1003) 0 --> (1203) 0:NM0, NI0, *, NI1
			8'd17 : rdata = 43'b0001110000000000101000000001010000000000000;
			// PEs: 34, 33 -> 33
			// srcs: (390, 16)(3) 1, (1004) 0 --> (1204) 0:NM0, PENB, *, PEGB1
			8'd18 : rdata = 43'b0001110000000000110111111100000000010010000;
			// PEs: 34, 34 -> 34
			// srcs: (392, 19)(398) 2, (1203) 0 --> (1403) 2:NW3, NI1, -, NW3
			8'd19 : rdata = 43'b0001001000000011101000000010001110000000000;
			// PEs: 34, 35 -> 34
			// srcs: (397, 20)(400) -2, (1205) 0 --> (1405) -2:NW2, PEGB3, -, NW2
			8'd20 : rdata = 43'b0001001000000010111000001100001100000000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 35) begin
	always @(*) begin
		case(address)
			// PEs: 35, 35 -> 39
			// srcs: (1, 0)(45) 0, (246) -2 --> (446) 0:ND0, NW0, *, PEGB7
			8'd0 : rdata = 43'b0001101100000000010000000000000000011110000;
			// PEs: 35, 35 -> 36
			// srcs: (2, 1)(123) 2, (324) 1 --> (524) 2:ND1, NW1, *, PENB
			8'd1 : rdata = 43'b0001101100000001010000000010000000100000000;
			// PEs: 35, 35 -> 36
			// srcs: (3, 2)(201) 2, (402) 2 --> (602) 4:ND2, NW2, *, PENB
			8'd2 : rdata = 43'b0001101100000010010000000100000000100000000;
			// PEs: 35, 35 -> 
			// srcs: (4, 3)(200) 0, (401) 0 --> (601) 0:ND3, NW3, *, 
			8'd3 : rdata = 43'b0001101100000011010000000110000000000000000;
			// PEs: 34, 35 -> 39
			// srcs: (9, 4)(794) 2, (601) 0 --> (795) 2:PENB, ALU, +, PEGB7
			8'd4 : rdata = 43'b0000111011111110001111111110000000011110000;
			// PEs: 32 -> 
			// srcs: (82, 5)(722) 6 --> (722) 6:PEGB0, pass, 
			8'd5 : rdata = 43'b1100011100000000000000000000000000000000000;
			// PEs: 35, 33 -> 32
			// srcs: (84, 6)(722) 6, (724) -3 --> (725) 3:ALU, PEGB1, +, PEGB0
			8'd6 : rdata = 43'b0000100111111111111000000100000000010000000;
			// PEs: 38, 35 -> 36
			// srcs: (234, 7)(809) 0, (45) 0 --> (851) 0:PEGB6, ND0, *, PENB
			8'd7 : rdata = 43'b0001111100001100011000000000000000100000000;
			// PEs: 35, 34 -> 34
			// srcs: (235, 11)(3) 1, (849) 0 --> (1049) 0:NM0, PENB, *, PEGB2
			8'd8 : rdata = 43'b0001110000000000110111111100000000010100000;
			// PEs: 35, 36 -> 35
			// srcs: (243, 16)(246) -2, (1051) 0 --> (1251) -2:NW0, PEGB4, -, NW0
			8'd9 : rdata = 43'b0001001000000000111000010000001000000000000;
			// PEs: 38, 35 -> 35
			// srcs: (312, 8)(809) 0, (123) 2 --> (929) 0:PEGB6, ND1, *, NI0
			8'd10 : rdata = 43'b0001111100001100011000000011000000000000000;
			// PEs: 35, 34 -> 34
			// srcs: (313, 12)(3) 1, (927) 0 --> (1127) 0:NM0, PENB, *, PEGB2
			8'd11 : rdata = 43'b0001110000000000110111111100000000010100000;
			// PEs: 35, 35 -> 
			// srcs: (315, 13)(3) 1, (929) 0 --> (1129) 0:NM0, NI0, *, 
			8'd12 : rdata = 43'b0001110000000000101000000000000000000000000;
			// PEs: 35, 35 -> 35
			// srcs: (318, 17)(324) 1, (1129) 0 --> (1329) 1:NW1, ALU, -, NW1
			8'd13 : rdata = 43'b0001001000000001001111111110001010000000000;
			// PEs: 38, 35 -> 35
			// srcs: (389, 9)(809) 0, (200) 0 --> (1006) 0:PEGB6, ND3, *, NI0
			8'd14 : rdata = 43'b0001111100001100011000000111000000000000000;
			// PEs: 38, 35 -> 36
			// srcs: (390, 10)(809) 0, (201) 2 --> (1007) 0:PEGB6, ND2, *, PENB
			8'd15 : rdata = 43'b0001111100001100011000000100000000100000000;
			// PEs: 35, 34 -> 34
			// srcs: (391, 14)(3) 1, (1005) 0 --> (1205) 0:NM0, PENB, *, PEGB2
			8'd16 : rdata = 43'b0001110000000000110111111100000000010100000;
			// PEs: 35, 35 -> 
			// srcs: (392, 15)(3) 1, (1006) 0 --> (1206) 0:NM0, NI0, *, 
			8'd17 : rdata = 43'b0001110000000000101000000000000000000000000;
			// PEs: 35, 35 -> 35
			// srcs: (395, 18)(401) 0, (1206) 0 --> (1406) 0:NW3, ALU, -, NW3
			8'd18 : rdata = 43'b0001001000000011001111111110001110000000000;
			// PEs: 35, 36 -> 35
			// srcs: (399, 19)(402) 2, (1207) 0 --> (1407) 2:NW2, PEGB4, -, NW2
			8'd19 : rdata = 43'b0001001000000010111000010000001100000000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 36) begin
	always @(*) begin
		case(address)
			// PEs: 36, 36 -> 39
			// srcs: (1, 0)(46) 2, (247) 2 --> (447) 4:ND0, NW0, *, PEGB7
			8'd0 : rdata = 43'b0001101100000000010000000000000000011110000;
			// PEs: 36, 36 -> 36
			// srcs: (2, 1)(124) -3, (325) -2 --> (525) 6:ND1, NW1, *, NI0
			8'd1 : rdata = 43'b0001101100000001010000000011000000000000000;
			// PEs: 36, 36 -> 36
			// srcs: (3, 2)(202) 0, (403) 1 --> (603) 0:ND2, NW2, *, NI1
			8'd2 : rdata = 43'b0001101100000010010000000101010000000000000;
			// PEs: 36, 36 -> 36
			// srcs: (4, 3)(203) 2, (404) -3 --> (604) -6:ND3, NW3, *, NI2
			8'd3 : rdata = 43'b0001101100000011010000000111100000000000000;
			// PEs: 35, 36 -> 32
			// srcs: (5, 4)(524) 2, (525) 6 --> (721) 8:PENB, NI0, +, PEGB0
			8'd4 : rdata = 43'b0000111011111110101000000000000000010000000;
			// PEs: 35, 36 -> 37
			// srcs: (6, 5)(602) 4, (603) 0 --> (796) 4:PENB, NI1, +, PENB
			8'd5 : rdata = 43'b0000111011111110101000000010000000100000000;
			// PEs: 36 -> 37
			// srcs: (13, 6)(604) -6 --> (604) -6:NI2, pass, PENB
			8'd6 : rdata = 43'b1100010100000010000000000000000000100000000;
			// PEs: 38, 36 -> 36
			// srcs: (235, 7)(809) 0, (46) 2 --> (852) 0:PEGB6, ND0, *, NI0
			8'd7 : rdata = 43'b0001111100001100011000000001000000000000000;
			// PEs: 36, 35 -> 35
			// srcs: (237, 11)(3) 1, (851) 0 --> (1051) 0:NM0, PENB, *, PEGB3
			8'd8 : rdata = 43'b0001110000000000110111111100000000010110000;
			// PEs: 36, 36 -> 
			// srcs: (238, 12)(3) 1, (852) 0 --> (1052) 0:NM0, NI0, *, 
			8'd9 : rdata = 43'b0001110000000000101000000000000000000000000;
			// PEs: 36, 36 -> 36
			// srcs: (241, 17)(247) 2, (1052) 0 --> (1252) 2:NW0, ALU, -, NW0
			8'd10 : rdata = 43'b0001001000000000001111111110001000000000000;
			// PEs: 38, 36 -> 
			// srcs: (313, 8)(809) 0, (124) -3 --> (930) 0:PEGB6, ND1, *, 
			8'd11 : rdata = 43'b0001111100001100011000000010000000000000000;
			// PEs: 36, 36 -> 
			// srcs: (316, 13)(3) 1, (930) 0 --> (1130) 0:NM0, ALU, *, 
			8'd12 : rdata = 43'b0001110000000000001111111110000000000000000;
			// PEs: 36, 36 -> 36
			// srcs: (319, 18)(325) -2, (1130) 0 --> (1330) -2:NW1, ALU, -, NW1
			8'd13 : rdata = 43'b0001001000000001001111111110001010000000000;
			// PEs: 38, 36 -> 36
			// srcs: (391, 9)(809) 0, (202) 0 --> (1008) 0:PEGB6, ND2, *, NI0
			8'd14 : rdata = 43'b0001111100001100011000000101000000000000000;
			// PEs: 38, 36 -> 36
			// srcs: (392, 10)(809) 0, (203) 2 --> (1009) 0:PEGB6, ND3, *, NI1
			8'd15 : rdata = 43'b0001111100001100011000000111010000000000000;
			// PEs: 36, 35 -> 35
			// srcs: (393, 14)(3) 1, (1007) 0 --> (1207) 0:NM0, PENB, *, PEGB3
			8'd16 : rdata = 43'b0001110000000000110111111100000000010110000;
			// PEs: 36, 36 -> 36
			// srcs: (394, 15)(3) 1, (1008) 0 --> (1208) 0:NM0, NI0, *, NI2
			8'd17 : rdata = 43'b0001110000000000101000000001100000000000000;
			// PEs: 36, 36 -> 36
			// srcs: (395, 16)(3) 1, (1009) 0 --> (1209) 0:NM0, NI1, *, NI0
			8'd18 : rdata = 43'b0001110000000000101000000011000000000000000;
			// PEs: 36, 36 -> 36
			// srcs: (397, 19)(403) 1, (1208) 0 --> (1408) 1:NW2, NI2, -, NW2
			8'd19 : rdata = 43'b0001001000000010101000000100001100000000000;
			// PEs: 36, 36 -> 36
			// srcs: (398, 20)(404) -3, (1209) 0 --> (1409) -3:NW3, NI0, -, NW3
			8'd20 : rdata = 43'b0001001000000011101000000000001110000000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 37) begin
	always @(*) begin
		case(address)
			// PEs: 37, 37 -> 38
			// srcs: (1, 0)(48) -3, (249) 1 --> (449) -3:ND0, NW0, *, PENB
			8'd0 : rdata = 43'b0001101100000000010000000000000000100000000;
			// PEs: 37, 37 -> 38
			// srcs: (2, 1)(126) -3, (327) 2 --> (527) -6:ND1, NW1, *, PENB
			8'd1 : rdata = 43'b0001101100000001010000000010000000100000000;
			// PEs: 37, 37 -> 32
			// srcs: (3, 2)(10) -3, (211) -2 --> (411) 6:ND2, NW2, *, PEGB0
			8'd2 : rdata = 43'b0001101100000010010000000100000000010000000;
			// PEs: 37, 37 -> 37
			// srcs: (4, 3)(805) 0, (204) -1 --> (806) 1:NM0, ND3, -, NI0
			8'd3 : rdata = 43'b0001010000000000011000000111000000000000000;
			// PEs: 36 -> 
			// srcs: (8, 4)(796) 4 --> (796) 4:PENB, pass, 
			8'd4 : rdata = 43'b1100011011111110000000000000000000000000000;
			// PEs: 37, 36 -> 39
			// srcs: (15, 5)(796) 4, (604) -6 --> (797) -2:ALU, PENB, +, PEGB7
			8'd5 : rdata = 43'b0000100111111111110111111100000000011110000;
			// PEs: 34 -> 
			// srcs: (99, 6)(793) -7 --> (793) -7:PEGB2, pass, 
			8'd6 : rdata = 43'b1100011100000100000000000000000000000000000;
			// PEs: 37, 39 -> 33
			// srcs: (102, 7)(793) -7, (798) 0 --> (799) -7:ALU, PEGB7, +, PEGB1
			8'd7 : rdata = 43'b0000100111111111111000011100000000010010000;
			// PEs: 37, 32 -> 38
			// srcs: (176, 8)(204) -1, (803) 92 --> (804) -92:ND3, PEGB0, *, PENB
			8'd8 : rdata = 43'b0001101100000011111000000000000000100000000;
			// PEs: 37 -> 38
			// srcs: (184, 9)(806) 1 --> (806) 1:NI0, pass, PENB
			8'd9 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 38, 37 -> 
			// srcs: (200, 10)(809) 0, (10) -3 --> (816) 0:PEGB6, ND2, *, 
			8'd10 : rdata = 43'b0001111100001100011000000100000000000000000;
			// PEs: 37, 37 -> 
			// srcs: (203, 13)(3) 1, (816) 0 --> (1016) 0:NM1, ALU, *, 
			8'd11 : rdata = 43'b0001110000000001001111111110000000000000000;
			// PEs: 37, 37 -> 37
			// srcs: (206, 16)(211) -2, (1016) 0 --> (1216) -2:NW2, ALU, -, NW2
			8'd12 : rdata = 43'b0001001000000010001111111110001100000000000;
			// PEs: 38, 37 -> 
			// srcs: (237, 11)(809) 0, (48) -3 --> (854) 0:PEGB6, ND0, *, 
			8'd13 : rdata = 43'b0001111100001100011000000000000000000000000;
			// PEs: 37, 37 -> 
			// srcs: (240, 14)(3) 1, (854) 0 --> (1054) 0:NM1, ALU, *, 
			8'd14 : rdata = 43'b0001110000000001001111111110000000000000000;
			// PEs: 37, 37 -> 37
			// srcs: (243, 17)(249) 1, (1054) 0 --> (1254) 1:NW0, ALU, -, NW0
			8'd15 : rdata = 43'b0001001000000000001111111110001000000000000;
			// PEs: 38, 37 -> 
			// srcs: (315, 12)(809) 0, (126) -3 --> (932) 0:PEGB6, ND1, *, 
			8'd16 : rdata = 43'b0001111100001100011000000010000000000000000;
			// PEs: 37, 37 -> 
			// srcs: (318, 15)(3) 1, (932) 0 --> (1132) 0:NM1, ALU, *, 
			8'd17 : rdata = 43'b0001110000000001001111111110000000000000000;
			// PEs: 37, 37 -> 37
			// srcs: (321, 18)(327) 2, (1132) 0 --> (1332) 2:NW1, ALU, -, NW1
			8'd18 : rdata = 43'b0001001000000001001111111110001010000000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 38) begin
	always @(*) begin
		case(address)
			// PEs: 38, 38 -> 38
			// srcs: (1, 0)(49) 1, (250) -2 --> (450) -2:ND0, NW0, *, NI0
			8'd0 : rdata = 43'b0001101100000000010000000001000000000000000;
			// PEs: 38, 38 -> 38
			// srcs: (2, 1)(127) -3, (328) -3 --> (528) 9:ND1, NW1, *, NI1
			8'd1 : rdata = 43'b0001101100000001010000000011010000000000000;
			// PEs: 38, 38 -> 33
			// srcs: (3, 2)(13) 2, (214) 0 --> (414) 0:ND2, NW2, *, PEGB1
			8'd2 : rdata = 43'b0001101100000010010000000100000000010010000;
			// PEs: 37, 38 -> 32
			// srcs: (4, 5)(449) -3, (450) -2 --> (646) -5:PENB, NI0, +, PEGB0
			8'd3 : rdata = 43'b0000111011111110101000000000000000010000000;
			// PEs: 37, 38 -> 33
			// srcs: (5, 6)(527) -6, (528) 9 --> (723) 3:PENB, NI1, +, PEGB1
			8'd4 : rdata = 43'b0000111011111110101000000010000000010010000;
			// PEs: 34 -> 
			// srcs: (6, 3)(444) 2 --> (444) 2:PEGB2, pass, 
			8'd5 : rdata = 43'b1100011100000100000000000000000000000000000;
			// PEs: 33, 38 -> 32
			// srcs: (9, 4)(443) 6, (444) 2 --> (641) 8:PEGB1, ALU, +, PEGB0
			8'd6 : rdata = 43'b0000111100000010001111111110000000010000000;
			// PEs: 37, 38 -> 
			// srcs: (179, 7)(804) -92, (807) 1 --> (808) 0:PENB, NM0, >, 
			8'd7 : rdata = 43'b0011111011111110100000000000000000000000000;
			// PEs: 38, 37 -> 39, 32, 38
			// srcs: (186, 8)(808) 0, (806) 1 --> (809) 0:ALU, PENB, *, NI0, PENB, PEGB0
			8'd8 : rdata = 43'b0001100111111111110111111101000000110000000;
			// PEs: 38 -> 32
			// srcs: (188, 9)(809) 0 --> (809) 0:ALU, pass, PEGB0
			8'd9 : rdata = 43'b1100000111111111000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (189, 10)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd10 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (190, 11)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd11 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (191, 12)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd12 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (192, 13)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd13 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 37
			// srcs: (193, 14)(809) 0 --> (809) 0:NI0, pass, PEGB5
			8'd14 : rdata = 43'b1100010100000000000000000000000000011010000;
			// PEs: 38 -> 32
			// srcs: (194, 15)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd15 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (195, 16)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd16 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38, 38 -> 39
			// srcs: (196, 17)(809) 0, (13) 2 --> (819) 0:NI0, ND2, *, PENB
			8'd17 : rdata = 43'b0001110100000000011000000100000000100000000;
			// PEs: 38 -> 32
			// srcs: (197, 18)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd18 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (198, 19)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd19 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (199, 20)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd20 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (200, 21)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd21 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (201, 22)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd22 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (202, 23)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd23 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (203, 24)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd24 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (204, 25)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd25 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (205, 26)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd26 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (206, 27)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd27 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (207, 28)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd28 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (208, 29)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd29 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (209, 30)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd30 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (210, 31)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd31 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (211, 32)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd32 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (212, 33)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd33 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (213, 34)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd34 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (214, 35)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd35 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (215, 36)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd36 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (216, 37)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd37 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (217, 38)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd38 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (218, 39)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd39 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (219, 40)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd40 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (220, 41)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd41 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (221, 42)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd42 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (222, 43)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd43 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (223, 44)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd44 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 33
			// srcs: (224, 45)(809) 0 --> (809) 0:NI0, pass, PEGB1
			8'd45 : rdata = 43'b1100010100000000000000000000000000010010000;
			// PEs: 38 -> 34
			// srcs: (225, 46)(809) 0 --> (809) 0:NI0, pass, PEGB2
			8'd46 : rdata = 43'b1100010100000000000000000000000000010100000;
			// PEs: 38 -> 32
			// srcs: (226, 47)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd47 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 35
			// srcs: (227, 48)(809) 0 --> (809) 0:NI0, pass, PEGB3
			8'd48 : rdata = 43'b1100010100000000000000000000000000010110000;
			// PEs: 38 -> 36
			// srcs: (228, 49)(809) 0 --> (809) 0:NI0, pass, PEGB4
			8'd49 : rdata = 43'b1100010100000000000000000000000000011000000;
			// PEs: 38 -> 32
			// srcs: (229, 50)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd50 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 37
			// srcs: (230, 51)(809) 0 --> (809) 0:NI0, pass, PEGB5
			8'd51 : rdata = 43'b1100010100000000000000000000000000011010000;
			// PEs: 38, 38 -> 39
			// srcs: (231, 52)(809) 0, (49) 1 --> (855) 0:NI0, ND0, *, PENB
			8'd52 : rdata = 43'b0001110100000000011000000000000000100000000;
			// PEs: 38 -> 32
			// srcs: (232, 53)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd53 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 39
			// srcs: (233, 54)(809) 0 --> (809) 0:NI0, pass, PENB
			8'd54 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 38 -> 32
			// srcs: (234, 55)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd55 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (235, 56)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd56 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (236, 57)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd57 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (237, 58)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd58 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (238, 59)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd59 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (239, 60)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd60 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (240, 61)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd61 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (241, 62)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd62 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (242, 63)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd63 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (243, 64)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd64 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (244, 65)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd65 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (245, 66)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd66 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (246, 67)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd67 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (247, 68)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd68 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (248, 69)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd69 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (249, 70)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd70 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (250, 71)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd71 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (251, 72)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd72 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (252, 73)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd73 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (253, 74)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd74 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (254, 75)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd75 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (255, 76)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd76 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (256, 77)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd77 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (257, 78)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd78 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (258, 79)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd79 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (259, 80)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd80 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (260, 81)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd81 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (261, 82)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd82 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (262, 83)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd83 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (263, 84)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd84 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (264, 85)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd85 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (265, 86)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd86 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (266, 87)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd87 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (267, 88)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd88 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (268, 89)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd89 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (269, 90)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd90 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (270, 91)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd91 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (271, 92)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd92 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (272, 93)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd93 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (273, 94)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd94 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (274, 95)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd95 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (275, 96)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd96 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (276, 97)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd97 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (277, 98)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd98 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (278, 99)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd99 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (279, 100)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd100 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (280, 101)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd101 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (281, 102)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd102 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (282, 103)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd103 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (283, 104)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd104 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (284, 105)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd105 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (285, 106)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd106 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (286, 107)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd107 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (287, 108)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd108 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (288, 109)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd109 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (289, 110)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd110 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (290, 111)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd111 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (291, 112)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd112 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (292, 113)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd113 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (293, 114)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd114 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (294, 115)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd115 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (295, 116)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd116 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (296, 117)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd117 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (297, 118)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd118 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (298, 119)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd119 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (299, 120)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd120 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (300, 121)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd121 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (301, 122)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd122 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 33
			// srcs: (302, 123)(809) 0 --> (809) 0:NI0, pass, PEGB1
			8'd123 : rdata = 43'b1100010100000000000000000000000000010010000;
			// PEs: 38 -> 34
			// srcs: (303, 124)(809) 0 --> (809) 0:NI0, pass, PEGB2
			8'd124 : rdata = 43'b1100010100000000000000000000000000010100000;
			// PEs: 38 -> 32
			// srcs: (304, 125)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd125 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 35
			// srcs: (305, 126)(809) 0 --> (809) 0:NI0, pass, PEGB3
			8'd126 : rdata = 43'b1100010100000000000000000000000000010110000;
			// PEs: 38 -> 36
			// srcs: (306, 127)(809) 0 --> (809) 0:NI0, pass, PEGB4
			8'd127 : rdata = 43'b1100010100000000000000000000000000011000000;
			// PEs: 38 -> 32
			// srcs: (307, 128)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd128 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 37
			// srcs: (308, 129)(809) 0 --> (809) 0:NI0, pass, PEGB5
			8'd129 : rdata = 43'b1100010100000000000000000000000000011010000;
			// PEs: 38, 38 -> 39
			// srcs: (309, 130)(809) 0, (127) -3 --> (933) 0:NI0, ND1, *, PENB
			8'd130 : rdata = 43'b0001110100000000011000000010000000100000000;
			// PEs: 38 -> 32
			// srcs: (310, 131)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd131 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 39
			// srcs: (311, 132)(809) 0 --> (809) 0:NI0, pass, PENB
			8'd132 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 38 -> 32
			// srcs: (312, 133)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd133 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (313, 134)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd134 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (314, 135)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd135 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (315, 136)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd136 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (316, 137)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd137 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (317, 138)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd138 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (318, 139)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd139 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (319, 140)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd140 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (320, 141)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd141 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (321, 142)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd142 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (322, 143)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd143 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (323, 144)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd144 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (324, 145)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd145 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (325, 146)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd146 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (326, 147)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd147 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (327, 148)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd148 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (328, 149)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd149 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (329, 150)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd150 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (330, 151)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd151 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (331, 152)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd152 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (332, 153)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd153 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (333, 154)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd154 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (334, 155)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd155 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (335, 156)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd156 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (336, 157)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd157 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (337, 158)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd158 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (338, 159)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd159 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (339, 160)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd160 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (340, 161)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd161 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (341, 162)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd162 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (342, 163)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd163 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (343, 164)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd164 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (344, 165)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd165 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (345, 166)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd166 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (346, 167)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd167 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (347, 168)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd168 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (348, 169)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd169 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (349, 170)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd170 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (350, 171)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd171 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (351, 172)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd172 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (352, 173)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd173 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (353, 174)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd174 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (354, 175)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd175 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (355, 176)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd176 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (356, 177)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd177 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (357, 178)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd178 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (358, 179)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd179 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (359, 180)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd180 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (360, 181)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd181 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (361, 182)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd182 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (362, 183)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd183 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (363, 184)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd184 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (364, 185)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd185 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (365, 186)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd186 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (366, 187)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd187 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (367, 188)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd188 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (368, 189)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd189 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (369, 190)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd190 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (370, 191)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd191 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (371, 192)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd192 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (372, 193)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd193 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (373, 194)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd194 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (374, 195)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd195 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (375, 196)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd196 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 33
			// srcs: (376, 197)(809) 0 --> (809) 0:NI0, pass, PEGB1
			8'd197 : rdata = 43'b1100010100000000000000000000000000010010000;
			// PEs: 38 -> 32
			// srcs: (377, 198)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd198 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 32
			// srcs: (378, 199)(809) 0 --> (809) 0:NI0, pass, PEGB0
			8'd199 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 38 -> 34
			// srcs: (379, 200)(809) 0 --> (809) 0:NI0, pass, PEGB2
			8'd200 : rdata = 43'b1100010100000000000000000000000000010100000;
			// PEs: 38 -> 33
			// srcs: (380, 201)(809) 0 --> (809) 0:NI0, pass, PEGB1
			8'd201 : rdata = 43'b1100010100000000000000000000000000010010000;
			// PEs: 38 -> 34
			// srcs: (381, 202)(809) 0 --> (809) 0:NI0, pass, PEGB2
			8'd202 : rdata = 43'b1100010100000000000000000000000000010100000;
			// PEs: 38 -> 35
			// srcs: (382, 203)(809) 0 --> (809) 0:NI0, pass, PEGB3
			8'd203 : rdata = 43'b1100010100000000000000000000000000010110000;
			// PEs: 38 -> 35
			// srcs: (383, 204)(809) 0 --> (809) 0:NI0, pass, PEGB3
			8'd204 : rdata = 43'b1100010100000000000000000000000000010110000;
			// PEs: 38 -> 36
			// srcs: (384, 205)(809) 0 --> (809) 0:NI0, pass, PEGB4
			8'd205 : rdata = 43'b1100010100000000000000000000000000011000000;
			// PEs: 38 -> 36
			// srcs: (385, 206)(809) 0 --> (809) 0:NI0, pass, PEGB4
			8'd206 : rdata = 43'b1100010100000000000000000000000000011000000;
			// PEs: 38, 39 -> 38
			// srcs: (386, 207)(214) 0, (1019) 0 --> (1219) 0:NW2, PEGB7, -, NW2
			8'd207 : rdata = 43'b0001001000000010111000011100001100000000000;
			// PEs: 38, 39 -> 38
			// srcs: (387, 208)(250) -2, (1055) 0 --> (1255) -2:NW0, PEGB7, -, NW0
			8'd208 : rdata = 43'b0001001000000000111000011100001000000000000;
			// PEs: 38, 39 -> 38
			// srcs: (388, 209)(328) -3, (1133) 0 --> (1333) -3:NW1, PEGB7, -, NW1
			8'd209 : rdata = 43'b0001001000000001111000011100001010000000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 39) begin
	always @(*) begin
		case(address)
			// PEs: 39, 39 -> 32
			// srcs: (1, 0)(51) 2, (252) -2 --> (452) -4:ND0, NW0, *, PENB
			8'd0 : rdata = 43'b0001101100000000010000000000000000100000000;
			// PEs: 39, 39 -> 32
			// srcs: (2, 1)(129) 1, (330) 1 --> (530) 1:ND1, NW1, *, PENB
			8'd1 : rdata = 43'b0001101100000001010000000010000000100000000;
			// PEs: 39, 39 -> 32
			// srcs: (3, 2)(16) -3, (217) 2 --> (417) -6:ND2, NW2, *, PENB
			8'd2 : rdata = 43'b0001101100000010010000000100000000100000000;
			// PEs: 36 -> 
			// srcs: (6, 3)(447) 4 --> (447) 4:PEGB4, pass, 
			8'd3 : rdata = 43'b1100011100001000000000000000000000000000000;
			// PEs: 35, 39 -> 32
			// srcs: (9, 4)(446) 0, (447) 4 --> (643) 4:PEGB3, ALU, +, PENB
			8'd4 : rdata = 43'b0000111100000110001111111110000000100000000;
			// PEs: 37 -> 
			// srcs: (20, 5)(797) -2 --> (797) -2:PEGB5, pass, 
			8'd5 : rdata = 43'b1100011100001010000000000000000000000000000;
			// PEs: 35, 39 -> 37
			// srcs: (23, 6)(795) 2, (797) -2 --> (798) 0:PEGB3, ALU, +, PEGB5
			8'd6 : rdata = 43'b0000111100000110001111111110000000011010000;
			// PEs: 38, 39 -> 
			// srcs: (189, 7)(809) 0, (16) -3 --> (822) 0:PENB, ND2, *, 
			8'd7 : rdata = 43'b0001111011111110011000000100000000000000000;
			// PEs: 39, 39 -> 
			// srcs: (192, 11)(3) 1, (822) 0 --> (1022) 0:NM0, ALU, *, 
			8'd8 : rdata = 43'b0001110000000000001111111110000000000000000;
			// PEs: 39, 39 -> 39
			// srcs: (195, 16)(217) 2, (1022) 0 --> (1222) 2:NW2, ALU, -, NW2
			8'd9 : rdata = 43'b0001001000000010001111111110001100000000000;
			// PEs: 39, 38 -> 38
			// srcs: (199, 10)(3) 1, (819) 0 --> (1019) 0:NM0, PENB, *, PEGB6
			8'd10 : rdata = 43'b0001110000000000110111111100000000011100000;
			// PEs: 39, 38 -> 38
			// srcs: (234, 12)(3) 1, (855) 0 --> (1055) 0:NM0, PENB, *, PEGB6
			8'd11 : rdata = 43'b0001110000000000110111111100000000011100000;
			// PEs: 38, 39 -> 
			// srcs: (237, 8)(809) 0, (51) 2 --> (857) 0:PENB, ND0, *, 
			8'd12 : rdata = 43'b0001111011111110011000000000000000000000000;
			// PEs: 39, 39 -> 
			// srcs: (240, 13)(3) 1, (857) 0 --> (1057) 0:NM0, ALU, *, 
			8'd13 : rdata = 43'b0001110000000000001111111110000000000000000;
			// PEs: 39, 39 -> 39
			// srcs: (243, 17)(252) -2, (1057) 0 --> (1257) -2:NW0, ALU, -, NW0
			8'd14 : rdata = 43'b0001001000000000001111111110001000000000000;
			// PEs: 39, 38 -> 38
			// srcs: (312, 14)(3) 1, (933) 0 --> (1133) 0:NM0, PENB, *, PEGB6
			8'd15 : rdata = 43'b0001110000000000110111111100000000011100000;
			// PEs: 38, 39 -> 
			// srcs: (315, 9)(809) 0, (129) 1 --> (935) 0:PENB, ND1, *, 
			8'd16 : rdata = 43'b0001111011111110011000000010000000000000000;
			// PEs: 39, 39 -> 
			// srcs: (318, 15)(3) 1, (935) 0 --> (1135) 0:NM0, ALU, *, 
			8'd17 : rdata = 43'b0001110000000000001111111110000000000000000;
			// PEs: 39, 39 -> 39
			// srcs: (321, 18)(330) 1, (1135) 0 --> (1335) 1:NW1, ALU, -, NW1
			8'd18 : rdata = 43'b0001001000000001001111111110001010000000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 40) begin
	always @(*) begin
		case(address)
			// PEs: 32 -> 41
			// srcs: (5, 0)(452) -4 --> (452) -4:PUNB, pass, PENB
			8'd0 : rdata = 43'b1100011011111111000000000000000000100000000;
			// PEs: 32 -> 41
			// srcs: (6, 1)(530) 1 --> (530) 1:PUNB, pass, PENB
			8'd1 : rdata = 43'b1100011011111111000000000000000000100000000;
			// PEs: 41 -> 32
			// srcs: (8, 2)(420) 3 --> (420) 3:PEGB1, pass, PUGB4
			8'd2 : rdata = 43'b1100011100000010000000000000000000000001100;
			// PEs: 43 -> 48
			// srcs: (9, 4)(426) -3 --> (426) -3:PEGB3, pass, PUNB
			8'd3 : rdata = 43'b1100011100000110000000000000000001000000000;
			// PEs: 44 -> 56
			// srcs: (10, 5)(429) 1 --> (429) 1:PEGB4, pass, PUGB7
			8'd4 : rdata = 43'b1100011100001000000000000000000000000001111;
			// PEs: 45 -> 0
			// srcs: (11, 6)(436) -1 --> (436) -1:PEGB5, pass, PUGB0
			8'd5 : rdata = 43'b1100011100001010000000000000000000000001000;
			// PEs: 46 -> 8
			// srcs: (12, 7)(439) 0 --> (439) 0:PEGB6, pass, PUGB1
			8'd6 : rdata = 43'b1100011100001100000000000000000000000001001;
			// PEs: 47 -> 32
			// srcs: (13, 8)(442) 0 --> (442) 0:PENB, pass, PUGB4
			8'd7 : rdata = 43'b1100011011111110000000000000000000000001100;
			// PEs: 41 -> 48
			// srcs: (14, 12)(648) -5 --> (648) -5:PEGB1, pass, PUNB
			8'd8 : rdata = 43'b1100011100000010000000000000000001000000000;
			// PEs: 47 -> 48
			// srcs: (15, 13)(657) -4 --> (657) -4:PENB, pass, PUNB
			8'd9 : rdata = 43'b1100011011111110000000000000000001000000000;
			// PEs: 47 -> 8
			// srcs: (16, 18)(734) -2 --> (734) -2:PENB, pass, PUGB1
			8'd10 : rdata = 43'b1100011011111110000000000000000000000001001;
			// PEs: 8 -> 41
			// srcs: (20, 3)(619) -2 --> (619) -2:PUGB1, pass, PENB
			8'd11 : rdata = 43'b1100011100000011000000000000000000100000000;
			// PEs: 32 -> 40
			// srcs: (21, 9)(646) -5 --> (646) -5:PUNB, pass, NI0
			8'd12 : rdata = 43'b1100011011111111000000000001000000000000000;
			// PEs: 48 -> 41
			// srcs: (22, 10)(451) -4 --> (451) -4:PUGB6, pass, PENB
			8'd13 : rdata = 43'b1100011100001101000000000000000000100000000;
			// PEs: 40 -> 41
			// srcs: (28, 11)(646) -5 --> (646) -5:NI0, pass, PENB
			8'd14 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 16 -> 40
			// srcs: (29, 14)(697) -1 --> (697) -1:PUGB2, pass, NI0
			8'd15 : rdata = 43'b1100011100000101000000000001000000000000000;
			// PEs: 0 -> 41
			// srcs: (30, 15)(504) 2 --> (504) 2:PUGB0, pass, PENB
			8'd16 : rdata = 43'b1100011100000001000000000000000000100000000;
			// PEs: 41 -> 48
			// srcs: (35, 26)(647) -9 --> (647) -9:PEGB1, pass, PUNB
			8'd17 : rdata = 43'b1100011100000010000000000000000001000000000;
			// PEs: 40 -> 41
			// srcs: (36, 16)(697) -1 --> (697) -1:NI0, pass, PENB
			8'd18 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 8 -> 41
			// srcs: (37, 17)(536) 0 --> (536) 0:PUGB1, pass, PENB
			8'd19 : rdata = 43'b1100011100000011000000000000000000100000000;
			// PEs: 56 -> 40
			// srcs: (38, 19)(747) 7 --> (747) 7:PUGB7, pass, NI0
			8'd20 : rdata = 43'b1100011100001111000000000001000000000000000;
			// PEs: 16 -> 41
			// srcs: (39, 20)(554) 0 --> (554) 0:PUGB2, pass, PENB
			8'd21 : rdata = 43'b1100011100000101000000000000000000100000000;
			// PEs: 42 -> 48
			// srcs: (40, 27)(656) 11 --> (656) 11:PEGB2, pass, PUNB
			8'd22 : rdata = 43'b1100011100000100000000000000000001000000000;
			// PEs: 41 -> 16
			// srcs: (43, 28)(698) 1 --> (698) 1:PEGB1, pass, PUGB2
			8'd23 : rdata = 43'b1100011100000010000000000000000000000001010;
			// PEs: 40 -> 41
			// srcs: (45, 21)(747) 7 --> (747) 7:NI0, pass, PENB
			8'd24 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 32 -> 40
			// srcs: (46, 22)(612) -3 --> (612) -3:PUNB, pass, NI0
			8'd25 : rdata = 43'b1100011011111111000000000001000000000000000;
			// PEs: 16 -> 41
			// srcs: (47, 23)(614) -2 --> (614) -2:PUGB2, pass, PENB
			8'd26 : rdata = 43'b1100011100000101000000000000000000100000000;
			// PEs: 32 -> 46
			// srcs: (48, 25)(618) 2 --> (618) 2:PUNB, pass, PEGB6
			8'd27 : rdata = 43'b1100011011111111000000000000000000011100000;
			// PEs: 41 -> 48
			// srcs: (52, 32)(748) 7 --> (748) 7:PEGB1, pass, PUNB
			8'd28 : rdata = 43'b1100011100000010000000000000000001000000000;
			// PEs: 40 -> 41
			// srcs: (53, 24)(612) -3 --> (612) -3:NI0, pass, PENB
			8'd29 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 44 -> 48
			// srcs: (54, 36)(733) 5 --> (733) 5:PEGB4, pass, PUNB
			8'd30 : rdata = 43'b1100011100001000000000000000000001000000000;
			// PEs: 16 -> 40
			// srcs: (57, 29)(717) 10 --> (717) 10:PUGB2, pass, NI0
			8'd31 : rdata = 43'b1100011100000101000000000001000000000000000;
			// PEs: 32 -> 41
			// srcs: (58, 30)(719) 5 --> (719) 5:PUNB, pass, PENB
			8'd32 : rdata = 43'b1100011011111111000000000000000000100000000;
			// PEs: 46 -> 56
			// srcs: (60, 34)(621) 4 --> (621) 4:PEGB6, pass, PUGB7
			8'd33 : rdata = 43'b1100011100001100000000000000000000000001111;
			// PEs: 40 -> 41
			// srcs: (64, 31)(717) 10 --> (717) 10:NI0, pass, PENB
			8'd34 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 48 -> 41
			// srcs: (65, 33)(610) 0 --> (610) 0:PUGB6, pass, PENB
			8'd35 : rdata = 43'b1100011100001101000000000000000000100000000;
			// PEs: 41 -> 8
			// srcs: (72, 37)(616) -5 --> (616) -5:PEGB1, pass, PUGB1
			8'd36 : rdata = 43'b1100011100000010000000000000000000000001001;
			// PEs: 32 -> 41
			// srcs: (91, 35)(725) 3 --> (725) 3:PUNB, pass, PENB
			8'd37 : rdata = 43'b1100011011111111000000000000000000100000000;
			// PEs: 56 -> 41
			// srcs: (92, 38)(715) 9 --> (715) 9:PUGB7, pass, PENB
			8'd38 : rdata = 43'b1100011100001111000000000000000000100000000;
			// PEs: 56 -> 41
			// srcs: (126, 39)(751) 29 --> (751) 29:PUGB7, pass, PENB
			8'd39 : rdata = 43'b1100011100001111000000000000000000100000000;
			// PEs: 41 -> 48
			// srcs: (134, 40)(752) 56 --> (752) 56:PEGB1, pass, PUNB
			8'd40 : rdata = 43'b1100011100000010000000000000000001000000000;
			// PEs: 32 -> 41
			// srcs: (210, 41)(809) 0 --> (809) 0:PUNB, pass, PENB
			8'd41 : rdata = 43'b1100011011111111000000000000000000100000000;
			// PEs: 32 -> 42
			// srcs: (213, 42)(809) 0 --> (809) 0:PUNB, pass, PEGB2
			8'd42 : rdata = 43'b1100011011111111000000000000000000010100000;
			// PEs: 32 -> 43
			// srcs: (216, 43)(809) 0 --> (809) 0:PUNB, pass, PEGB3
			8'd43 : rdata = 43'b1100011011111111000000000000000000010110000;
			// PEs: 32 -> 44
			// srcs: (219, 44)(809) 0 --> (809) 0:PUNB, pass, PEGB4
			8'd44 : rdata = 43'b1100011011111111000000000000000000011000000;
			// PEs: 32 -> 45
			// srcs: (226, 45)(809) 0 --> (809) 0:PUNB, pass, PEGB5
			8'd45 : rdata = 43'b1100011011111111000000000000000000011010000;
			// PEs: 32 -> 46
			// srcs: (229, 46)(809) 0 --> (809) 0:PUNB, pass, PEGB6
			8'd46 : rdata = 43'b1100011011111111000000000000000000011100000;
			// PEs: 32 -> 47
			// srcs: (232, 47)(809) 0 --> (809) 0:PUNB, pass, PEGB7
			8'd47 : rdata = 43'b1100011011111111000000000000000000011110000;
			// PEs: 32 -> 41
			// srcs: (243, 48)(809) 0 --> (809) 0:PUNB, pass, PENB
			8'd48 : rdata = 43'b1100011011111111000000000000000000100000000;
			// PEs: 32 -> 42
			// srcs: (245, 49)(809) 0 --> (809) 0:PUNB, pass, PEGB2
			8'd49 : rdata = 43'b1100011011111111000000000000000000010100000;
			// PEs: 32 -> 43
			// srcs: (246, 50)(809) 0 --> (809) 0:PUNB, pass, PEGB3
			8'd50 : rdata = 43'b1100011011111111000000000000000000010110000;
			// PEs: 32 -> 44
			// srcs: (247, 51)(809) 0 --> (809) 0:PUNB, pass, PEGB4
			8'd51 : rdata = 43'b1100011011111111000000000000000000011000000;
			// PEs: 32 -> 45
			// srcs: (248, 52)(809) 0 --> (809) 0:PUNB, pass, PEGB5
			8'd52 : rdata = 43'b1100011011111111000000000000000000011010000;
			// PEs: 32 -> 46
			// srcs: (249, 53)(809) 0 --> (809) 0:PUNB, pass, PEGB6
			8'd53 : rdata = 43'b1100011011111111000000000000000000011100000;
			// PEs: 32 -> 47
			// srcs: (250, 54)(809) 0 --> (809) 0:PUNB, pass, PEGB7
			8'd54 : rdata = 43'b1100011011111111000000000000000000011110000;
			// PEs: 32 -> 41
			// srcs: (321, 55)(809) 0 --> (809) 0:PUNB, pass, PENB
			8'd55 : rdata = 43'b1100011011111111000000000000000000100000000;
			// PEs: 32 -> 42
			// srcs: (322, 56)(809) 0 --> (809) 0:PUNB, pass, PEGB2
			8'd56 : rdata = 43'b1100011011111111000000000000000000010100000;
			// PEs: 32 -> 43
			// srcs: (323, 57)(809) 0 --> (809) 0:PUNB, pass, PEGB3
			8'd57 : rdata = 43'b1100011011111111000000000000000000010110000;
			// PEs: 32 -> 44
			// srcs: (324, 58)(809) 0 --> (809) 0:PUNB, pass, PEGB4
			8'd58 : rdata = 43'b1100011011111111000000000000000000011000000;
			// PEs: 32 -> 45
			// srcs: (325, 59)(809) 0 --> (809) 0:PUNB, pass, PEGB5
			8'd59 : rdata = 43'b1100011011111111000000000000000000011010000;
			// PEs: 32 -> 46
			// srcs: (327, 60)(809) 0 --> (809) 0:PUNB, pass, PEGB6
			8'd60 : rdata = 43'b1100011011111111000000000000000000011100000;
			// PEs: 32 -> 47
			// srcs: (328, 61)(809) 0 --> (809) 0:PUNB, pass, PEGB7
			8'd61 : rdata = 43'b1100011011111111000000000000000000011110000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 41) begin
	always @(*) begin
		case(address)
			// PEs: 41, 41 -> 41
			// srcs: (1, 0)(52) 1, (253) -1 --> (453) -1:ND0, NW0, *, NI0
			8'd0 : rdata = 43'b0001101100000000010000000001000000000000000;
			// PEs: 41, 41 -> 41
			// srcs: (2, 1)(130) 2, (331) 0 --> (531) 0:ND1, NW1, *, NI1
			8'd1 : rdata = 43'b0001101100000001010000000011010000000000000;
			// PEs: 41, 41 -> 40
			// srcs: (3, 2)(19) -3, (220) -1 --> (420) 3:ND2, NW2, *, PEGB0
			8'd2 : rdata = 43'b0001101100000010010000000100000000010000000;
			// PEs: 40, 41 -> 40
			// srcs: (8, 3)(452) -4, (453) -1 --> (648) -5:PENB, NI0, +, PEGB0
			8'd3 : rdata = 43'b0000111011111110101000000000000000010000000;
			// PEs: 40, 41 -> 44
			// srcs: (9, 4)(530) 1, (531) 0 --> (728) 1:PENB, NI1, +, PEGB4
			8'd4 : rdata = 43'b0000111011111110101000000010000000011000000;
			// PEs: 40, 42 -> 46
			// srcs: (22, 5)(619) -2, (423) 4 --> (620) 2:PENB, PEGB2, +, PEGB6
			8'd5 : rdata = 43'b0000111011111110111000001000000000011100000;
			// PEs: 40 -> 
			// srcs: (24, 6)(451) -4 --> (451) -4:PENB, pass, 
			8'd6 : rdata = 43'b1100011011111110000000000000000000000000000;
			// PEs: 40, 41 -> 40
			// srcs: (30, 7)(646) -5, (451) -4 --> (647) -9:PENB, ALU, +, PEGB0
			8'd7 : rdata = 43'b0000111011111110001111111110000000010000000;
			// PEs: 40 -> 
			// srcs: (32, 8)(504) 2 --> (504) 2:PENB, pass, 
			8'd8 : rdata = 43'b1100011011111110000000000000000000000000000;
			// PEs: 40, 41 -> 40
			// srcs: (38, 9)(697) -1, (504) 2 --> (698) 1:PENB, ALU, +, PEGB0
			8'd9 : rdata = 43'b0000111011111110001111111110000000010000000;
			// PEs: 45, 40 -> 44
			// srcs: (39, 10)(731) 6, (536) 0 --> (732) 6:PEGB5, PENB, +, PEGB4
			8'd10 : rdata = 43'b0000111100001010110111111100000000011000000;
			// PEs: 40 -> 
			// srcs: (41, 11)(554) 0 --> (554) 0:PENB, pass, 
			8'd11 : rdata = 43'b1100011011111110000000000000000000000000000;
			// PEs: 40, 41 -> 40
			// srcs: (47, 12)(747) 7, (554) 0 --> (748) 7:PENB, ALU, +, PEGB0
			8'd12 : rdata = 43'b0000111011111110001111111110000000010000000;
			// PEs: 40 -> 
			// srcs: (49, 13)(614) -2 --> (614) -2:PENB, pass, 
			8'd13 : rdata = 43'b1100011011111110000000000000000000000000000;
			// PEs: 40, 41 -> 41
			// srcs: (55, 14)(612) -3, (614) -2 --> (615) -5:PENB, ALU, +, NI0
			8'd14 : rdata = 43'b0000111011111110001111111111000000000000000;
			// PEs: 40 -> 
			// srcs: (60, 15)(719) 5 --> (719) 5:PENB, pass, 
			8'd15 : rdata = 43'b1100011011111110000000000000000000000000000;
			// PEs: 40, 41 -> 41
			// srcs: (66, 16)(717) 10, (719) 5 --> (720) 15:PENB, ALU, +, NI1
			8'd16 : rdata = 43'b0000111011111110001111111111010000000000000;
			// PEs: 40, 41 -> 40
			// srcs: (67, 17)(610) 0, (615) -5 --> (616) -5:PENB, NI0, +, PEGB0
			8'd17 : rdata = 43'b0000111011111110101000000000000000010000000;
			// PEs: 41, 40 -> 
			// srcs: (94, 18)(720) 15, (725) 3 --> (726) 18:NI1, PENB, +, 
			8'd18 : rdata = 43'b0000110100000001110111111100000000000000000;
			// PEs: 40, 41 -> 
			// srcs: (107, 19)(715) 9, (726) 18 --> (727) 27:PENB, ALU, +, 
			8'd19 : rdata = 43'b0000111011111110001111111110000000000000000;
			// PEs: 41, 40 -> 40
			// srcs: (129, 20)(727) 27, (751) 29 --> (752) 56:ALU, PENB, +, PEGB0
			8'd20 : rdata = 43'b0000100111111111110111111100000000010000000;
			// PEs: 40, 41 -> 42
			// srcs: (212, 21)(809) 0, (19) -3 --> (825) 0:PENB, ND2, *, PENB
			8'd21 : rdata = 43'b0001111011111110011000000100000000100000000;
			// PEs: 41, 42 -> 41
			// srcs: (221, 24)(220) -1, (1025) 0 --> (1225) -1:NW2, PEGB2, -, NW2
			8'd22 : rdata = 43'b0001001000000010111000001000001100000000000;
			// PEs: 40, 41 -> 42
			// srcs: (245, 22)(809) 0, (52) 1 --> (858) 0:PENB, ND0, *, PENB
			8'd23 : rdata = 43'b0001111011111110011000000000000000100000000;
			// PEs: 41, 42 -> 41
			// srcs: (254, 25)(253) -1, (1058) 0 --> (1258) -1:NW0, PEGB2, -, NW0
			8'd24 : rdata = 43'b0001001000000000111000001000001000000000000;
			// PEs: 40, 41 -> 42
			// srcs: (323, 23)(809) 0, (130) 2 --> (936) 0:PENB, ND1, *, PENB
			8'd25 : rdata = 43'b0001111011111110011000000010000000100000000;
			// PEs: 41, 42 -> 41
			// srcs: (332, 26)(331) 0, (1136) 0 --> (1336) 0:NW1, PEGB2, -, NW1
			8'd26 : rdata = 43'b0001001000000001111000001000001010000000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 42) begin
	always @(*) begin
		case(address)
			// PEs: 42, 42 -> 43
			// srcs: (1, 0)(54) 2, (255) 1 --> (455) 2:ND0, NW0, *, PENB
			8'd0 : rdata = 43'b0001101100000000010000000000000000100000000;
			// PEs: 42, 42 -> 43
			// srcs: (2, 1)(131) 1, (332) -3 --> (532) -3:ND1, NW1, *, PENB
			8'd1 : rdata = 43'b0001101100000001010000000010000000100000000;
			// PEs: 42, 42 -> 41
			// srcs: (3, 2)(22) 2, (223) 2 --> (423) 4:ND2, NW2, *, PEGB1
			8'd2 : rdata = 43'b0001101100000010010000000100000000010010000;
			// PEs: 45 -> 
			// srcs: (9, 3)(655) 9 --> (655) 9:PEGB5, pass, 
			8'd3 : rdata = 43'b1100011100001010000000000000000000000000000;
			// PEs: 43, 42 -> 40
			// srcs: (12, 4)(654) 2, (655) 9 --> (656) 11:PEGB3, ALU, +, PEGB0
			8'd4 : rdata = 43'b0000111100000110001111111110000000010000000;
			// PEs: 42, 41 -> 41
			// srcs: (215, 8)(3) 1, (825) 0 --> (1025) 0:NM0, PENB, *, PEGB1
			8'd5 : rdata = 43'b0001110000000000110111111100000000010010000;
			// PEs: 40, 42 -> 
			// srcs: (218, 5)(809) 0, (22) 2 --> (828) 0:PEGB0, ND2, *, 
			8'd6 : rdata = 43'b0001111100000000011000000100000000000000000;
			// PEs: 42, 42 -> 
			// srcs: (221, 9)(3) 1, (828) 0 --> (1028) 0:NM0, ALU, *, 
			8'd7 : rdata = 43'b0001110000000000001111111110000000000000000;
			// PEs: 42, 42 -> 42
			// srcs: (224, 12)(223) 2, (1028) 0 --> (1228) 2:NW2, ALU, -, NW2
			8'd8 : rdata = 43'b0001001000000010001111111110001100000000000;
			// PEs: 42, 41 -> 41
			// srcs: (248, 10)(3) 1, (858) 0 --> (1058) 0:NM0, PENB, *, PEGB1
			8'd9 : rdata = 43'b0001110000000000110111111100000000010010000;
			// PEs: 40, 42 -> 43
			// srcs: (250, 6)(809) 0, (54) 2 --> (860) 0:PEGB0, ND0, *, PENB
			8'd10 : rdata = 43'b0001111100000000011000000000000000100000000;
			// PEs: 42, 43 -> 42
			// srcs: (259, 13)(255) 1, (1060) 0 --> (1260) 1:NW0, PEGB3, -, NW0
			8'd11 : rdata = 43'b0001001000000000111000001100001000000000000;
			// PEs: 42, 41 -> 41
			// srcs: (326, 11)(3) 1, (936) 0 --> (1136) 0:NM0, PENB, *, PEGB1
			8'd12 : rdata = 43'b0001110000000000110111111100000000010010000;
			// PEs: 40, 42 -> 43
			// srcs: (327, 7)(809) 0, (131) 1 --> (937) 0:PEGB0, ND1, *, PENB
			8'd13 : rdata = 43'b0001111100000000011000000010000000100000000;
			// PEs: 42, 43 -> 42
			// srcs: (336, 14)(332) -3, (1137) 0 --> (1337) -3:NW1, PEGB3, -, NW1
			8'd14 : rdata = 43'b0001001000000001111000001100001010000000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 43) begin
	always @(*) begin
		case(address)
			// PEs: 43, 43 -> 43
			// srcs: (1, 0)(55) 0, (256) -1 --> (456) 0:ND0, NW0, *, NI0
			8'd0 : rdata = 43'b0001101100000000010000000001000000000000000;
			// PEs: 43, 43 -> 43
			// srcs: (2, 1)(132) -1, (333) -1 --> (533) 1:ND1, NW1, *, NI1
			8'd1 : rdata = 43'b0001101100000001010000000011010000000000000;
			// PEs: 43, 43 -> 40
			// srcs: (3, 2)(25) 1, (226) -3 --> (426) -3:ND2, NW2, *, PEGB0
			8'd2 : rdata = 43'b0001101100000010010000000100000000010000000;
			// PEs: 42, 43 -> 42
			// srcs: (4, 3)(455) 2, (456) 0 --> (654) 2:PENB, NI0, +, PEGB2
			8'd3 : rdata = 43'b0000111011111110101000000000000000010100000;
			// PEs: 42, 43 -> 44
			// srcs: (5, 4)(532) -3, (533) 1 --> (729) -2:PENB, NI1, +, PENB
			8'd4 : rdata = 43'b0000111011111110101000000010000000100000000;
			// PEs: 40, 43 -> 
			// srcs: (221, 5)(809) 0, (25) 1 --> (831) 0:PEGB0, ND2, *, 
			8'd5 : rdata = 43'b0001111100000000011000000100000000000000000;
			// PEs: 43, 43 -> 
			// srcs: (224, 8)(3) 1, (831) 0 --> (1031) 0:NM0, ALU, *, 
			8'd6 : rdata = 43'b0001110000000000001111111110000000000000000;
			// PEs: 43, 43 -> 43
			// srcs: (227, 11)(226) -3, (1031) 0 --> (1231) -3:NW2, ALU, -, NW2
			8'd7 : rdata = 43'b0001001000000010001111111110001100000000000;
			// PEs: 40, 43 -> 44
			// srcs: (251, 6)(809) 0, (55) 0 --> (861) 0:PEGB0, ND0, *, PENB
			8'd8 : rdata = 43'b0001111100000000011000000000000000100000000;
			// PEs: 43, 42 -> 42
			// srcs: (253, 9)(3) 1, (860) 0 --> (1060) 0:NM0, PENB, *, PEGB2
			8'd9 : rdata = 43'b0001110000000000110111111100000000010100000;
			// PEs: 43, 44 -> 43
			// srcs: (260, 12)(256) -1, (1061) 0 --> (1261) -1:NW0, PEGB4, -, NW0
			8'd10 : rdata = 43'b0001001000000000111000010000001000000000000;
			// PEs: 40, 43 -> 44
			// srcs: (328, 7)(809) 0, (132) -1 --> (938) 0:PEGB0, ND1, *, PENB
			8'd11 : rdata = 43'b0001111100000000011000000010000000100000000;
			// PEs: 43, 42 -> 42
			// srcs: (330, 10)(3) 1, (937) 0 --> (1137) 0:NM0, PENB, *, PEGB2
			8'd12 : rdata = 43'b0001110000000000110111111100000000010100000;
			// PEs: 43, 44 -> 43
			// srcs: (337, 13)(333) -1, (1138) 0 --> (1338) -1:NW1, PEGB4, -, NW1
			8'd13 : rdata = 43'b0001001000000001111000010000001010000000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 44) begin
	always @(*) begin
		case(address)
			// PEs: 44, 44 -> 45
			// srcs: (1, 0)(56) -3, (257) -2 --> (457) 6:ND0, NW0, *, PENB
			8'd0 : rdata = 43'b0001101100000000010000000000000000100000000;
			// PEs: 44, 44 -> 45
			// srcs: (2, 1)(133) -3, (334) -3 --> (534) 9:ND1, NW1, *, PENB
			8'd1 : rdata = 43'b0001101100000001010000000010000000100000000;
			// PEs: 44, 44 -> 40
			// srcs: (3, 2)(28) 1, (229) 1 --> (429) 1:ND2, NW2, *, PEGB0
			8'd2 : rdata = 43'b0001101100000010010000000100000000010000000;
			// PEs: 41, 43 -> 
			// srcs: (15, 3)(728) 1, (729) -2 --> (730) -1:PEGB1, PENB, +, 
			8'd3 : rdata = 43'b0000111100000010110111111100000000000000000;
			// PEs: 44, 41 -> 40
			// srcs: (45, 4)(730) -1, (732) 6 --> (733) 5:ALU, PEGB1, +, PEGB0
			8'd4 : rdata = 43'b0000100111111111111000000100000000010000000;
			// PEs: 40, 44 -> 
			// srcs: (224, 5)(809) 0, (28) 1 --> (834) 0:PEGB0, ND2, *, 
			8'd5 : rdata = 43'b0001111100000000011000000100000000000000000;
			// PEs: 44, 44 -> 
			// srcs: (227, 8)(3) 1, (834) 0 --> (1034) 0:NM0, ALU, *, 
			8'd6 : rdata = 43'b0001110000000000001111111110000000000000000;
			// PEs: 44, 44 -> 44
			// srcs: (230, 11)(229) 1, (1034) 0 --> (1234) 1:NW2, ALU, -, NW2
			8'd7 : rdata = 43'b0001001000000010001111111110001100000000000;
			// PEs: 40, 44 -> 45
			// srcs: (252, 6)(809) 0, (56) -3 --> (862) 0:PEGB0, ND0, *, PENB
			8'd8 : rdata = 43'b0001111100000000011000000000000000100000000;
			// PEs: 44, 43 -> 43
			// srcs: (254, 9)(3) 1, (861) 0 --> (1061) 0:NM0, PENB, *, PEGB3
			8'd9 : rdata = 43'b0001110000000000110111111100000000010110000;
			// PEs: 44, 45 -> 44
			// srcs: (261, 12)(257) -2, (1062) 0 --> (1262) -2:NW0, PEGB5, -, NW0
			8'd10 : rdata = 43'b0001001000000000111000010100001000000000000;
			// PEs: 40, 44 -> 45
			// srcs: (329, 7)(809) 0, (133) -3 --> (939) 0:PEGB0, ND1, *, PENB
			8'd11 : rdata = 43'b0001111100000000011000000010000000100000000;
			// PEs: 44, 43 -> 43
			// srcs: (331, 10)(3) 1, (938) 0 --> (1138) 0:NM0, PENB, *, PEGB3
			8'd12 : rdata = 43'b0001110000000000110111111100000000010110000;
			// PEs: 44, 45 -> 44
			// srcs: (338, 13)(334) -3, (1139) 0 --> (1339) -3:NW1, PEGB5, -, NW1
			8'd13 : rdata = 43'b0001001000000001111000010100001010000000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 45) begin
	always @(*) begin
		case(address)
			// PEs: 45, 45 -> 45
			// srcs: (1, 0)(57) -1, (258) -3 --> (458) 3:ND0, NW0, *, NI0
			8'd0 : rdata = 43'b0001101100000000010000000001000000000000000;
			// PEs: 45, 45 -> 45
			// srcs: (2, 1)(134) -3, (335) 1 --> (535) -3:ND1, NW1, *, NI1
			8'd1 : rdata = 43'b0001101100000001010000000011010000000000000;
			// PEs: 45, 45 -> 40
			// srcs: (3, 2)(35) 1, (236) -1 --> (436) -1:ND2, NW2, *, PEGB0
			8'd2 : rdata = 43'b0001101100000010010000000100000000010000000;
			// PEs: 44, 45 -> 42
			// srcs: (4, 4)(457) 6, (458) 3 --> (655) 9:PENB, NI0, +, PEGB2
			8'd3 : rdata = 43'b0000111011111110101000000000000000010100000;
			// PEs: 44, 45 -> 41
			// srcs: (5, 3)(534) 9, (535) -3 --> (731) 6:PENB, NI1, +, PEGB1
			8'd4 : rdata = 43'b0000111011111110101000000010000000010010000;
			// PEs: 40, 45 -> 
			// srcs: (231, 5)(809) 0, (35) 1 --> (841) 0:PEGB0, ND2, *, 
			8'd5 : rdata = 43'b0001111100000000011000000100000000000000000;
			// PEs: 45, 45 -> 
			// srcs: (234, 8)(3) 1, (841) 0 --> (1041) 0:NM0, ALU, *, 
			8'd6 : rdata = 43'b0001110000000000001111111110000000000000000;
			// PEs: 45, 45 -> 45
			// srcs: (237, 11)(236) -1, (1041) 0 --> (1241) -1:NW2, ALU, -, NW2
			8'd7 : rdata = 43'b0001001000000010001111111110001100000000000;
			// PEs: 40, 45 -> 46
			// srcs: (253, 6)(809) 0, (57) -1 --> (863) 0:PEGB0, ND0, *, PENB
			8'd8 : rdata = 43'b0001111100000000011000000000000000100000000;
			// PEs: 45, 44 -> 44
			// srcs: (255, 9)(3) 1, (862) 0 --> (1062) 0:NM0, PENB, *, PEGB4
			8'd9 : rdata = 43'b0001110000000000110111111100000000011000000;
			// PEs: 45, 46 -> 45
			// srcs: (262, 12)(258) -3, (1063) 0 --> (1263) -3:NW0, PEGB6, -, NW0
			8'd10 : rdata = 43'b0001001000000000111000011000001000000000000;
			// PEs: 40, 45 -> 46
			// srcs: (330, 7)(809) 0, (134) -3 --> (940) 0:PEGB0, ND1, *, PENB
			8'd11 : rdata = 43'b0001111100000000011000000010000000100000000;
			// PEs: 45, 44 -> 44
			// srcs: (332, 10)(3) 1, (939) 0 --> (1139) 0:NM0, PENB, *, PEGB4
			8'd12 : rdata = 43'b0001110000000000110111111100000000011000000;
			// PEs: 45, 46 -> 45
			// srcs: (339, 13)(335) 1, (1140) 0 --> (1340) 1:NW1, PEGB6, -, NW1
			8'd13 : rdata = 43'b0001001000000001111000011000001010000000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 46) begin
	always @(*) begin
		case(address)
			// PEs: 46, 46 -> 47
			// srcs: (1, 0)(58) 1, (259) -1 --> (459) -1:ND0, NW0, *, PENB
			8'd0 : rdata = 43'b0001101100000000010000000000000000100000000;
			// PEs: 46, 46 -> 47
			// srcs: (2, 1)(136) 0, (337) 1 --> (537) 0:ND1, NW1, *, PENB
			8'd1 : rdata = 43'b0001101100000001010000000010000000100000000;
			// PEs: 46, 46 -> 40
			// srcs: (3, 2)(38) 0, (239) 0 --> (439) 0:ND2, NW2, *, PEGB0
			8'd2 : rdata = 43'b0001101100000010010000000100000000010000000;
			// PEs: 40 -> 
			// srcs: (53, 3)(618) 2 --> (618) 2:PEGB0, pass, 
			8'd3 : rdata = 43'b1100011100000000000000000000000000000000000;
			// PEs: 46, 41 -> 40
			// srcs: (55, 4)(618) 2, (620) 2 --> (621) 4:ALU, PEGB1, +, PEGB0
			8'd4 : rdata = 43'b0000100111111111111000000100000000010000000;
			// PEs: 40, 46 -> 
			// srcs: (234, 5)(809) 0, (38) 0 --> (844) 0:PEGB0, ND2, *, 
			8'd5 : rdata = 43'b0001111100000000011000000100000000000000000;
			// PEs: 46, 46 -> 
			// srcs: (237, 8)(3) 1, (844) 0 --> (1044) 0:NM0, ALU, *, 
			8'd6 : rdata = 43'b0001110000000000001111111110000000000000000;
			// PEs: 46, 46 -> 46
			// srcs: (240, 12)(239) 0, (1044) 0 --> (1244) 0:NW2, ALU, -, NW2
			8'd7 : rdata = 43'b0001001000000010001111111110001100000000000;
			// PEs: 40, 46 -> 47
			// srcs: (254, 6)(809) 0, (58) 1 --> (864) 0:PEGB0, ND0, *, PENB
			8'd8 : rdata = 43'b0001111100000000011000000000000000100000000;
			// PEs: 46, 45 -> 45
			// srcs: (256, 9)(3) 1, (863) 0 --> (1063) 0:NM0, PENB, *, PEGB5
			8'd9 : rdata = 43'b0001110000000000110111111100000000011010000;
			// PEs: 46, 47 -> 46
			// srcs: (263, 13)(259) -1, (1064) 0 --> (1264) -1:NW0, PEGB7, -, NW0
			8'd10 : rdata = 43'b0001001000000000111000011100001000000000000;
			// PEs: 40, 46 -> 46
			// srcs: (332, 7)(809) 0, (136) 0 --> (942) 0:PEGB0, ND1, *, NI0
			8'd11 : rdata = 43'b0001111100000000011000000011000000000000000;
			// PEs: 46, 45 -> 45
			// srcs: (333, 10)(3) 1, (940) 0 --> (1140) 0:NM0, PENB, *, PEGB5
			8'd12 : rdata = 43'b0001110000000000110111111100000000011010000;
			// PEs: 46, 46 -> 
			// srcs: (335, 11)(3) 1, (942) 0 --> (1142) 0:NM0, NI0, *, 
			8'd13 : rdata = 43'b0001110000000000101000000000000000000000000;
			// PEs: 46, 46 -> 46
			// srcs: (338, 14)(337) 1, (1142) 0 --> (1342) 1:NW1, ALU, -, NW1
			8'd14 : rdata = 43'b0001001000000001001111111110001010000000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 47) begin
	always @(*) begin
		case(address)
			// PEs: 47, 47 -> 47
			// srcs: (1, 0)(59) -3, (260) 1 --> (460) -3:ND0, NW0, *, NI0
			8'd0 : rdata = 43'b0001101100000000010000000001000000000000000;
			// PEs: 47, 47 -> 47
			// srcs: (2, 1)(137) -1, (338) 2 --> (538) -2:ND1, NW1, *, NI1
			8'd1 : rdata = 43'b0001101100000001010000000011010000000000000;
			// PEs: 47, 47 -> 40
			// srcs: (3, 2)(41) -2, (242) 0 --> (442) 0:ND2, NW2, *, PENB
			8'd2 : rdata = 43'b0001101100000010010000000100000000100000000;
			// PEs: 46, 47 -> 40
			// srcs: (4, 3)(459) -1, (460) -3 --> (657) -4:PENB, NI0, +, PENB
			8'd3 : rdata = 43'b0000111011111110101000000000000000100000000;
			// PEs: 46, 47 -> 40
			// srcs: (5, 4)(537) 0, (538) -2 --> (734) -2:PENB, NI1, +, PENB
			8'd4 : rdata = 43'b0000111011111110101000000010000000100000000;
			// PEs: 40, 47 -> 
			// srcs: (237, 5)(809) 0, (41) -2 --> (847) 0:PEGB0, ND2, *, 
			8'd5 : rdata = 43'b0001111100000000011000000100000000000000000;
			// PEs: 47, 47 -> 
			// srcs: (240, 8)(3) 1, (847) 0 --> (1047) 0:NM0, ALU, *, 
			8'd6 : rdata = 43'b0001110000000000001111111110000000000000000;
			// PEs: 47, 47 -> 47
			// srcs: (243, 12)(242) 0, (1047) 0 --> (1247) 0:NW2, ALU, -, NW2
			8'd7 : rdata = 43'b0001001000000010001111111110001100000000000;
			// PEs: 40, 47 -> 47
			// srcs: (255, 6)(809) 0, (59) -3 --> (865) 0:PEGB0, ND0, *, NI0
			8'd8 : rdata = 43'b0001111100000000011000000001000000000000000;
			// PEs: 47, 46 -> 46
			// srcs: (257, 9)(3) 1, (864) 0 --> (1064) 0:NM0, PENB, *, PEGB6
			8'd9 : rdata = 43'b0001110000000000110111111100000000011100000;
			// PEs: 47, 47 -> 
			// srcs: (258, 10)(3) 1, (865) 0 --> (1065) 0:NM0, NI0, *, 
			8'd10 : rdata = 43'b0001110000000000101000000000000000000000000;
			// PEs: 47, 47 -> 47
			// srcs: (261, 13)(260) 1, (1065) 0 --> (1265) 1:NW0, ALU, -, NW0
			8'd11 : rdata = 43'b0001001000000000001111111110001000000000000;
			// PEs: 40, 47 -> 
			// srcs: (333, 7)(809) 0, (137) -1 --> (943) 0:PEGB0, ND1, *, 
			8'd12 : rdata = 43'b0001111100000000011000000010000000000000000;
			// PEs: 47, 47 -> 
			// srcs: (336, 11)(3) 1, (943) 0 --> (1143) 0:NM0, ALU, *, 
			8'd13 : rdata = 43'b0001110000000000001111111110000000000000000;
			// PEs: 47, 47 -> 47
			// srcs: (339, 14)(338) 2, (1143) 0 --> (1343) 2:NW1, ALU, -, NW1
			8'd14 : rdata = 43'b0001001000000001001111111110001010000000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 48) begin
	always @(*) begin
		case(address)
			// PEs: 55 -> 56
			// srcs: (3, 0)(471) 2 --> (471) 2:PENB, pass, PUNB
			8'd0 : rdata = 43'b1100011011111110000000000000000001000000000;
			// PEs: 55 -> 56
			// srcs: (4, 1)(549) -6 --> (549) -6:PENB, pass, PUNB
			8'd1 : rdata = 43'b1100011011111110000000000000000001000000000;
			// PEs: 49 -> 16
			// srcs: (8, 8)(445) 4 --> (445) 4:PEGB1, pass, PUGB2
			8'd2 : rdata = 43'b1100011100000010000000000000000000000001010;
			// PEs: 51 -> 40
			// srcs: (9, 10)(451) -4 --> (451) -4:PEGB3, pass, PUGB5
			8'd3 : rdata = 43'b1100011100000110000000000000000000000001101;
			// PEs: 54 -> 56
			// srcs: (10, 13)(666) 0 --> (666) 0:PEGB6, pass, PUNB
			8'd4 : rdata = 43'b1100011100001100000000000000000001000000000;
			// PEs: 52 -> 56
			// srcs: (11, 15)(740) 1 --> (740) 1:PEGB4, pass, PUNB
			8'd5 : rdata = 43'b1100011100001000000000000000000001000000000;
			// PEs: 54 -> 32
			// srcs: (12, 16)(742) 9 --> (742) 9:PEGB6, pass, PUGB4
			8'd6 : rdata = 43'b1100011100001100000000000000000000000001100;
			// PEs: 32 -> 48
			// srcs: (13, 3)(411) 6 --> (411) 6:PUGB4, pass, NI0
			8'd7 : rdata = 43'b1100011100001001000000000001000000000000000;
			// PEs: 0 -> 49
			// srcs: (19, 2)(608) -4 --> (608) -4:PUGB0, pass, PENB
			8'd8 : rdata = 43'b1100011100000001000000000000000000100000000;
			// PEs: 0 -> 55
			// srcs: (22, 20)(607) -2 --> (607) -2:PUGB0, pass, PEGB7
			8'd9 : rdata = 43'b1100011100000001000000000000000000011110000;
			// PEs: 48 -> 49
			// srcs: (26, 4)(411) 6 --> (411) 6:NI0, pass, PENB
			8'd10 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 16 -> 48
			// srcs: (27, 5)(622) 1 --> (622) 1:PUGB2, pass, NI0
			8'd11 : rdata = 43'b1100011100000101000000000001000000000000000;
			// PEs: 40 -> 49
			// srcs: (28, 6)(426) -3 --> (426) -3:PUNB, pass, PENB
			8'd12 : rdata = 43'b1100011011111111000000000000000000100000000;
			// PEs: 48 -> 49
			// srcs: (34, 7)(622) 1 --> (622) 1:NI0, pass, PENB
			8'd13 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 32 -> 49
			// srcs: (35, 9)(643) 4 --> (643) 4:PUGB4, pass, PENB
			8'd14 : rdata = 43'b1100011100001001000000000000000000100000000;
			// PEs: 40 -> 49
			// srcs: (36, 11)(648) -5 --> (648) -5:PUNB, pass, PENB
			8'd15 : rdata = 43'b1100011011111111000000000000000000100000000;
			// PEs: 40 -> 49
			// srcs: (37, 12)(657) -4 --> (657) -4:PUNB, pass, PENB
			8'd16 : rdata = 43'b1100011011111111000000000000000000100000000;
			// PEs: 8 -> 49
			// srcs: (38, 14)(542) 0 --> (542) 0:PUGB1, pass, PENB
			8'd17 : rdata = 43'b1100011100000011000000000000000000100000000;
			// PEs: 56 -> 48
			// srcs: (39, 17)(745) -2 --> (745) -2:PUGB7, pass, NI0
			8'd18 : rdata = 43'b1100011100001111000000000001000000000000000;
			// PEs: 49 -> 56
			// srcs: (41, 21)(623) -2 --> (623) -2:PEGB1, pass, PUNB
			8'd19 : rdata = 43'b1100011100000010000000000000000001000000000;
			// PEs: 49 -> 0
			// srcs: (42, 25)(644) 10 --> (644) 10:PEGB1, pass, PUGB0
			8'd20 : rdata = 43'b1100011100000010000000000000000000000001000;
			// PEs: 16 -> 49
			// srcs: (43, 18)(551) 9 --> (551) 9:PUGB2, pass, PENB
			8'd21 : rdata = 43'b1100011100000101000000000000000000100000000;
			// PEs: 49 -> 16
			// srcs: (45, 28)(737) 1 --> (737) 1:PEGB1, pass, PUGB2
			8'd22 : rdata = 43'b1100011100000010000000000000000000000001010;
			// PEs: 55 -> 40
			// srcs: (46, 30)(610) 0 --> (610) 0:PENB, pass, PUGB5
			8'd23 : rdata = 43'b1100011011111110000000000000000000000001101;
			// PEs: 48 -> 49
			// srcs: (49, 19)(745) -2 --> (745) -2:NI0, pass, PENB
			8'd24 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 24 -> 48
			// srcs: (50, 22)(631) -3 --> (631) -3:PUGB3, pass, NI0
			8'd25 : rdata = 43'b1100011100000111000000000001000000000000000;
			// PEs: 0 -> 49
			// srcs: (51, 23)(633) 1 --> (633) 1:PUGB0, pass, PENB
			8'd26 : rdata = 43'b1100011100000001000000000000000000100000000;
			// PEs: 48 -> 49
			// srcs: (57, 24)(631) -3 --> (631) -3:NI0, pass, PENB
			8'd27 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 40 -> 49
			// srcs: (58, 26)(647) -9 --> (647) -9:PUNB, pass, PENB
			8'd28 : rdata = 43'b1100011011111111000000000000000000100000000;
			// PEs: 40 -> 49
			// srcs: (59, 27)(656) 11 --> (656) 11:PUNB, pass, PENB
			8'd29 : rdata = 43'b1100011011111111000000000000000000100000000;
			// PEs: 40 -> 53
			// srcs: (60, 29)(748) 7 --> (748) 7:PUNB, pass, PEGB5
			8'd30 : rdata = 43'b1100011011111111000000000000000000011010000;
			// PEs: 49 -> 8
			// srcs: (64, 31)(634) -2 --> (634) -2:PEGB1, pass, PUGB1
			8'd31 : rdata = 43'b1100011100000010000000000000000000000001001;
			// PEs: 0 -> 49
			// srcs: (67, 32)(645) 22 --> (645) 22:PUGB0, pass, PENB
			8'd32 : rdata = 43'b1100011100000001000000000000000000100000000;
			// PEs: 40 -> 48
			// srcs: (68, 33)(733) 5 --> (733) 5:PUNB, pass, NI0
			8'd33 : rdata = 43'b1100011011111111000000000001000000000000000;
			// PEs: 53 -> 56
			// srcs: (72, 36)(749) 14 --> (749) 14:PEGB5, pass, PUNB
			8'd34 : rdata = 43'b1100011100001010000000000000000001000000000;
			// PEs: 50 -> 56
			// srcs: (73, 38)(665) 6 --> (665) 6:PEGB2, pass, PUNB
			8'd35 : rdata = 43'b1100011100000100000000000000000001000000000;
			// PEs: 16 -> 49
			// srcs: (75, 34)(738) 3 --> (738) 3:PUGB2, pass, PENB
			8'd36 : rdata = 43'b1100011100000101000000000000000000100000000;
			// PEs: 49 -> 16
			// srcs: (78, 37)(651) 10 --> (651) 10:PEGB1, pass, PUGB2
			8'd37 : rdata = 43'b1100011100000010000000000000000000000001010;
			// PEs: 48 -> 49
			// srcs: (82, 35)(733) 5 --> (733) 5:NI0, pass, PENB
			8'd38 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 49 -> 56
			// srcs: (89, 39)(739) 8 --> (739) 8:PEGB1, pass, PUNB
			8'd39 : rdata = 43'b1100011100000010000000000000000001000000000;
			// PEs: 0 -> 48
			// srcs: (119, 40)(776) 21 --> (776) 21:PUGB0, pass, NI0
			8'd40 : rdata = 43'b1100011100000001000000000001000000000000000;
			// PEs: 32 -> 49
			// srcs: (122, 41)(800) -20 --> (800) -20:PUGB4, pass, PENB
			8'd41 : rdata = 43'b1100011100001001000000000000000000100000000;
			// PEs: 48 -> 49
			// srcs: (129, 42)(776) 21 --> (776) 21:NI0, pass, PENB
			8'd42 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 40 -> 49
			// srcs: (136, 43)(752) 56 --> (752) 56:PUNB, pass, PENB
			8'd43 : rdata = 43'b1100011011111111000000000000000000100000000;
			// PEs: 49 -> 0
			// srcs: (146, 44)(802) 57 --> (802) 57:PEGB1, pass, PUGB0
			8'd44 : rdata = 43'b1100011100000010000000000000000000000001000;
			// PEs: 32 -> 49
			// srcs: (238, 45)(809) 0 --> (809) 0:PUGB4, pass, PENB
			8'd45 : rdata = 43'b1100011100001001000000000000000000100000000;
			// PEs: 32 -> 50
			// srcs: (241, 46)(809) 0 --> (809) 0:PUGB4, pass, PEGB2
			8'd46 : rdata = 43'b1100011100001001000000000000000000010100000;
			// PEs: 32 -> 51
			// srcs: (244, 47)(809) 0 --> (809) 0:PUGB4, pass, PEGB3
			8'd47 : rdata = 43'b1100011100001001000000000000000000010110000;
			// PEs: 32 -> 52
			// srcs: (247, 48)(809) 0 --> (809) 0:PUGB4, pass, PEGB4
			8'd48 : rdata = 43'b1100011100001001000000000000000000011000000;
			// PEs: 32 -> 53
			// srcs: (254, 49)(809) 0 --> (809) 0:PUGB4, pass, PEGB5
			8'd49 : rdata = 43'b1100011100001001000000000000000000011010000;
			// PEs: 32 -> 49
			// srcs: (255, 50)(809) 0 --> (809) 0:PUGB4, pass, PENB
			8'd50 : rdata = 43'b1100011100001001000000000000000000100000000;
			// PEs: 32 -> 50
			// srcs: (256, 51)(809) 0 --> (809) 0:PUGB4, pass, PEGB2
			8'd51 : rdata = 43'b1100011100001001000000000000000000010100000;
			// PEs: 32 -> 54
			// srcs: (257, 52)(809) 0 --> (809) 0:PUGB4, pass, PEGB6
			8'd52 : rdata = 43'b1100011100001001000000000000000000011100000;
			// PEs: 32 -> 51
			// srcs: (258, 53)(809) 0 --> (809) 0:PUGB4, pass, PEGB3
			8'd53 : rdata = 43'b1100011100001001000000000000000000010110000;
			// PEs: 32 -> 52
			// srcs: (259, 54)(809) 0 --> (809) 0:PUGB4, pass, PEGB4
			8'd54 : rdata = 43'b1100011100001001000000000000000000011000000;
			// PEs: 32 -> 55
			// srcs: (260, 55)(809) 0 --> (809) 0:PUGB4, pass, PEGB7
			8'd55 : rdata = 43'b1100011100001001000000000000000000011110000;
			// PEs: 32 -> 53
			// srcs: (261, 56)(809) 0 --> (809) 0:PUGB4, pass, PEGB5
			8'd56 : rdata = 43'b1100011100001001000000000000000000011010000;
			// PEs: 32 -> 54
			// srcs: (262, 57)(809) 0 --> (809) 0:PUGB4, pass, PEGB6
			8'd57 : rdata = 43'b1100011100001001000000000000000000011100000;
			// PEs: 32 -> 55
			// srcs: (264, 58)(809) 0 --> (809) 0:PUGB4, pass, PEGB7
			8'd58 : rdata = 43'b1100011100001001000000000000000000011110000;
			// PEs: 32 -> 49
			// srcs: (333, 59)(809) 0 --> (809) 0:PUGB4, pass, PENB
			8'd59 : rdata = 43'b1100011100001001000000000000000000100000000;
			// PEs: 32 -> 50
			// srcs: (334, 60)(809) 0 --> (809) 0:PUGB4, pass, PEGB2
			8'd60 : rdata = 43'b1100011100001001000000000000000000010100000;
			// PEs: 32 -> 51
			// srcs: (336, 61)(809) 0 --> (809) 0:PUGB4, pass, PEGB3
			8'd61 : rdata = 43'b1100011100001001000000000000000000010110000;
			// PEs: 32 -> 52
			// srcs: (337, 62)(809) 0 --> (809) 0:PUGB4, pass, PEGB4
			8'd62 : rdata = 43'b1100011100001001000000000000000000011000000;
			// PEs: 32 -> 53
			// srcs: (339, 63)(809) 0 --> (809) 0:PUGB4, pass, PEGB5
			8'd63 : rdata = 43'b1100011100001001000000000000000000011010000;
			// PEs: 32 -> 54
			// srcs: (340, 64)(809) 0 --> (809) 0:PUGB4, pass, PEGB6
			8'd64 : rdata = 43'b1100011100001001000000000000000000011100000;
			// PEs: 32 -> 55
			// srcs: (342, 65)(809) 0 --> (809) 0:PUGB4, pass, PEGB7
			8'd65 : rdata = 43'b1100011100001001000000000000000000011110000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 49) begin
	always @(*) begin
		case(address)
			// PEs: 49, 49 -> 50
			// srcs: (1, 0)(61) 1, (262) -2 --> (462) -2:ND0, NW0, *, PENB
			8'd0 : rdata = 43'b0001101100000000010000000000000000100000000;
			// PEs: 49, 49 -> 50
			// srcs: (2, 1)(139) 0, (340) 0 --> (540) 0:ND1, NW1, *, PENB
			8'd1 : rdata = 43'b0001101100000001010000000010000000100000000;
			// PEs: 49, 49 -> 48
			// srcs: (3, 2)(44) -2, (245) -2 --> (445) 4:ND2, NW2, *, PEGB0
			8'd2 : rdata = 43'b0001101100000010010000000100000000010000000;
			// PEs: 48 -> 
			// srcs: (21, 3)(608) -4 --> (608) -4:PENB, pass, 
			8'd3 : rdata = 43'b1100011011111110000000000000000000000000000;
			// PEs: 49, 48 -> 55
			// srcs: (28, 4)(608) -4, (411) 6 --> (609) 2:ALU, PENB, +, PEGB7
			8'd4 : rdata = 43'b0000100111111111110111111100000000011110000;
			// PEs: 48 -> 
			// srcs: (30, 5)(426) -3 --> (426) -3:PENB, pass, 
			8'd5 : rdata = 43'b1100011011111110000000000000000000000000000;
			// PEs: 48, 49 -> 48
			// srcs: (36, 6)(622) 1, (426) -3 --> (623) -2:PENB, ALU, +, PEGB0
			8'd6 : rdata = 43'b0000111011111110001111111110000000010000000;
			// PEs: 48, 50 -> 48
			// srcs: (37, 7)(643) 4, (448) 6 --> (644) 10:PENB, PEGB2, +, PEGB0
			8'd7 : rdata = 43'b0000111011111110111000001000000000010000000;
			// PEs: 48, 52 -> 49
			// srcs: (38, 8)(648) -5, (454) 2 --> (649) -3:PENB, PEGB4, +, NI0
			8'd8 : rdata = 43'b0000111011111110111000010001000000000000000;
			// PEs: 48, 53 -> 49
			// srcs: (39, 9)(657) -4, (461) 0 --> (658) -4:PENB, PEGB5, +, NI1
			8'd9 : rdata = 43'b0000111011111110111000010101010000000000000;
			// PEs: 50, 48 -> 48
			// srcs: (40, 10)(736) 1, (542) 0 --> (737) 1:PEGB2, PENB, +, PEGB0
			8'd10 : rdata = 43'b0000111100000100110111111100000000010000000;
			// PEs: 48 -> 
			// srcs: (45, 11)(551) 9 --> (551) 9:PENB, pass, 
			8'd11 : rdata = 43'b1100011011111110000000000000000000000000000;
			// PEs: 48, 49 -> 53
			// srcs: (51, 12)(745) -2, (551) 9 --> (746) 7:PENB, ALU, +, PEGB5
			8'd12 : rdata = 43'b0000111011111110001111111110000000011010000;
			// PEs: 48 -> 
			// srcs: (53, 13)(633) 1 --> (633) 1:PENB, pass, 
			8'd13 : rdata = 43'b1100011011111110000000000000000000000000000;
			// PEs: 48, 49 -> 48
			// srcs: (59, 14)(631) -3, (633) 1 --> (634) -2:PENB, ALU, +, PEGB0
			8'd14 : rdata = 43'b0000111011111110001111111110000000010000000;
			// PEs: 48, 49 -> 49
			// srcs: (60, 15)(647) -9, (649) -3 --> (650) -12:PENB, NI0, +, NI2
			8'd15 : rdata = 43'b0000111011111110101000000001100000000000000;
			// PEs: 48, 49 -> 50
			// srcs: (61, 16)(656) 11, (658) -4 --> (659) 7:PENB, NI1, +, PENB
			8'd16 : rdata = 43'b0000111011111110101000000010000000100000000;
			// PEs: 48, 49 -> 48
			// srcs: (73, 17)(645) 22, (650) -12 --> (651) 10:PENB, NI2, +, PEGB0
			8'd17 : rdata = 43'b0000111011111110101000000100000000010000000;
			// PEs: 48 -> 
			// srcs: (77, 18)(738) 3 --> (738) 3:PENB, pass, 
			8'd18 : rdata = 43'b1100011011111110000000000000000000000000000;
			// PEs: 48, 49 -> 48
			// srcs: (84, 19)(733) 5, (738) 3 --> (739) 8:PENB, ALU, +, PEGB0
			8'd19 : rdata = 43'b0000111011111110001111111110000000010000000;
			// PEs: 48 -> 
			// srcs: (124, 20)(800) -20 --> (800) -20:PENB, pass, 
			8'd20 : rdata = 43'b1100011011111110000000000000000000000000000;
			// PEs: 48, 49 -> 
			// srcs: (131, 21)(776) 21, (800) -20 --> (801) 1:PENB, ALU, +, 
			8'd21 : rdata = 43'b0000111011111110001111111110000000000000000;
			// PEs: 48, 49 -> 48
			// srcs: (141, 22)(752) 56, (801) 1 --> (802) 57:PENB, ALU, +, PEGB0
			8'd22 : rdata = 43'b0000111011111110001111111110000000010000000;
			// PEs: 48, 49 -> 50
			// srcs: (240, 23)(809) 0, (44) -2 --> (850) 0:PENB, ND2, *, PENB
			8'd23 : rdata = 43'b0001111011111110011000000100000000100000000;
			// PEs: 49, 50 -> 49
			// srcs: (249, 26)(245) -2, (1050) 0 --> (1250) -2:NW2, PEGB2, -, NW2
			8'd24 : rdata = 43'b0001001000000010111000001000001100000000000;
			// PEs: 48, 49 -> 50
			// srcs: (257, 24)(809) 0, (61) 1 --> (867) 0:PENB, ND0, *, PENB
			8'd25 : rdata = 43'b0001111011111110011000000000000000100000000;
			// PEs: 49, 50 -> 49
			// srcs: (266, 27)(262) -2, (1067) 0 --> (1267) -2:NW0, PEGB2, -, NW0
			8'd26 : rdata = 43'b0001001000000000111000001000001000000000000;
			// PEs: 48, 49 -> 50
			// srcs: (335, 25)(809) 0, (139) 0 --> (945) 0:PENB, ND1, *, PENB
			8'd27 : rdata = 43'b0001111011111110011000000010000000100000000;
			// PEs: 49, 50 -> 49
			// srcs: (344, 28)(340) 0, (1145) 0 --> (1345) 0:NW1, PEGB2, -, NW1
			8'd28 : rdata = 43'b0001001000000001111000001000001010000000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 50) begin
	always @(*) begin
		case(address)
			// PEs: 50, 50 -> 50
			// srcs: (1, 0)(62) -3, (263) 2 --> (463) -6:ND0, NW0, *, NI0
			8'd0 : rdata = 43'b0001101100000000010000000001000000000000000;
			// PEs: 50, 50 -> 50
			// srcs: (2, 1)(140) 1, (341) 1 --> (541) 1:ND1, NW1, *, NI1
			8'd1 : rdata = 43'b0001101100000001010000000011010000000000000;
			// PEs: 50, 50 -> 49
			// srcs: (3, 2)(47) -2, (248) -3 --> (448) 6:ND2, NW2, *, PEGB1
			8'd2 : rdata = 43'b0001101100000010010000000100000000010010000;
			// PEs: 49, 50 -> 51
			// srcs: (4, 3)(462) -2, (463) -6 --> (660) -8:PENB, NI0, +, PENB
			8'd3 : rdata = 43'b0000111011111110101000000000000000100000000;
			// PEs: 49, 50 -> 49
			// srcs: (5, 4)(540) 0, (541) 1 --> (736) 1:PENB, NI1, +, PEGB1
			8'd4 : rdata = 43'b0000111011111110101000000010000000010010000;
			// PEs: 49, 51 -> 48
			// srcs: (67, 5)(659) 7, (664) -1 --> (665) 6:PENB, PEGB3, +, PEGB0
			8'd5 : rdata = 43'b0000111011111110111000001100000000010000000;
			// PEs: 50, 49 -> 49
			// srcs: (243, 9)(3) 1, (850) 0 --> (1050) 0:NM0, PENB, *, PEGB1
			8'd6 : rdata = 43'b0001110000000000110111111100000000010010000;
			// PEs: 48, 50 -> 
			// srcs: (246, 6)(809) 0, (47) -2 --> (853) 0:PEGB0, ND2, *, 
			8'd7 : rdata = 43'b0001111100000000011000000100000000000000000;
			// PEs: 50, 50 -> 
			// srcs: (249, 10)(3) 1, (853) 0 --> (1053) 0:NM0, ALU, *, 
			8'd8 : rdata = 43'b0001110000000000001111111110000000000000000;
			// PEs: 50, 50 -> 50
			// srcs: (252, 13)(248) -3, (1053) 0 --> (1253) -3:NW2, ALU, -, NW2
			8'd9 : rdata = 43'b0001001000000010001111111110001100000000000;
			// PEs: 50, 49 -> 49
			// srcs: (260, 11)(3) 1, (867) 0 --> (1067) 0:NM0, PENB, *, PEGB1
			8'd10 : rdata = 43'b0001110000000000110111111100000000010010000;
			// PEs: 48, 50 -> 51
			// srcs: (261, 7)(809) 0, (62) -3 --> (868) 0:PEGB0, ND0, *, PENB
			8'd11 : rdata = 43'b0001111100000000011000000000000000100000000;
			// PEs: 50, 51 -> 50
			// srcs: (270, 14)(263) 2, (1068) 0 --> (1268) 2:NW0, PEGB3, -, NW0
			8'd12 : rdata = 43'b0001001000000000111000001100001000000000000;
			// PEs: 50, 49 -> 49
			// srcs: (338, 12)(3) 1, (945) 0 --> (1145) 0:NM0, PENB, *, PEGB1
			8'd13 : rdata = 43'b0001110000000000110111111100000000010010000;
			// PEs: 48, 50 -> 51
			// srcs: (339, 8)(809) 0, (140) 1 --> (946) 0:PEGB0, ND1, *, PENB
			8'd14 : rdata = 43'b0001111100000000011000000010000000100000000;
			// PEs: 50, 51 -> 50
			// srcs: (348, 15)(341) 1, (1146) 0 --> (1346) 1:NW1, PEGB3, -, NW1
			8'd15 : rdata = 43'b0001001000000001111000001100001010000000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 51) begin
	always @(*) begin
		case(address)
			// PEs: 51, 51 -> 52
			// srcs: (1, 0)(64) -1, (265) -1 --> (465) 1:ND0, NW0, *, PENB
			8'd0 : rdata = 43'b0001101100000000010000000000000000100000000;
			// PEs: 51, 51 -> 52
			// srcs: (2, 1)(142) -1, (343) -1 --> (543) 1:ND1, NW1, *, PENB
			8'd1 : rdata = 43'b0001101100000001010000000010000000100000000;
			// PEs: 51, 51 -> 48
			// srcs: (3, 2)(50) -2, (251) 2 --> (451) -4:ND2, NW2, *, PEGB0
			8'd2 : rdata = 43'b0001101100000010010000000100000000010000000;
			// PEs: 50, 54 -> 
			// srcs: (10, 3)(660) -8, (464) 6 --> (661) -2:PENB, PEGB6, +, 
			8'd3 : rdata = 43'b0000111011111110111000011000000000000000000;
			// PEs: 51, 53 -> 50
			// srcs: (16, 4)(661) -2, (663) 1 --> (664) -1:ALU, PEGB5, +, PEGB2
			8'd4 : rdata = 43'b0000100111111111111000010100000000010100000;
			// PEs: 48, 51 -> 
			// srcs: (249, 5)(809) 0, (50) -2 --> (856) 0:PEGB0, ND2, *, 
			8'd5 : rdata = 43'b0001111100000000011000000100000000000000000;
			// PEs: 51, 51 -> 
			// srcs: (252, 8)(3) 1, (856) 0 --> (1056) 0:NM0, ALU, *, 
			8'd6 : rdata = 43'b0001110000000000001111111110000000000000000;
			// PEs: 51, 51 -> 51
			// srcs: (255, 12)(251) 2, (1056) 0 --> (1256) 2:NW2, ALU, -, NW2
			8'd7 : rdata = 43'b0001001000000010001111111110001100000000000;
			// PEs: 48, 51 -> 52
			// srcs: (263, 6)(809) 0, (64) -1 --> (870) 0:PEGB0, ND0, *, PENB
			8'd8 : rdata = 43'b0001111100000000011000000000000000100000000;
			// PEs: 51, 50 -> 50
			// srcs: (264, 9)(3) 1, (868) 0 --> (1068) 0:NM0, PENB, *, PEGB2
			8'd9 : rdata = 43'b0001110000000000110111111100000000010100000;
			// PEs: 51, 52 -> 51
			// srcs: (272, 13)(265) -1, (1070) 0 --> (1270) -1:NW0, PEGB4, -, NW0
			8'd10 : rdata = 43'b0001001000000000111000010000001000000000000;
			// PEs: 48, 51 -> 51
			// srcs: (341, 7)(809) 0, (142) -1 --> (948) 0:PEGB0, ND1, *, NI0
			8'd11 : rdata = 43'b0001111100000000011000000011000000000000000;
			// PEs: 51, 50 -> 50
			// srcs: (342, 10)(3) 1, (946) 0 --> (1146) 0:NM0, PENB, *, PEGB2
			8'd12 : rdata = 43'b0001110000000000110111111100000000010100000;
			// PEs: 51, 51 -> 
			// srcs: (344, 11)(3) 1, (948) 0 --> (1148) 0:NM0, NI0, *, 
			8'd13 : rdata = 43'b0001110000000000101000000000000000000000000;
			// PEs: 51, 51 -> 51
			// srcs: (347, 14)(343) -1, (1148) 0 --> (1348) -1:NW1, ALU, -, NW1
			8'd14 : rdata = 43'b0001001000000001001111111110001010000000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 52) begin
	always @(*) begin
		case(address)
			// PEs: 52, 52 -> 52
			// srcs: (1, 0)(65) 2, (266) 0 --> (466) 0:ND0, NW0, *, NI0
			8'd0 : rdata = 43'b0001101100000000010000000001000000000000000;
			// PEs: 52, 52 -> 52
			// srcs: (2, 1)(143) 0, (344) 2 --> (544) 0:ND1, NW1, *, NI1
			8'd1 : rdata = 43'b0001101100000001010000000011010000000000000;
			// PEs: 52, 52 -> 49
			// srcs: (3, 2)(53) -2, (254) -1 --> (454) 2:ND2, NW2, *, PEGB1
			8'd2 : rdata = 43'b0001101100000010010000000100000000010010000;
			// PEs: 51, 52 -> 53
			// srcs: (4, 3)(465) 1, (466) 0 --> (662) 1:PENB, NI0, +, PENB
			8'd3 : rdata = 43'b0000111011111110101000000000000000100000000;
			// PEs: 51, 52 -> 48
			// srcs: (5, 4)(543) 1, (544) 0 --> (740) 1:PENB, NI1, +, PEGB0
			8'd4 : rdata = 43'b0000111011111110101000000010000000010000000;
			// PEs: 48, 52 -> 
			// srcs: (252, 5)(809) 0, (53) -2 --> (859) 0:PEGB0, ND2, *, 
			8'd5 : rdata = 43'b0001111100000000011000000100000000000000000;
			// PEs: 52, 52 -> 
			// srcs: (255, 8)(3) 1, (859) 0 --> (1059) 0:NM0, ALU, *, 
			8'd6 : rdata = 43'b0001110000000000001111111110000000000000000;
			// PEs: 52, 52 -> 52
			// srcs: (258, 11)(254) -1, (1059) 0 --> (1259) -1:NW2, ALU, -, NW2
			8'd7 : rdata = 43'b0001001000000010001111111110001100000000000;
			// PEs: 48, 52 -> 52
			// srcs: (264, 6)(809) 0, (65) 2 --> (871) 0:PEGB0, ND0, *, NI0
			8'd8 : rdata = 43'b0001111100000000011000000001000000000000000;
			// PEs: 52, 51 -> 51
			// srcs: (266, 9)(3) 1, (870) 0 --> (1070) 0:NM0, PENB, *, PEGB3
			8'd9 : rdata = 43'b0001110000000000110111111100000000010110000;
			// PEs: 52, 52 -> 
			// srcs: (267, 10)(3) 1, (871) 0 --> (1071) 0:NM0, NI0, *, 
			8'd10 : rdata = 43'b0001110000000000101000000000000000000000000;
			// PEs: 52, 52 -> 52
			// srcs: (270, 12)(266) 0, (1071) 0 --> (1271) 0:NW0, ALU, -, NW0
			8'd11 : rdata = 43'b0001001000000000001111111110001000000000000;
			// PEs: 48, 52 -> 53
			// srcs: (342, 7)(809) 0, (143) 0 --> (949) 0:PEGB0, ND1, *, PENB
			8'd12 : rdata = 43'b0001111100000000011000000010000000100000000;
			// PEs: 52, 53 -> 52
			// srcs: (351, 13)(344) 2, (1149) 0 --> (1349) 2:NW1, PEGB5, -, NW1
			8'd13 : rdata = 43'b0001001000000001111000010100001010000000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 53) begin
	always @(*) begin
		case(address)
			// PEs: 53, 53 -> 54
			// srcs: (1, 0)(67) -3, (268) 0 --> (468) 0:ND0, NW0, *, PENB
			8'd0 : rdata = 43'b0001101100000000010000000000000000100000000;
			// PEs: 53, 53 -> 54
			// srcs: (2, 1)(145) -3, (346) -3 --> (546) 9:ND1, NW1, *, PENB
			8'd1 : rdata = 43'b0001101100000001010000000010000000100000000;
			// PEs: 53, 53 -> 49
			// srcs: (3, 2)(60) 0, (261) 1 --> (461) 0:ND2, NW2, *, PEGB1
			8'd2 : rdata = 43'b0001101100000010010000000100000000010010000;
			// PEs: 52, 55 -> 51
			// srcs: (10, 3)(662) 1, (467) 0 --> (663) 1:PENB, PEGB7, +, PEGB3
			8'd3 : rdata = 43'b0000111011111110111000011100000000010110000;
			// PEs: 48 -> 
			// srcs: (65, 4)(748) 7 --> (748) 7:PEGB0, pass, 
			8'd4 : rdata = 43'b1100011100000000000000000000000000000000000;
			// PEs: 49, 53 -> 48
			// srcs: (67, 5)(746) 7, (748) 7 --> (749) 14:PEGB1, ALU, +, PEGB0
			8'd5 : rdata = 43'b0000111100000010001111111110000000010000000;
			// PEs: 48, 53 -> 
			// srcs: (259, 6)(809) 0, (60) 0 --> (866) 0:PEGB0, ND2, *, 
			8'd6 : rdata = 43'b0001111100000000011000000100000000000000000;
			// PEs: 53, 53 -> 
			// srcs: (262, 9)(3) 1, (866) 0 --> (1066) 0:NM0, ALU, *, 
			8'd7 : rdata = 43'b0001110000000000001111111110000000000000000;
			// PEs: 53, 53 -> 53
			// srcs: (265, 11)(261) 1, (1066) 0 --> (1266) 1:NW2, ALU, -, NW2
			8'd8 : rdata = 43'b0001001000000010001111111110001100000000000;
			// PEs: 48, 53 -> 54
			// srcs: (266, 7)(809) 0, (67) -3 --> (873) 0:PEGB0, ND0, *, PENB
			8'd9 : rdata = 43'b0001111100000000011000000000000000100000000;
			// PEs: 53, 54 -> 53
			// srcs: (275, 12)(268) 0, (1073) 0 --> (1273) 0:NW0, PEGB6, -, NW0
			8'd10 : rdata = 43'b0001001000000000111000011000001000000000000;
			// PEs: 48, 53 -> 54
			// srcs: (344, 8)(809) 0, (145) -3 --> (951) 0:PEGB0, ND1, *, PENB
			8'd11 : rdata = 43'b0001111100000000011000000010000000100000000;
			// PEs: 53, 52 -> 52
			// srcs: (345, 10)(3) 1, (949) 0 --> (1149) 0:NM0, PENB, *, PEGB4
			8'd12 : rdata = 43'b0001110000000000110111111100000000011000000;
			// PEs: 53, 54 -> 53
			// srcs: (353, 13)(346) -3, (1151) 0 --> (1351) -3:NW1, PEGB6, -, NW1
			8'd13 : rdata = 43'b0001001000000001111000011000001010000000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 54) begin
	always @(*) begin
		case(address)
			// PEs: 54, 54 -> 54
			// srcs: (1, 0)(68) 0, (269) -2 --> (469) 0:ND0, NW0, *, NI0
			8'd0 : rdata = 43'b0001101100000000010000000001000000000000000;
			// PEs: 54, 54 -> 54
			// srcs: (2, 1)(146) 0, (347) 2 --> (547) 0:ND1, NW1, *, NI1
			8'd1 : rdata = 43'b0001101100000001010000000011010000000000000;
			// PEs: 54, 54 -> 51
			// srcs: (3, 2)(63) -2, (264) -3 --> (464) 6:ND2, NW2, *, PEGB3
			8'd2 : rdata = 43'b0001101100000010010000000100000000010110000;
			// PEs: 53, 54 -> 48
			// srcs: (4, 3)(468) 0, (469) 0 --> (666) 0:PENB, NI0, +, PEGB0
			8'd3 : rdata = 43'b0000111011111110101000000000000000010000000;
			// PEs: 53, 54 -> 48
			// srcs: (5, 4)(546) 9, (547) 0 --> (742) 9:PENB, NI1, +, PEGB0
			8'd4 : rdata = 43'b0000111011111110101000000010000000010000000;
			// PEs: 48, 54 -> 
			// srcs: (262, 5)(809) 0, (63) -2 --> (869) 0:PEGB0, ND2, *, 
			8'd5 : rdata = 43'b0001111100000000011000000100000000000000000;
			// PEs: 54, 54 -> 54
			// srcs: (265, 8)(3) 1, (869) 0 --> (1069) 0:NM0, ALU, *, NI0
			8'd6 : rdata = 43'b0001110000000000001111111111000000000000000;
			// PEs: 48, 54 -> 55
			// srcs: (267, 6)(809) 0, (68) 0 --> (874) 0:PEGB0, ND0, *, PENB
			8'd7 : rdata = 43'b0001111100000000011000000000000000100000000;
			// PEs: 54, 54 -> 54
			// srcs: (268, 12)(264) -3, (1069) 0 --> (1269) -3:NW2, NI0, -, NW2
			8'd8 : rdata = 43'b0001001000000010101000000000001100000000000;
			// PEs: 54, 53 -> 53
			// srcs: (269, 9)(3) 1, (873) 0 --> (1073) 0:NM0, PENB, *, PEGB5
			8'd9 : rdata = 43'b0001110000000000110111111100000000011010000;
			// PEs: 54, 55 -> 54
			// srcs: (276, 13)(269) -2, (1074) 0 --> (1274) -2:NW0, PEGB7, -, NW0
			8'd10 : rdata = 43'b0001001000000000111000011100001000000000000;
			// PEs: 48, 54 -> 54
			// srcs: (345, 7)(809) 0, (146) 0 --> (952) 0:PEGB0, ND1, *, NI0
			8'd11 : rdata = 43'b0001111100000000011000000011000000000000000;
			// PEs: 54, 53 -> 53
			// srcs: (347, 10)(3) 1, (951) 0 --> (1151) 0:NM0, PENB, *, PEGB5
			8'd12 : rdata = 43'b0001110000000000110111111100000000011010000;
			// PEs: 54, 54 -> 
			// srcs: (348, 11)(3) 1, (952) 0 --> (1152) 0:NM0, NI0, *, 
			8'd13 : rdata = 43'b0001110000000000101000000000000000000000000;
			// PEs: 54, 54 -> 54
			// srcs: (351, 14)(347) 2, (1152) 0 --> (1352) 2:NW1, ALU, -, NW1
			8'd14 : rdata = 43'b0001001000000001001111111110001010000000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 55) begin
	always @(*) begin
		case(address)
			// PEs: 55, 55 -> 48
			// srcs: (1, 0)(70) -1, (271) -2 --> (471) 2:ND0, NW0, *, PENB
			8'd0 : rdata = 43'b0001101100000000010000000000000000100000000;
			// PEs: 55, 55 -> 48
			// srcs: (2, 1)(148) -3, (349) 2 --> (549) -6:ND1, NW1, *, PENB
			8'd1 : rdata = 43'b0001101100000001010000000010000000100000000;
			// PEs: 55, 55 -> 53
			// srcs: (3, 2)(66) -1, (267) 0 --> (467) 0:ND2, NW2, *, PEGB5
			8'd2 : rdata = 43'b0001101100000010010000000100000000011010000;
			// PEs: 49 -> 
			// srcs: (33, 3)(609) 2 --> (609) 2:PEGB1, pass, 
			8'd3 : rdata = 43'b1100011100000010000000000000000000000000000;
			// PEs: 48, 55 -> 48
			// srcs: (43, 4)(607) -2, (609) 2 --> (610) 0:PEGB0, ALU, +, PENB
			8'd4 : rdata = 43'b0000111100000000001111111110000000100000000;
			// PEs: 48, 55 -> 
			// srcs: (265, 5)(809) 0, (66) -1 --> (872) 0:PEGB0, ND2, *, 
			8'd5 : rdata = 43'b0001111100000000011000000100000000000000000;
			// PEs: 55, 55 -> 55
			// srcs: (268, 8)(3) 1, (872) 0 --> (1072) 0:NM0, ALU, *, NI0
			8'd6 : rdata = 43'b0001110000000000001111111111000000000000000;
			// PEs: 48, 55 -> 55
			// srcs: (269, 6)(809) 0, (70) -1 --> (876) 0:PEGB0, ND0, *, NI1
			8'd7 : rdata = 43'b0001111100000000011000000001010000000000000;
			// PEs: 55, 54 -> 54
			// srcs: (270, 9)(3) 1, (874) 0 --> (1074) 0:NM0, PENB, *, PEGB6
			8'd8 : rdata = 43'b0001110000000000110111111100000000011100000;
			// PEs: 55, 55 -> 55
			// srcs: (271, 12)(267) 0, (1072) 0 --> (1272) 0:NW2, NI0, -, NW2
			8'd9 : rdata = 43'b0001001000000010101000000000001100000000000;
			// PEs: 55, 55 -> 
			// srcs: (272, 10)(3) 1, (876) 0 --> (1076) 0:NM0, NI1, *, 
			8'd10 : rdata = 43'b0001110000000000101000000010000000000000000;
			// PEs: 55, 55 -> 55
			// srcs: (275, 13)(271) -2, (1076) 0 --> (1276) -2:NW0, ALU, -, NW0
			8'd11 : rdata = 43'b0001001000000000001111111110001000000000000;
			// PEs: 48, 55 -> 
			// srcs: (347, 7)(809) 0, (148) -3 --> (954) 0:PEGB0, ND1, *, 
			8'd12 : rdata = 43'b0001111100000000011000000010000000000000000;
			// PEs: 55, 55 -> 
			// srcs: (350, 11)(3) 1, (954) 0 --> (1154) 0:NM0, ALU, *, 
			8'd13 : rdata = 43'b0001110000000000001111111110000000000000000;
			// PEs: 55, 55 -> 55
			// srcs: (353, 14)(349) 2, (1154) 0 --> (1354) 2:NW1, ALU, -, NW1
			8'd14 : rdata = 43'b0001001000000001001111111110001010000000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 56) begin
	always @(*) begin
		case(address)
			// PEs: 48 -> 57
			// srcs: (5, 0)(471) 2 --> (471) 2:PUNB, pass, PENB
			8'd0 : rdata = 43'b1100011011111111000000000000000000100000000;
			// PEs: 48 -> 57
			// srcs: (6, 1)(549) -6 --> (549) -6:PUNB, pass, PENB
			8'd1 : rdata = 43'b1100011011111111000000000000000000100000000;
			// PEs: 63 -> 0
			// srcs: (7, 6)(678) -1 --> (678) -1:PENB, pass, PUNB
			8'd2 : rdata = 43'b1100011011111110000000000000000001000000000;
			// PEs: 61 -> 0
			// srcs: (8, 7)(486) 6 --> (486) 6:PEGB5, pass, PUNB
			8'd3 : rdata = 43'b1100011100001010000000000000000001000000000;
			// PEs: 62 -> 0
			// srcs: (9, 8)(489) -6 --> (489) -6:PEGB6, pass, PUNB
			8'd4 : rdata = 43'b1100011100001100000000000000000001000000000;
			// PEs: 59 -> 40
			// srcs: (10, 17)(747) 7 --> (747) 7:PEGB3, pass, PUGB5
			8'd5 : rdata = 43'b1100011100000110000000000000000000000001101;
			// PEs: 63 -> 8
			// srcs: (14, 9)(492) 2 --> (492) 2:PENB, pass, PUGB1
			8'd6 : rdata = 43'b1100011011111110000000000000000000000001001;
			// PEs: 57 -> 48
			// srcs: (15, 16)(745) -2 --> (745) -2:PEGB1, pass, PUGB6
			8'd7 : rdata = 43'b1100011100000010000000000000000000000001110;
			// PEs: 62 -> 0
			// srcs: (16, 24)(755) 16 --> (755) 16:PEGB6, pass, PUNB
			8'd8 : rdata = 43'b1100011100001100000000000000000001000000000;
			// PEs: 16 -> 56
			// srcs: (20, 2)(624) 2 --> (624) 2:PUGB2, pass, NI0
			8'd9 : rdata = 43'b1100011100000101000000000001000000000000000;
			// PEs: 40 -> 57
			// srcs: (21, 3)(429) 1 --> (429) 1:PUGB5, pass, PENB
			8'd10 : rdata = 43'b1100011100001011000000000000000000100000000;
			// PEs: 56 -> 57
			// srcs: (27, 4)(624) 2 --> (624) 2:NI0, pass, PENB
			8'd11 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 48 -> 57
			// srcs: (28, 5)(666) 0 --> (666) 0:PUNB, pass, PENB
			8'd12 : rdata = 43'b1100011011111111000000000000000000100000000;
			// PEs: 24 -> 56
			// srcs: (29, 10)(707) -4 --> (707) -4:PUGB3, pass, NI0
			8'd13 : rdata = 43'b1100011100000111000000000001000000000000000;
			// PEs: 0 -> 57
			// srcs: (30, 11)(511) 4 --> (511) 4:PUGB0, pass, PENB
			8'd14 : rdata = 43'b1100011100000001000000000000000000100000000;
			// PEs: 56 -> 57
			// srcs: (36, 12)(707) -4 --> (707) -4:NI0, pass, PENB
			8'd15 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 48 -> 56
			// srcs: (37, 13)(740) 1 --> (740) 1:PUNB, pass, NI0
			8'd16 : rdata = 43'b1100011011111111000000000001000000000000000;
			// PEs: 16 -> 57
			// srcs: (42, 14)(545) -3 --> (545) -3:PUGB2, pass, PENB
			8'd17 : rdata = 43'b1100011100000101000000000000000000100000000;
			// PEs: 56 -> 57
			// srcs: (48, 15)(740) 1 --> (740) 1:NI0, pass, PENB
			8'd18 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 56
			// srcs: (49, 18)(759) 2 --> (759) 2:PUGB0, pass, NI0
			8'd19 : rdata = 43'b1100011100000001000000000001000000000000000;
			// PEs: 16 -> 57
			// srcs: (50, 19)(564) -4 --> (564) -4:PUGB2, pass, PENB
			8'd20 : rdata = 43'b1100011100000101000000000000000000100000000;
			// PEs: 57 -> 24
			// srcs: (55, 23)(741) -2 --> (741) -2:PEGB1, pass, PUGB3
			8'd21 : rdata = 43'b1100011100000010000000000000000000000001011;
			// PEs: 56 -> 57
			// srcs: (56, 20)(759) 2 --> (759) 2:NI0, pass, PENB
			8'd22 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 48 -> 57
			// srcs: (57, 21)(623) -2 --> (623) -2:PUNB, pass, PENB
			8'd23 : rdata = 43'b1100011011111111000000000000000000100000000;
			// PEs: 57 -> 0
			// srcs: (63, 25)(760) -2 --> (760) -2:PEGB1, pass, PUNB
			8'd24 : rdata = 43'b1100011100000010000000000000000001000000000;
			// PEs: 16 -> 57
			// srcs: (67, 22)(706) 1 --> (706) 1:PUGB2, pass, PENB
			8'd25 : rdata = 43'b1100011100000101000000000000000000100000000;
			// PEs: 40 -> 57
			// srcs: (68, 26)(621) 4 --> (621) 4:PUGB5, pass, PENB
			8'd26 : rdata = 43'b1100011100001011000000000000000000100000000;
			// PEs: 24 -> 57
			// srcs: (69, 27)(714) 8 --> (714) 8:PUGB3, pass, PENB
			8'd27 : rdata = 43'b1100011100000111000000000000000000100000000;
			// PEs: 57 -> 8
			// srcs: (77, 31)(627) 5 --> (627) 5:PEGB1, pass, PUGB1
			8'd28 : rdata = 43'b1100011100000010000000000000000000000001001;
			// PEs: 57 -> 40
			// srcs: (87, 33)(715) 9 --> (715) 9:PEGB1, pass, PUGB5
			8'd29 : rdata = 43'b1100011100000010000000000000000000000001101;
			// PEs: 24 -> 56
			// srcs: (97, 28)(744) 7 --> (744) 7:PUGB3, pass, NI0
			8'd30 : rdata = 43'b1100011100000111000000000001000000000000000;
			// PEs: 48 -> 57
			// srcs: (98, 29)(749) 14 --> (749) 14:PUNB, pass, PENB
			8'd31 : rdata = 43'b1100011011111111000000000000000000100000000;
			// PEs: 56 -> 57
			// srcs: (104, 30)(744) 7 --> (744) 7:NI0, pass, PENB
			8'd32 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 48 -> 57
			// srcs: (105, 32)(665) 6 --> (665) 6:PUNB, pass, PENB
			8'd33 : rdata = 43'b1100011011111111000000000000000000100000000;
			// PEs: 48 -> 57
			// srcs: (106, 34)(739) 8 --> (739) 8:PUNB, pass, PENB
			8'd34 : rdata = 43'b1100011011111111000000000000000000100000000;
			// PEs: 57 -> 24
			// srcs: (112, 35)(677) 16 --> (677) 16:PEGB1, pass, PUGB3
			8'd35 : rdata = 43'b1100011100000010000000000000000000000001011;
			// PEs: 57 -> 40
			// srcs: (121, 36)(751) 29 --> (751) 29:PEGB1, pass, PUGB5
			8'd36 : rdata = 43'b1100011100000010000000000000000000000001101;
			// PEs: 32 -> 57
			// srcs: (263, 37)(809) 0 --> (809) 0:PUGB4, pass, PENB
			8'd37 : rdata = 43'b1100011100001001000000000000000000100000000;
			// PEs: 32 -> 57
			// srcs: (265, 38)(809) 0 --> (809) 0:PUGB4, pass, PENB
			8'd38 : rdata = 43'b1100011100001001000000000000000000100000000;
			// PEs: 32 -> 58
			// srcs: (266, 39)(809) 0 --> (809) 0:PUGB4, pass, PEGB2
			8'd39 : rdata = 43'b1100011100001001000000000000000000010100000;
			// PEs: 32 -> 58
			// srcs: (267, 40)(809) 0 --> (809) 0:PUGB4, pass, PEGB2
			8'd40 : rdata = 43'b1100011100001001000000000000000000010100000;
			// PEs: 32 -> 59
			// srcs: (268, 41)(809) 0 --> (809) 0:PUGB4, pass, PEGB3
			8'd41 : rdata = 43'b1100011100001001000000000000000000010110000;
			// PEs: 32 -> 59
			// srcs: (269, 42)(809) 0 --> (809) 0:PUGB4, pass, PEGB3
			8'd42 : rdata = 43'b1100011100001001000000000000000000010110000;
			// PEs: 32 -> 60
			// srcs: (270, 43)(809) 0 --> (809) 0:PUGB4, pass, PEGB4
			8'd43 : rdata = 43'b1100011100001001000000000000000000011000000;
			// PEs: 32 -> 61
			// srcs: (271, 44)(809) 0 --> (809) 0:PUGB4, pass, PEGB5
			8'd44 : rdata = 43'b1100011100001001000000000000000000011010000;
			// PEs: 32 -> 60
			// srcs: (272, 45)(809) 0 --> (809) 0:PUGB4, pass, PEGB4
			8'd45 : rdata = 43'b1100011100001001000000000000000000011000000;
			// PEs: 32 -> 62
			// srcs: (273, 46)(809) 0 --> (809) 0:PUGB4, pass, PEGB6
			8'd46 : rdata = 43'b1100011100001001000000000000000000011100000;
			// PEs: 32 -> 63
			// srcs: (274, 47)(809) 0 --> (809) 0:PUGB4, pass, PEGB7
			8'd47 : rdata = 43'b1100011100001001000000000000000000011110000;
			// PEs: 32 -> 61
			// srcs: (279, 48)(809) 0 --> (809) 0:PUGB4, pass, PEGB5
			8'd48 : rdata = 43'b1100011100001001000000000000000000011010000;
			// PEs: 32 -> 62
			// srcs: (282, 49)(809) 0 --> (809) 0:PUGB4, pass, PEGB6
			8'd49 : rdata = 43'b1100011100001001000000000000000000011100000;
			// PEs: 32 -> 63
			// srcs: (285, 50)(809) 0 --> (809) 0:PUGB4, pass, PEGB7
			8'd50 : rdata = 43'b1100011100001001000000000000000000011110000;
			// PEs: 32 -> 57
			// srcs: (343, 51)(809) 0 --> (809) 0:PUGB4, pass, PENB
			8'd51 : rdata = 43'b1100011100001001000000000000000000100000000;
			// PEs: 32 -> 58
			// srcs: (345, 52)(809) 0 --> (809) 0:PUGB4, pass, PEGB2
			8'd52 : rdata = 43'b1100011100001001000000000000000000010100000;
			// PEs: 32 -> 59
			// srcs: (346, 53)(809) 0 --> (809) 0:PUGB4, pass, PEGB3
			8'd53 : rdata = 43'b1100011100001001000000000000000000010110000;
			// PEs: 32 -> 60
			// srcs: (348, 54)(809) 0 --> (809) 0:PUGB4, pass, PEGB4
			8'd54 : rdata = 43'b1100011100001001000000000000000000011000000;
			// PEs: 32 -> 61
			// srcs: (349, 55)(809) 0 --> (809) 0:PUGB4, pass, PEGB5
			8'd55 : rdata = 43'b1100011100001001000000000000000000011010000;
			// PEs: 32 -> 62
			// srcs: (350, 56)(809) 0 --> (809) 0:PUGB4, pass, PEGB6
			8'd56 : rdata = 43'b1100011100001001000000000000000000011100000;
			// PEs: 32 -> 63
			// srcs: (351, 57)(809) 0 --> (809) 0:PUGB4, pass, PEGB7
			8'd57 : rdata = 43'b1100011100001001000000000000000000011110000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 57) begin
	always @(*) begin
		case(address)
			// PEs: 57, 57 -> 57
			// srcs: (1, 0)(71) 0, (272) -3 --> (472) 0:ND0, NW0, *, NI0
			8'd0 : rdata = 43'b0001101100000000010000000001000000000000000;
			// PEs: 57, 57 -> 57
			// srcs: (2, 1)(149) -2, (350) -2 --> (550) 4:ND1, NW1, *, NI1
			8'd1 : rdata = 43'b0001101100000001010000000011010000000000000;
			// PEs: 57, 57 -> 57
			// srcs: (3, 2)(69) -1, (270) -3 --> (470) 3:ND2, NW2, *, NI2
			8'd2 : rdata = 43'b0001101100000010010000000101100000000000000;
			// PEs: 56, 57 -> 58
			// srcs: (8, 3)(471) 2, (472) 0 --> (668) 2:PENB, NI0, +, PENB
			8'd3 : rdata = 43'b0000111011111110101000000000000000100000000;
			// PEs: 56, 57 -> 56
			// srcs: (9, 4)(549) -6, (550) 4 --> (745) -2:PENB, NI1, +, PEGB0
			8'd4 : rdata = 43'b0000111011111110101000000010000000010000000;
			// PEs: 56 -> 
			// srcs: (23, 5)(429) 1 --> (429) 1:PENB, pass, 
			8'd5 : rdata = 43'b1100011011111110000000000000000000000000000;
			// PEs: 56, 57 -> 57
			// srcs: (29, 6)(624) 2, (429) 1 --> (625) 3:PENB, ALU, +, NI0
			8'd6 : rdata = 43'b0000111011111110001111111111000000000000000;
			// PEs: 56, 57 -> 58
			// srcs: (30, 7)(666) 0, (470) 3 --> (667) 3:PENB, NI2, +, PENB
			8'd7 : rdata = 43'b0000111011111110101000000100000000100000000;
			// PEs: 56 -> 
			// srcs: (32, 8)(511) 4 --> (511) 4:PENB, pass, 
			8'd8 : rdata = 43'b1100011011111110000000000000000000000000000;
			// PEs: 56, 57 -> 57
			// srcs: (38, 9)(707) -4, (511) 4 --> (708) 0:PENB, ALU, +, NI1
			8'd9 : rdata = 43'b0000111011111110001111111111010000000000000;
			// PEs: 56 -> 
			// srcs: (44, 10)(545) -3 --> (545) -3:PENB, pass, 
			8'd10 : rdata = 43'b1100011011111110000000000000000000000000000;
			// PEs: 56, 57 -> 56
			// srcs: (50, 11)(740) 1, (545) -3 --> (741) -2:PENB, ALU, +, PEGB0
			8'd11 : rdata = 43'b0000111011111110001111111110000000010000000;
			// PEs: 56 -> 
			// srcs: (52, 12)(564) -4 --> (564) -4:PENB, pass, 
			8'd12 : rdata = 43'b1100011011111110000000000000000000000000000;
			// PEs: 56, 57 -> 56
			// srcs: (58, 13)(759) 2, (564) -4 --> (760) -2:PENB, ALU, +, PEGB0
			8'd13 : rdata = 43'b0000111011111110001111111110000000010000000;
			// PEs: 56, 57 -> 57
			// srcs: (59, 14)(623) -2, (625) 3 --> (626) 1:PENB, NI0, +, NI2
			8'd14 : rdata = 43'b0000111011111110101000000001100000000000000;
			// PEs: 56, 57 -> 57
			// srcs: (69, 15)(706) 1, (708) 0 --> (709) 1:PENB, NI1, +, NI0
			8'd15 : rdata = 43'b0000111011111110101000000011000000000000000;
			// PEs: 56, 57 -> 56
			// srcs: (72, 16)(621) 4, (626) 1 --> (627) 5:PENB, NI2, +, PEGB0
			8'd16 : rdata = 43'b0000111011111110101000000100000000010000000;
			// PEs: 57, 56 -> 56
			// srcs: (82, 17)(709) 1, (714) 8 --> (715) 9:NI0, PENB, +, PEGB0
			8'd17 : rdata = 43'b0000110100000000110111111100000000010000000;
			// PEs: 56 -> 
			// srcs: (100, 18)(749) 14 --> (749) 14:PENB, pass, 
			8'd18 : rdata = 43'b1100011011111110000000000000000000000000000;
			// PEs: 56, 57 -> 57
			// srcs: (106, 19)(744) 7, (749) 14 --> (750) 21:PENB, ALU, +, NI0
			8'd19 : rdata = 43'b0000111011111110001111111111000000000000000;
			// PEs: 56, 62 -> 56
			// srcs: (107, 20)(665) 6, (676) 10 --> (677) 16:PENB, PEGB6, +, PEGB0
			8'd20 : rdata = 43'b0000111011111110111000011000000000010000000;
			// PEs: 56, 57 -> 56
			// srcs: (116, 21)(739) 8, (750) 21 --> (751) 29:PENB, NI0, +, PEGB0
			8'd21 : rdata = 43'b0000111011111110101000000000000000010000000;
			// PEs: 56, 57 -> 58
			// srcs: (265, 22)(809) 0, (69) -1 --> (875) 0:PENB, ND2, *, PENB
			8'd22 : rdata = 43'b0001111011111110011000000100000000100000000;
			// PEs: 56, 57 -> 58
			// srcs: (267, 23)(809) 0, (71) 0 --> (877) 0:PENB, ND0, *, PENB
			8'd23 : rdata = 43'b0001111011111110011000000000000000100000000;
			// PEs: 57, 58 -> 57
			// srcs: (274, 25)(270) -3, (1075) 0 --> (1275) -3:NW2, PEGB2, -, NW2
			8'd24 : rdata = 43'b0001001000000010111000001000001100000000000;
			// PEs: 57, 58 -> 57
			// srcs: (276, 26)(272) -3, (1077) 0 --> (1277) -3:NW0, PEGB2, -, NW0
			8'd25 : rdata = 43'b0001001000000000111000001000001000000000000;
			// PEs: 56, 57 -> 58
			// srcs: (345, 24)(809) 0, (149) -2 --> (955) 0:PENB, ND1, *, PENB
			8'd26 : rdata = 43'b0001111011111110011000000010000000100000000;
			// PEs: 57, 58 -> 57
			// srcs: (354, 27)(350) -2, (1155) 0 --> (1355) -2:NW1, PEGB2, -, NW1
			8'd27 : rdata = 43'b0001001000000001111000001000001010000000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 58) begin
	always @(*) begin
		case(address)
			// PEs: 58, 58 -> 59
			// srcs: (1, 0)(73) -3, (274) -2 --> (474) 6:ND0, NW0, *, PENB
			8'd0 : rdata = 43'b0001101100000000010000000000000000100000000;
			// PEs: 58, 58 -> 59
			// srcs: (2, 1)(151) 2, (352) -1 --> (552) -2:ND1, NW1, *, PENB
			8'd1 : rdata = 43'b0001101100000001010000000010000000100000000;
			// PEs: 58, 58 -> 
			// srcs: (3, 2)(72) 1, (273) -2 --> (473) -2:ND2, NW2, *, 
			8'd2 : rdata = 43'b0001101100000010010000000100000000000000000;
			// PEs: 57, 58 -> 
			// srcs: (11, 3)(668) 2, (473) -2 --> (669) 0:PENB, ALU, +, 
			8'd3 : rdata = 43'b0000111011111110001111111110000000000000000;
			// PEs: 57, 58 -> 62
			// srcs: (33, 4)(667) 3, (669) 0 --> (670) 3:PENB, ALU, +, PEGB6
			8'd4 : rdata = 43'b0000111011111110001111111110000000011100000;
			// PEs: 58, 57 -> 57
			// srcs: (268, 8)(3) 1, (875) 0 --> (1075) 0:NM0, PENB, *, PEGB1
			8'd5 : rdata = 43'b0001110000000000110111111100000000010010000;
			// PEs: 58, 57 -> 57
			// srcs: (270, 9)(3) 1, (877) 0 --> (1077) 0:NM0, PENB, *, PEGB1
			8'd6 : rdata = 43'b0001110000000000110111111100000000010010000;
			// PEs: 56, 58 -> 58
			// srcs: (271, 5)(809) 0, (72) 1 --> (878) 0:PEGB0, ND2, *, NI0
			8'd7 : rdata = 43'b0001111100000000011000000101000000000000000;
			// PEs: 56, 58 -> 59
			// srcs: (272, 6)(809) 0, (73) -3 --> (879) 0:PEGB0, ND0, *, PENB
			8'd8 : rdata = 43'b0001111100000000011000000000000000100000000;
			// PEs: 58, 58 -> 
			// srcs: (274, 10)(3) 1, (878) 0 --> (1078) 0:NM0, NI0, *, 
			8'd9 : rdata = 43'b0001110000000000101000000000000000000000000;
			// PEs: 58, 58 -> 58
			// srcs: (277, 12)(273) -2, (1078) 0 --> (1278) -2:NW2, ALU, -, NW2
			8'd10 : rdata = 43'b0001001000000010001111111110001100000000000;
			// PEs: 58, 59 -> 58
			// srcs: (281, 13)(274) -2, (1079) 0 --> (1279) -2:NW0, PEGB3, -, NW0
			8'd11 : rdata = 43'b0001001000000000111000001100001000000000000;
			// PEs: 58, 57 -> 57
			// srcs: (348, 11)(3) 1, (955) 0 --> (1155) 0:NM0, PENB, *, PEGB1
			8'd12 : rdata = 43'b0001110000000000110111111100000000010010000;
			// PEs: 56, 58 -> 59
			// srcs: (350, 7)(809) 0, (151) 2 --> (957) 0:PEGB0, ND1, *, PENB
			8'd13 : rdata = 43'b0001111100000000011000000010000000100000000;
			// PEs: 58, 59 -> 58
			// srcs: (359, 14)(352) -1, (1157) 0 --> (1357) -1:NW1, PEGB3, -, NW1
			8'd14 : rdata = 43'b0001001000000001111000001100001010000000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 59) begin
	always @(*) begin
		case(address)
			// PEs: 59, 59 -> 59
			// srcs: (1, 0)(74) -1, (275) 0 --> (475) 0:ND0, NW0, *, NI0
			8'd0 : rdata = 43'b0001101100000000010000000001000000000000000;
			// PEs: 59, 59 -> 59
			// srcs: (2, 1)(152) -3, (353) -3 --> (553) 9:ND1, NW1, *, NI1
			8'd1 : rdata = 43'b0001101100000001010000000011010000000000000;
			// PEs: 59, 59 -> 59
			// srcs: (3, 2)(75) 2, (276) 2 --> (476) 4:ND2, NW2, *, NI2
			8'd2 : rdata = 43'b0001101100000010010000000101100000000000000;
			// PEs: 58, 59 -> 60
			// srcs: (4, 3)(474) 6, (475) 0 --> (671) 6:PENB, NI0, +, PENB
			8'd3 : rdata = 43'b0000111011111110101000000000000000100000000;
			// PEs: 58, 59 -> 56
			// srcs: (5, 4)(552) -2, (553) 9 --> (747) 7:PENB, NI1, +, PEGB0
			8'd4 : rdata = 43'b0000111011111110101000000010000000010000000;
			// PEs: 59 -> 60
			// srcs: (11, 5)(476) 4 --> (476) 4:NI2, pass, PENB
			8'd5 : rdata = 43'b1100010100000010000000000000000000100000000;
			// PEs: 56, 59 -> 60
			// srcs: (273, 6)(809) 0, (74) -1 --> (880) 0:PEGB0, ND0, *, PENB
			8'd6 : rdata = 43'b0001111100000000011000000000000000100000000;
			// PEs: 56, 59 -> 59
			// srcs: (274, 7)(809) 0, (75) 2 --> (881) 0:PEGB0, ND2, *, NI0
			8'd7 : rdata = 43'b0001111100000000011000000101000000000000000;
			// PEs: 59, 58 -> 58
			// srcs: (275, 9)(3) 1, (879) 0 --> (1079) 0:NM0, PENB, *, PEGB2
			8'd8 : rdata = 43'b0001110000000000110111111100000000010100000;
			// PEs: 59, 59 -> 
			// srcs: (277, 10)(3) 1, (881) 0 --> (1081) 0:NM0, NI0, *, 
			8'd9 : rdata = 43'b0001110000000000101000000000000000000000000;
			// PEs: 59, 59 -> 59
			// srcs: (280, 13)(276) 2, (1081) 0 --> (1281) 2:NW2, ALU, -, NW2
			8'd10 : rdata = 43'b0001001000000010001111111110001100000000000;
			// PEs: 59, 60 -> 59
			// srcs: (282, 12)(275) 0, (1080) 0 --> (1280) 0:NW0, PEGB4, -, NW0
			8'd11 : rdata = 43'b0001001000000000111000010000001000000000000;
			// PEs: 56, 59 -> 60
			// srcs: (351, 8)(809) 0, (152) -3 --> (958) 0:PEGB0, ND1, *, PENB
			8'd12 : rdata = 43'b0001111100000000011000000010000000100000000;
			// PEs: 59, 58 -> 58
			// srcs: (353, 11)(3) 1, (957) 0 --> (1157) 0:NM0, PENB, *, PEGB2
			8'd13 : rdata = 43'b0001110000000000110111111100000000010100000;
			// PEs: 59, 60 -> 59
			// srcs: (360, 14)(353) -3, (1158) 0 --> (1358) -3:NW1, PEGB4, -, NW1
			8'd14 : rdata = 43'b0001001000000001111000010000001010000000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 60) begin
	always @(*) begin
		case(address)
			// PEs: 60, 60 -> 61
			// srcs: (1, 0)(76) 0, (277) -1 --> (477) 0:ND0, NW0, *, PENB
			8'd0 : rdata = 43'b0001101100000000010000000000000000100000000;
			// PEs: 60, 60 -> 61
			// srcs: (2, 1)(154) 2, (355) 2 --> (555) 4:ND1, NW1, *, PENB
			8'd1 : rdata = 43'b0001101100000001010000000010000000100000000;
			// PEs: 60, 60 -> 61
			// srcs: (3, 2)(78) -2, (279) 0 --> (479) 0:ND2, NW2, *, PENB
			8'd2 : rdata = 43'b0001101100000010010000000100000000100000000;
			// PEs: 59 -> 
			// srcs: (6, 3)(671) 6 --> (671) 6:PENB, pass, 
			8'd3 : rdata = 43'b1100011011111110000000000000000000000000000;
			// PEs: 60, 59 -> 61
			// srcs: (13, 4)(671) 6, (476) 4 --> (672) 10:ALU, PENB, +, PENB
			8'd4 : rdata = 43'b0000100111111111110111111100000000100000000;
			// PEs: 56, 60 -> 60
			// srcs: (275, 5)(809) 0, (76) 0 --> (882) 0:PEGB0, ND0, *, NI0
			8'd5 : rdata = 43'b0001111100000000011000000001000000000000000;
			// PEs: 60, 59 -> 59
			// srcs: (276, 8)(3) 1, (880) 0 --> (1080) 0:NM0, PENB, *, PEGB3
			8'd6 : rdata = 43'b0001110000000000110111111100000000010110000;
			// PEs: 56, 60 -> 60
			// srcs: (277, 6)(809) 0, (78) -2 --> (884) 0:PEGB0, ND2, *, NI1
			8'd7 : rdata = 43'b0001111100000000011000000101010000000000000;
			// PEs: 60, 60 -> 60
			// srcs: (278, 9)(3) 1, (882) 0 --> (1082) 0:NM0, NI0, *, NI2
			8'd8 : rdata = 43'b0001110000000000101000000001100000000000000;
			// PEs: 60, 60 -> 60
			// srcs: (280, 10)(3) 1, (884) 0 --> (1084) 0:NM0, NI1, *, NI0
			8'd9 : rdata = 43'b0001110000000000101000000011000000000000000;
			// PEs: 60, 60 -> 60
			// srcs: (281, 12)(277) -1, (1082) 0 --> (1282) -1:NW0, NI2, -, NW0
			8'd10 : rdata = 43'b0001001000000000101000000100001000000000000;
			// PEs: 60, 60 -> 60
			// srcs: (283, 13)(279) 0, (1084) 0 --> (1284) 0:NW2, NI0, -, NW2
			8'd11 : rdata = 43'b0001001000000010101000000000001100000000000;
			// PEs: 56, 60 -> 61
			// srcs: (353, 7)(809) 0, (154) 2 --> (960) 0:PEGB0, ND1, *, PENB
			8'd12 : rdata = 43'b0001111100000000011000000010000000100000000;
			// PEs: 60, 59 -> 59
			// srcs: (354, 11)(3) 1, (958) 0 --> (1158) 0:NM0, PENB, *, PEGB3
			8'd13 : rdata = 43'b0001110000000000110111111100000000010110000;
			// PEs: 60, 61 -> 60
			// srcs: (362, 14)(355) 2, (1160) 0 --> (1360) 2:NW1, PEGB5, -, NW1
			8'd14 : rdata = 43'b0001001000000001111000010100001010000000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 61) begin
	always @(*) begin
		case(address)
			// PEs: 61, 61 -> 61
			// srcs: (1, 0)(77) -3, (278) 1 --> (478) -3:ND0, NW0, *, NI0
			8'd0 : rdata = 43'b0001101100000000010000000001000000000000000;
			// PEs: 61, 61 -> 61
			// srcs: (2, 1)(155) -3, (356) -2 --> (556) 6:ND1, NW1, *, NI1
			8'd1 : rdata = 43'b0001101100000001010000000011010000000000000;
			// PEs: 61, 61 -> 56
			// srcs: (3, 2)(85) -2, (286) -3 --> (486) 6:ND2, NW2, *, PEGB0
			8'd2 : rdata = 43'b0001101100000010010000000100000000010000000;
			// PEs: 60, 61 -> 61
			// srcs: (4, 3)(477) 0, (478) -3 --> (673) -3:PENB, NI0, +, NI2
			8'd3 : rdata = 43'b0000111011111110101000000001100000000000000;
			// PEs: 60, 61 -> 62
			// srcs: (5, 4)(555) 4, (556) 6 --> (753) 10:PENB, NI1, +, PENB
			8'd4 : rdata = 43'b0000111011111110101000000010000000100000000;
			// PEs: 61, 60 -> 
			// srcs: (7, 5)(673) -3, (479) 0 --> (674) -3:NI2, PENB, +, 
			8'd5 : rdata = 43'b0000110100000010110111111100000000000000000;
			// PEs: 60, 61 -> 62
			// srcs: (16, 6)(672) 10, (674) -3 --> (675) 7:PENB, ALU, +, PENB
			8'd6 : rdata = 43'b0000111011111110001111111110000000100000000;
			// PEs: 56, 61 -> 62
			// srcs: (276, 7)(809) 0, (77) -3 --> (883) 0:PEGB0, ND0, *, PENB
			8'd7 : rdata = 43'b0001111100000000011000000000000000100000000;
			// PEs: 56, 61 -> 61
			// srcs: (284, 8)(809) 0, (85) -2 --> (891) 0:PEGB0, ND2, *, NI0
			8'd8 : rdata = 43'b0001111100000000011000000101000000000000000;
			// PEs: 61, 62 -> 61
			// srcs: (285, 12)(278) 1, (1083) 0 --> (1283) 1:NW0, PEGB6, -, NW0
			8'd9 : rdata = 43'b0001001000000000111000011000001000000000000;
			// PEs: 61, 61 -> 
			// srcs: (287, 10)(3) 1, (891) 0 --> (1091) 0:NM0, NI0, *, 
			8'd10 : rdata = 43'b0001110000000000101000000000000000000000000;
			// PEs: 61, 61 -> 61
			// srcs: (290, 13)(286) -3, (1091) 0 --> (1291) -3:NW2, ALU, -, NW2
			8'd11 : rdata = 43'b0001001000000010001111111110001100000000000;
			// PEs: 56, 61 -> 62
			// srcs: (354, 9)(809) 0, (155) -3 --> (961) 0:PEGB0, ND1, *, PENB
			8'd12 : rdata = 43'b0001111100000000011000000010000000100000000;
			// PEs: 61, 60 -> 60
			// srcs: (356, 11)(3) 1, (960) 0 --> (1160) 0:NM0, PENB, *, PEGB4
			8'd13 : rdata = 43'b0001110000000000110111111100000000011000000;
			// PEs: 61, 62 -> 61
			// srcs: (363, 14)(356) -2, (1161) 0 --> (1361) -2:NW1, PEGB6, -, NW1
			8'd14 : rdata = 43'b0001001000000001111000011000001010000000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 62) begin
	always @(*) begin
		case(address)
			// PEs: 62, 62 -> 63
			// srcs: (1, 0)(79) -2, (280) 2 --> (480) -4:ND0, NW0, *, PENB
			8'd0 : rdata = 43'b0001101100000000010000000000000000100000000;
			// PEs: 62, 62 -> 63
			// srcs: (2, 1)(156) -2, (357) -3 --> (557) 6:ND1, NW1, *, PENB
			8'd1 : rdata = 43'b0001101100000001010000000010000000100000000;
			// PEs: 62, 62 -> 56
			// srcs: (3, 2)(88) 2, (289) -3 --> (489) -6:ND2, NW2, *, PEGB0
			8'd2 : rdata = 43'b0001101100000010010000000100000000010000000;
			// PEs: 61, 63 -> 56
			// srcs: (11, 3)(753) 10, (754) 6 --> (755) 16:PENB, PEGB7, +, PEGB0
			8'd3 : rdata = 43'b0000111011111110111000011100000000010000000;
			// PEs: 58, 61 -> 57
			// srcs: (39, 4)(670) 3, (675) 7 --> (676) 10:PEGB2, PENB, +, PEGB1
			8'd4 : rdata = 43'b0000111100000100110111111100000000010010000;
			// PEs: 56, 62 -> 62
			// srcs: (278, 5)(809) 0, (79) -2 --> (885) 0:PEGB0, ND0, *, NI0
			8'd5 : rdata = 43'b0001111100000000011000000001000000000000000;
			// PEs: 62, 61 -> 61
			// srcs: (279, 8)(3) 1, (883) 0 --> (1083) 0:NM0, PENB, *, PEGB5
			8'd6 : rdata = 43'b0001110000000000110111111100000000011010000;
			// PEs: 62, 62 -> 
			// srcs: (281, 9)(3) 1, (885) 0 --> (1085) 0:NM0, NI0, *, 
			8'd7 : rdata = 43'b0001110000000000101000000000000000000000000;
			// PEs: 62, 62 -> 62
			// srcs: (284, 12)(280) 2, (1085) 0 --> (1285) 2:NW0, ALU, -, NW0
			8'd8 : rdata = 43'b0001001000000000001111111110001000000000000;
			// PEs: 56, 62 -> 
			// srcs: (287, 6)(809) 0, (88) 2 --> (894) 0:PEGB0, ND2, *, 
			8'd9 : rdata = 43'b0001111100000000011000000100000000000000000;
			// PEs: 62, 62 -> 
			// srcs: (290, 10)(3) 1, (894) 0 --> (1094) 0:NM0, ALU, *, 
			8'd10 : rdata = 43'b0001110000000000001111111110000000000000000;
			// PEs: 62, 62 -> 62
			// srcs: (293, 13)(289) -3, (1094) 0 --> (1294) -3:NW2, ALU, -, NW2
			8'd11 : rdata = 43'b0001001000000010001111111110001100000000000;
			// PEs: 56, 62 -> 63
			// srcs: (355, 7)(809) 0, (156) -2 --> (962) 0:PEGB0, ND1, *, PENB
			8'd12 : rdata = 43'b0001111100000000011000000010000000100000000;
			// PEs: 62, 61 -> 61
			// srcs: (357, 11)(3) 1, (961) 0 --> (1161) 0:NM0, PENB, *, PEGB5
			8'd13 : rdata = 43'b0001110000000000110111111100000000011010000;
			// PEs: 62, 63 -> 62
			// srcs: (364, 14)(357) -3, (1162) 0 --> (1362) -3:NW1, PEGB7, -, NW1
			8'd14 : rdata = 43'b0001001000000001111000011100001010000000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 63) begin
	always @(*) begin
		case(address)
			// PEs: 63, 63 -> 63
			// srcs: (1, 0)(80) -1, (281) -3 --> (481) 3:ND0, NW0, *, NI0
			8'd0 : rdata = 43'b0001101100000000010000000001000000000000000;
			// PEs: 63, 63 -> 63
			// srcs: (2, 1)(157) 0, (358) -3 --> (558) 0:ND1, NW1, *, NI1
			8'd1 : rdata = 43'b0001101100000001010000000011010000000000000;
			// PEs: 63, 63 -> 63
			// srcs: (3, 2)(91) -2, (292) -1 --> (492) 2:ND2, NW2, *, NI2
			8'd2 : rdata = 43'b0001101100000010010000000101100000000000000;
			// PEs: 62, 63 -> 56
			// srcs: (4, 3)(480) -4, (481) 3 --> (678) -1:PENB, NI0, +, PENB
			8'd3 : rdata = 43'b0000111011111110101000000000000000100000000;
			// PEs: 62, 63 -> 62
			// srcs: (5, 4)(557) 6, (558) 0 --> (754) 6:PENB, NI1, +, PEGB6
			8'd4 : rdata = 43'b0000111011111110101000000010000000011100000;
			// PEs: 63 -> 56
			// srcs: (12, 5)(492) 2 --> (492) 2:NI2, pass, PENB
			8'd5 : rdata = 43'b1100010100000010000000000000000000100000000;
			// PEs: 56, 63 -> 
			// srcs: (279, 6)(809) 0, (80) -1 --> (886) 0:PEGB0, ND0, *, 
			8'd6 : rdata = 43'b0001111100000000011000000000000000000000000;
			// PEs: 63, 63 -> 
			// srcs: (282, 9)(3) 1, (886) 0 --> (1086) 0:NM0, ALU, *, 
			8'd7 : rdata = 43'b0001110000000000001111111110000000000000000;
			// PEs: 63, 63 -> 63
			// srcs: (285, 13)(281) -3, (1086) 0 --> (1286) -3:NW0, ALU, -, NW0
			8'd8 : rdata = 43'b0001001000000000001111111110001000000000000;
			// PEs: 56, 63 -> 
			// srcs: (290, 7)(809) 0, (91) -2 --> (897) 0:PEGB0, ND2, *, 
			8'd9 : rdata = 43'b0001111100000000011000000100000000000000000;
			// PEs: 63, 63 -> 
			// srcs: (293, 10)(3) 1, (897) 0 --> (1097) 0:NM0, ALU, *, 
			8'd10 : rdata = 43'b0001110000000000001111111110000000000000000;
			// PEs: 63, 63 -> 63
			// srcs: (296, 14)(292) -1, (1097) 0 --> (1297) -1:NW2, ALU, -, NW2
			8'd11 : rdata = 43'b0001001000000010001111111110001100000000000;
			// PEs: 56, 63 -> 63
			// srcs: (356, 8)(809) 0, (157) 0 --> (963) 0:PEGB0, ND1, *, NI0
			8'd12 : rdata = 43'b0001111100000000011000000011000000000000000;
			// PEs: 63, 62 -> 62
			// srcs: (358, 11)(3) 1, (962) 0 --> (1162) 0:NM0, PENB, *, PEGB6
			8'd13 : rdata = 43'b0001110000000000110111111100000000011100000;
			// PEs: 63, 63 -> 
			// srcs: (359, 12)(3) 1, (963) 0 --> (1163) 0:NM0, NI0, *, 
			8'd14 : rdata = 43'b0001110000000000101000000000000000000000000;
			// PEs: 63, 63 -> 63
			// srcs: (362, 15)(358) -3, (1163) 0 --> (1363) -3:NW1, ALU, -, NW1
			8'd15 : rdata = 43'b0001001000000001001111111110001010000000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

endgenerate
/*****************************************************************************/
endmodule
