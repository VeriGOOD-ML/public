`define  `PIPE 6
`define  `SIZE 10
`define  `BITWIDTH 32
`define  `INPUT_BITWIDTH 16
