//WEIGHT_COUNT
//LANE0
`define WEIGHT_COUNT_PE_0 16'h0
`define WEIGHT_COUNT_PE_16 16'h0
`define WEIGHT_COUNT_PE_32 16'h0
`define WEIGHT_COUNT_PE_48 16'h0
`define WEIGHT_COUNT_LANE_0 16'h0
//LANE1
`define WEIGHT_COUNT_PE_1 16'he
`define WEIGHT_COUNT_PE_17 16'he
`define WEIGHT_COUNT_PE_33 16'he
`define WEIGHT_COUNT_PE_49 16'he
`define WEIGHT_COUNT_LANE_1 16'h38
//LANE2
`define WEIGHT_COUNT_PE_2 16'he
`define WEIGHT_COUNT_PE_18 16'he
`define WEIGHT_COUNT_PE_34 16'he
`define WEIGHT_COUNT_PE_50 16'he
`define WEIGHT_COUNT_LANE_2 16'h38
//LANE3
`define WEIGHT_COUNT_PE_3 16'he
`define WEIGHT_COUNT_PE_19 16'he
`define WEIGHT_COUNT_PE_35 16'he
`define WEIGHT_COUNT_PE_51 16'he
`define WEIGHT_COUNT_LANE_3 16'h38
//LANE4
`define WEIGHT_COUNT_PE_4 16'he
`define WEIGHT_COUNT_PE_20 16'he
`define WEIGHT_COUNT_PE_36 16'he
`define WEIGHT_COUNT_PE_52 16'he
`define WEIGHT_COUNT_LANE_4 16'h38
//LANE5
`define WEIGHT_COUNT_PE_5 16'he
`define WEIGHT_COUNT_PE_21 16'he
`define WEIGHT_COUNT_PE_37 16'he
`define WEIGHT_COUNT_PE_53 16'he
`define WEIGHT_COUNT_LANE_5 16'h38
//LANE6
`define WEIGHT_COUNT_PE_6 16'he
`define WEIGHT_COUNT_PE_22 16'he
`define WEIGHT_COUNT_PE_38 16'he
`define WEIGHT_COUNT_PE_54 16'he
`define WEIGHT_COUNT_LANE_6 16'h38
//LANE7
`define WEIGHT_COUNT_PE_7 16'he
`define WEIGHT_COUNT_PE_23 16'he
`define WEIGHT_COUNT_PE_39 16'he
`define WEIGHT_COUNT_PE_55 16'he
`define WEIGHT_COUNT_LANE_7 16'h38
//LANE8
`define WEIGHT_COUNT_PE_8 16'h0
`define WEIGHT_COUNT_PE_24 16'h0
`define WEIGHT_COUNT_PE_40 16'h0
`define WEIGHT_COUNT_PE_56 16'h0
`define WEIGHT_COUNT_LANE_8 16'h0
//LANE9
`define WEIGHT_COUNT_PE_9 16'he
`define WEIGHT_COUNT_PE_25 16'he
`define WEIGHT_COUNT_PE_41 16'he
`define WEIGHT_COUNT_PE_57 16'he
`define WEIGHT_COUNT_LANE_9 16'h38
//LANE10
`define WEIGHT_COUNT_PE_10 16'he
`define WEIGHT_COUNT_PE_26 16'he
`define WEIGHT_COUNT_PE_42 16'he
`define WEIGHT_COUNT_PE_58 16'he
`define WEIGHT_COUNT_LANE_10 16'h38
//LANE11
`define WEIGHT_COUNT_PE_11 16'he
`define WEIGHT_COUNT_PE_27 16'he
`define WEIGHT_COUNT_PE_43 16'he
`define WEIGHT_COUNT_PE_59 16'he
`define WEIGHT_COUNT_LANE_11 16'h38
//LANE12
`define WEIGHT_COUNT_PE_12 16'he
`define WEIGHT_COUNT_PE_28 16'he
`define WEIGHT_COUNT_PE_44 16'he
`define WEIGHT_COUNT_PE_60 16'he
`define WEIGHT_COUNT_LANE_12 16'h38
//LANE13
`define WEIGHT_COUNT_PE_13 16'he
`define WEIGHT_COUNT_PE_29 16'he
`define WEIGHT_COUNT_PE_45 16'he
`define WEIGHT_COUNT_PE_61 16'he
`define WEIGHT_COUNT_LANE_13 16'h38
//LANE14
`define WEIGHT_COUNT_PE_14 16'he
`define WEIGHT_COUNT_PE_30 16'he
`define WEIGHT_COUNT_PE_46 16'he
`define WEIGHT_COUNT_PE_62 16'he
`define WEIGHT_COUNT_LANE_14 16'h38
//LANE15
`define WEIGHT_COUNT_PE_15 16'he
`define WEIGHT_COUNT_PE_31 16'he
`define WEIGHT_COUNT_PE_47 16'he
`define WEIGHT_COUNT_PE_63 16'he
`define WEIGHT_COUNT_LANE_15 16'h38
