
`timescale 1ns/1ps
module instruction_memory #(
    parameter integer addrLen = 5,
    parameter integer dataLen = 32,
    parameter integer peId  = 1
)(
    input clk,
    input rstn,
    
    input stall,
    input start,
    input restart,
    
    output reg [dataLen - 1: 0] data_out
);
//--------------------------------------------------------------------------------------
//reg [dataLen - 1: 0] mem  [0: (1 << addrLen) - 1];
reg [addrLen-1:0]        address;
reg enable;
reg [dataLen - 1: 0] rdata;
wire end_of_instruction;
always @(posedge clk or negedge rstn)
    if(~rstn)
        enable <= 1'b0;
    else if(start)
        enable <= 1'b1;
    else if(end_of_instruction)
       enable <= 1'b0;
always @(posedge clk or negedge rstn) begin
    if(~rstn)
        address <= {addrLen{1'b0}};
    else begin
        if(end_of_instruction)
            address <= {addrLen{1'b0}};
        else if(~stall && enable )
            address <= address + {{addrLen-1{1'b0}},1'b1};   
    end     
end
always @(posedge clk or negedge rstn) begin
    if(~rstn)
        data_out <= {1'b1,{dataLen-1{1'b0}}};
    else if((~stall && enable && ~end_of_instruction)||(end_of_instruction && start))
       data_out <= rdata;
end
    
assign end_of_instruction = (data_out[dataLen-1:dataLen-5] == 5'b0);
/****************************************************************************/
generate
if(peId == 0) begin
	always @(*) begin
		case(address)
			// PEs: 7 -> 8
			// srcs: (3, 0)(412) 14 --> (412) 14:PENB, pass, PUNB
			8'd0 : rdata = 44'b11000110111111100000000000000000001000000000;
			// PEs: 7 -> 8
			// srcs: (4, 1)(490) 36 --> (490) 36:PENB, pass, PUNB
			8'd1 : rdata = 44'b11000110111111100000000000000000001000000000;
			// PEs: 7 -> 8
			// srcs: (5, 2)(568) 2 --> (568) 2:PENB, pass, PUNB
			8'd2 : rdata = 44'b11000110111111100000000000000000001000000000;
			// PEs: 7 -> 24
			// srcs: (6, 16)(517) 0 --> (517) 0:PENB, pass, PUGB3
			8'd3 : rdata = 44'b11000110111111100000000000000000000000001011;
			// PEs: 1 -> 8
			// srcs: (9, 10)(495) 4 --> (495) 4:PEGB1, pass, PUNB
			8'd4 : rdata = 44'b11000111000000100000000000000000001000000000;
			// PEs: 2 -> 8
			// srcs: (10, 11)(498) 40 --> (498) 40:PEGB2, pass, PUNB
			8'd5 : rdata = 44'b11000111000001000000000000000000001000000000;
			// PEs: 4 -> 40
			// srcs: (11, 13)(504) 5 --> (504) 5:PEGB4, pass, PUGB5
			8'd6 : rdata = 44'b11000111000010000000000000000000000000001101;
			// PEs: 5 -> 56
			// srcs: (12, 14)(511) 14 --> (511) 14:PEGB5, pass, PUGB7
			8'd7 : rdata = 44'b11000111000010100000000000000000000000001111;
			// PEs: 6 -> 16
			// srcs: (13, 15)(514) 20 --> (514) 20:PEGB6, pass, PUGB2
			8'd8 : rdata = 44'b11000111000011000000000000000000000000001010;
			// PEs: 1 -> 48
			// srcs: (14, 3)(608) 0 --> (608) 0:PEGB1, pass, PUGB6
			8'd9 : rdata = 44'b11000111000000100000000000000000000000001110;
			// PEs: 4 -> 56
			// srcs: (15, 18)(759) 57 --> (759) 57:PEGB4, pass, PUGB7
			8'd10 : rdata = 44'b11000111000010000000000000000000000000001111;
			// PEs: 40 -> 0
			// srcs: (16, 5)(436) 9 --> (436) 9:PUGB5, pass, NI0
			8'd11 : rdata = 44'b11000111000010110000000000010000000000000000;
			// PEs: 7 -> 48
			// srcs: (17, 20)(607) 74 --> (607) 74:PENB, pass, PUGB6
			8'd12 : rdata = 44'b11000110111111100000000000000000000000001110;
			// PEs: 24 -> 1
			// srcs: (19, 4)(632) 75 --> (632) 75:PUGB3, pass, PENB
			8'd13 : rdata = 44'b11000111000001110000000000000000000100000000;
			// PEs: 0 -> 1
			// srcs: (26, 6)(436) 9 --> (436) 9:NI0, pass, PENB
			8'd14 : rdata = 44'b11000101000000000000000000000000000100000000;
			// PEs: 56 -> 1
			// srcs: (27, 7)(678) 62 --> (678) 62:PUNB, pass, PENB
			8'd15 : rdata = 44'b11000110111111110000000000000000000100000000;
			// PEs: 56 -> 1
			// srcs: (28, 8)(486) 72 --> (486) 72:PUNB, pass, PENB
			8'd16 : rdata = 44'b11000110111111110000000000000000000100000000;
			// PEs: 56 -> 1
			// srcs: (29, 9)(489) 32 --> (489) 32:PUNB, pass, PENB
			8'd17 : rdata = 44'b11000110111111110000000000000000000100000000;
			// PEs: 8 -> 1
			// srcs: (30, 12)(695) 65 --> (695) 65:PUGB1, pass, PENB
			8'd18 : rdata = 44'b11000111000000110000000000000000000100000000;
			// PEs: 16 -> 1
			// srcs: (31, 17)(561) 18 --> (561) 18:PUGB2, pass, PENB
			8'd19 : rdata = 44'b11000111000001010000000000000000000100000000;
			// PEs: 1 -> 48
			// srcs: (33, 21)(633) 84 --> (633) 84:PEGB1, pass, PUGB6
			8'd20 : rdata = 44'b11000111000000100000000000000000000000001110;
			// PEs: 1 -> 8
			// srcs: (36, 25)(685) 58 --> (685) 58:PEGB1, pass, PUNB
			8'd21 : rdata = 44'b11000111000000100000000000000000001000000000;
			// PEs: 1 -> 16
			// srcs: (37, 26)(696) 77 --> (696) 77:PEGB1, pass, PUGB2
			8'd22 : rdata = 44'b11000111000000100000000000000000000000001010;
			// PEs: 2 -> 8
			// srcs: (44, 30)(683) 297 --> (683) 297:PEGB2, pass, PUNB
			8'd23 : rdata = 44'b11000111000001000000000000000000001000000000;
			// PEs: 16 -> 1
			// srcs: (47, 19)(567) 7 --> (567) 7:PUGB2, pass, PENB
			8'd24 : rdata = 44'b11000111000001010000000000000000000100000000;
			// PEs: 16 -> 0
			// srcs: (48, 22)(642) 81 --> (642) 81:PUGB2, pass, NI0
			8'd25 : rdata = 44'b11000111000001010000000000010000000000000000;
			// PEs: 48 -> 1
			// srcs: (49, 23)(644) 99 --> (644) 99:PUGB6, pass, PENB
			8'd26 : rdata = 44'b11000111000011010000000000000000000100000000;
			// PEs: 0 -> 1
			// srcs: (55, 24)(642) 81 --> (642) 81:NI0, pass, PENB
			8'd27 : rdata = 44'b11000101000000000000000000000000000100000000;
			// PEs: 56 -> 1
			// srcs: (56, 27)(755) 48 --> (755) 48:PUNB, pass, PENB
			8'd28 : rdata = 44'b11000110111111110000000000000000000100000000;
			// PEs: 1 -> 48
			// srcs: (62, 29)(645) 180 --> (645) 180:PEGB1, pass, PUGB6
			8'd29 : rdata = 44'b11000111000000100000000000000000000000001110;
			// PEs: 56 -> 1
			// srcs: (65, 28)(760) 57 --> (760) 57:PUNB, pass, PENB
			8'd30 : rdata = 44'b11000110111111110000000000000000000100000000;
			// PEs: 32 -> 1
			// srcs: (106, 31)(775) 272 --> (775) 272:PUGB4, pass, PENB
			8'd31 : rdata = 44'b11000111000010010000000000000000000100000000;
			// PEs: 1 -> 48
			// srcs: (114, 32)(776) 448 --> (776) 448:PEGB1, pass, PUGB6
			8'd32 : rdata = 44'b11000111000000100000000000000000000000001110;
			// PEs: 24 -> 0
			// srcs: (146, 33)(703) 2052 --> (703) 2052:PUGB3, pass, NI0
			8'd33 : rdata = 44'b11000111000001110000000000010000000000000000;
			// PEs: 48 -> 1
			// srcs: (149, 34)(802) 2056 --> (802) 2056:PUGB6, pass, PENB
			8'd34 : rdata = 44'b11000111000011010000000000000000000100000000;
			// PEs: 0 -> 1
			// srcs: (156, 35)(703) 2052 --> (703) 2052:NI0, pass, PENB
			8'd35 : rdata = 44'b11000101000000000000000000000000000100000000;
			// PEs: 2 -> 32
			// srcs: (175, 36)(805) -9 --> (805) -9:PEGB2, pass, PUGB4
			8'd36 : rdata = 44'b11000111000001000000000000000000000000001100;
			// PEs: 2 -> 8
			// srcs: (177, 37)(805) -9 --> (805) -9:PEGB2, pass, PUNB
			8'd37 : rdata = 44'b11000111000001000000000000000000001000000000;
			// PEs: 2 -> 32
			// srcs: (178, 38)(805) -9 --> (805) -9:PEGB2, pass, PUGB4
			8'd38 : rdata = 44'b11000111000001000000000000000000000000001100;
			// PEs: 2 -> 8
			// srcs: (179, 39)(805) -9 --> (805) -9:PEGB2, pass, PUNB
			8'd39 : rdata = 44'b11000111000001000000000000000000001000000000;
			// PEs: 2 -> 8
			// srcs: (180, 40)(805) -9 --> (805) -9:PEGB2, pass, PUNB
			8'd40 : rdata = 44'b11000111000001000000000000000000001000000000;
			// PEs: 2 -> 32
			// srcs: (181, 41)(805) -9 --> (805) -9:PEGB2, pass, PUGB4
			8'd41 : rdata = 44'b11000111000001000000000000000000000000001100;
			// PEs: 2 -> 8
			// srcs: (182, 42)(805) -9 --> (805) -9:PEGB2, pass, PUNB
			8'd42 : rdata = 44'b11000111000001000000000000000000001000000000;
			// PEs: 2 -> 8
			// srcs: (183, 43)(805) -9 --> (805) -9:PEGB2, pass, PUNB
			8'd43 : rdata = 44'b11000111000001000000000000000000001000000000;
			// PEs: 2 -> 40
			// srcs: (184, 44)(805) -9 --> (805) -9:PEGB2, pass, PUGB5
			8'd44 : rdata = 44'b11000111000001000000000000000000000000001101;
			// PEs: 2 -> 8
			// srcs: (185, 45)(805) -9 --> (805) -9:PEGB2, pass, PUNB
			8'd45 : rdata = 44'b11000111000001000000000000000000001000000000;
			// PEs: 2 -> 8
			// srcs: (186, 46)(805) -9 --> (805) -9:PEGB2, pass, PUNB
			8'd46 : rdata = 44'b11000111000001000000000000000000001000000000;
			// PEs: 2 -> 40
			// srcs: (187, 47)(805) -9 --> (805) -9:PEGB2, pass, PUGB5
			8'd47 : rdata = 44'b11000111000001000000000000000000000000001101;
			// PEs: 2 -> 16
			// srcs: (188, 48)(805) -9 --> (805) -9:PEGB2, pass, PUGB2
			8'd48 : rdata = 44'b11000111000001000000000000000000000000001010;
			// PEs: 2 -> 16
			// srcs: (189, 49)(805) -9 --> (805) -9:PEGB2, pass, PUGB2
			8'd49 : rdata = 44'b11000111000001000000000000000000000000001010;
			// PEs: 2 -> 40
			// srcs: (190, 50)(805) -9 --> (805) -9:PEGB2, pass, PUGB5
			8'd50 : rdata = 44'b11000111000001000000000000000000000000001101;
			// PEs: 2 -> 16
			// srcs: (191, 51)(805) -9 --> (805) -9:PEGB2, pass, PUGB2
			8'd51 : rdata = 44'b11000111000001000000000000000000000000001010;
			// PEs: 2 -> 16
			// srcs: (192, 52)(805) -9 --> (805) -9:PEGB2, pass, PUGB2
			8'd52 : rdata = 44'b11000111000001000000000000000000000000001010;
			// PEs: 2 -> 40
			// srcs: (193, 53)(805) -9 --> (805) -9:PEGB2, pass, PUGB5
			8'd53 : rdata = 44'b11000111000001000000000000000000000000001101;
			// PEs: 2 -> 16
			// srcs: (194, 54)(805) -9 --> (805) -9:PEGB2, pass, PUGB2
			8'd54 : rdata = 44'b11000111000001000000000000000000000000001010;
			// PEs: 2 -> 16
			// srcs: (195, 55)(805) -9 --> (805) -9:PEGB2, pass, PUGB2
			8'd55 : rdata = 44'b11000111000001000000000000000000000000001010;
			// PEs: 2 -> 16
			// srcs: (196, 56)(805) -9 --> (805) -9:PEGB2, pass, PUGB2
			8'd56 : rdata = 44'b11000111000001000000000000000000000000001010;
			// PEs: 2 -> 24
			// srcs: (197, 57)(805) -9 --> (805) -9:PEGB2, pass, PUGB3
			8'd57 : rdata = 44'b11000111000001000000000000000000000000001011;
			// PEs: 2 -> 24
			// srcs: (198, 58)(805) -9 --> (805) -9:PEGB2, pass, PUGB3
			8'd58 : rdata = 44'b11000111000001000000000000000000000000001011;
			// PEs: 2 -> 24
			// srcs: (199, 59)(805) -9 --> (805) -9:PEGB2, pass, PUGB3
			8'd59 : rdata = 44'b11000111000001000000000000000000000000001011;
			// PEs: 2 -> 40
			// srcs: (200, 60)(805) -9 --> (805) -9:PEGB2, pass, PUGB5
			8'd60 : rdata = 44'b11000111000001000000000000000000000000001101;
			// PEs: 2 -> 24
			// srcs: (201, 61)(805) -9 --> (805) -9:PEGB2, pass, PUGB3
			8'd61 : rdata = 44'b11000111000001000000000000000000000000001011;
			// PEs: 2 -> 24
			// srcs: (202, 62)(805) -9 --> (805) -9:PEGB2, pass, PUGB3
			8'd62 : rdata = 44'b11000111000001000000000000000000000000001011;
			// PEs: 2 -> 40
			// srcs: (203, 63)(805) -9 --> (805) -9:PEGB2, pass, PUGB5
			8'd63 : rdata = 44'b11000111000001000000000000000000000000001101;
			// PEs: 2 -> 24
			// srcs: (204, 64)(805) -9 --> (805) -9:PEGB2, pass, PUGB3
			8'd64 : rdata = 44'b11000111000001000000000000000000000000001011;
			// PEs: 2 -> 24
			// srcs: (205, 65)(805) -9 --> (805) -9:PEGB2, pass, PUGB3
			8'd65 : rdata = 44'b11000111000001000000000000000000000000001011;
			// PEs: 2 -> 40
			// srcs: (206, 66)(805) -9 --> (805) -9:PEGB2, pass, PUGB5
			8'd66 : rdata = 44'b11000111000001000000000000000000000000001101;
			// PEs: 2 -> 32
			// srcs: (207, 67)(805) -9 --> (805) -9:PEGB2, pass, PUGB4
			8'd67 : rdata = 44'b11000111000001000000000000000000000000001100;
			// PEs: 2 -> 32
			// srcs: (208, 68)(805) -9 --> (805) -9:PEGB2, pass, PUGB4
			8'd68 : rdata = 44'b11000111000001000000000000000000000000001100;
			// PEs: 2 -> 48
			// srcs: (209, 69)(805) -9 --> (805) -9:PEGB2, pass, PUGB6
			8'd69 : rdata = 44'b11000111000001000000000000000000000000001110;
			// PEs: 2 -> 32
			// srcs: (210, 70)(805) -9 --> (805) -9:PEGB2, pass, PUGB4
			8'd70 : rdata = 44'b11000111000001000000000000000000000000001100;
			// PEs: 2 -> 32
			// srcs: (211, 71)(805) -9 --> (805) -9:PEGB2, pass, PUGB4
			8'd71 : rdata = 44'b11000111000001000000000000000000000000001100;
			// PEs: 2 -> 48
			// srcs: (212, 72)(805) -9 --> (805) -9:PEGB2, pass, PUGB6
			8'd72 : rdata = 44'b11000111000001000000000000000000000000001110;
			// PEs: 2 -> 32
			// srcs: (213, 73)(805) -9 --> (805) -9:PEGB2, pass, PUGB4
			8'd73 : rdata = 44'b11000111000001000000000000000000000000001100;
			// PEs: 2 -> 32
			// srcs: (214, 74)(805) -9 --> (805) -9:PEGB2, pass, PUGB4
			8'd74 : rdata = 44'b11000111000001000000000000000000000000001100;
			// PEs: 2 -> 48
			// srcs: (215, 75)(805) -9 --> (805) -9:PEGB2, pass, PUGB6
			8'd75 : rdata = 44'b11000111000001000000000000000000000000001110;
			// PEs: 2 -> 32
			// srcs: (216, 76)(805) -9 --> (805) -9:PEGB2, pass, PUGB4
			8'd76 : rdata = 44'b11000111000001000000000000000000000000001100;
			// PEs: 2 -> 40
			// srcs: (217, 77)(805) -9 --> (805) -9:PEGB2, pass, PUGB5
			8'd77 : rdata = 44'b11000111000001000000000000000000000000001101;
			// PEs: 2 -> 48
			// srcs: (218, 78)(805) -9 --> (805) -9:PEGB2, pass, PUGB6
			8'd78 : rdata = 44'b11000111000001000000000000000000000000001110;
			// PEs: 2 -> 40
			// srcs: (219, 79)(805) -9 --> (805) -9:PEGB2, pass, PUGB5
			8'd79 : rdata = 44'b11000111000001000000000000000000000000001101;
			// PEs: 2 -> 40
			// srcs: (220, 80)(805) -9 --> (805) -9:PEGB2, pass, PUGB5
			8'd80 : rdata = 44'b11000111000001000000000000000000000000001101;
			// PEs: 2 -> 40
			// srcs: (221, 81)(805) -9 --> (805) -9:PEGB2, pass, PUGB5
			8'd81 : rdata = 44'b11000111000001000000000000000000000000001101;
			// PEs: 2 -> 40
			// srcs: (222, 82)(805) -9 --> (805) -9:PEGB2, pass, PUGB5
			8'd82 : rdata = 44'b11000111000001000000000000000000000000001101;
			// PEs: 2 -> 40
			// srcs: (223, 83)(805) -9 --> (805) -9:PEGB2, pass, PUGB5
			8'd83 : rdata = 44'b11000111000001000000000000000000000000001101;
			// PEs: 2 -> 40
			// srcs: (224, 84)(805) -9 --> (805) -9:PEGB2, pass, PUGB5
			8'd84 : rdata = 44'b11000111000001000000000000000000000000001101;
			// PEs: 2 -> 48
			// srcs: (225, 85)(805) -9 --> (805) -9:PEGB2, pass, PUGB6
			8'd85 : rdata = 44'b11000111000001000000000000000000000000001110;
			// PEs: 2 -> 48
			// srcs: (226, 86)(805) -9 --> (805) -9:PEGB2, pass, PUGB6
			8'd86 : rdata = 44'b11000111000001000000000000000000000000001110;
			// PEs: 2 -> 48
			// srcs: (227, 87)(805) -9 --> (805) -9:PEGB2, pass, PUGB6
			8'd87 : rdata = 44'b11000111000001000000000000000000000000001110;
			// PEs: 2 -> 48
			// srcs: (228, 88)(805) -9 --> (805) -9:PEGB2, pass, PUGB6
			8'd88 : rdata = 44'b11000111000001000000000000000000000000001110;
			// PEs: 2 -> 48
			// srcs: (229, 89)(805) -9 --> (805) -9:PEGB2, pass, PUGB6
			8'd89 : rdata = 44'b11000111000001000000000000000000000000001110;
			// PEs: 2 -> 48
			// srcs: (230, 90)(805) -9 --> (805) -9:PEGB2, pass, PUGB6
			8'd90 : rdata = 44'b11000111000001000000000000000000000000001110;
			// PEs: 2 -> 48
			// srcs: (231, 91)(805) -9 --> (805) -9:PEGB2, pass, PUGB6
			8'd91 : rdata = 44'b11000111000001000000000000000000000000001110;
			// PEs: 2 -> 48
			// srcs: (232, 92)(805) -9 --> (805) -9:PEGB2, pass, PUGB6
			8'd92 : rdata = 44'b11000111000001000000000000000000000000001110;
			// PEs: 2 -> 48
			// srcs: (233, 93)(805) -9 --> (805) -9:PEGB2, pass, PUGB6
			8'd93 : rdata = 44'b11000111000001000000000000000000000000001110;
			// PEs: 2 -> 56
			// srcs: (234, 94)(805) -9 --> (805) -9:PEGB2, pass, PUGB7
			8'd94 : rdata = 44'b11000111000001000000000000000000000000001111;
			// PEs: 2 -> 48
			// srcs: (235, 95)(805) -9 --> (805) -9:PEGB2, pass, PUGB6
			8'd95 : rdata = 44'b11000111000001000000000000000000000000001110;
			// PEs: 2 -> 56
			// srcs: (236, 96)(805) -9 --> (805) -9:PEGB2, pass, PUGB7
			8'd96 : rdata = 44'b11000111000001000000000000000000000000001111;
			// PEs: 2 -> 56
			// srcs: (237, 97)(805) -9 --> (805) -9:PEGB2, pass, PUGB7
			8'd97 : rdata = 44'b11000111000001000000000000000000000000001111;
			// PEs: 2 -> 56
			// srcs: (238, 98)(805) -9 --> (805) -9:PEGB2, pass, PUGB7
			8'd98 : rdata = 44'b11000111000001000000000000000000000000001111;
			// PEs: 2 -> 56
			// srcs: (239, 99)(805) -9 --> (805) -9:PEGB2, pass, PUGB7
			8'd99 : rdata = 44'b11000111000001000000000000000000000000001111;
			// PEs: 2 -> 56
			// srcs: (240, 100)(805) -9 --> (805) -9:PEGB2, pass, PUGB7
			8'd100 : rdata = 44'b11000111000001000000000000000000000000001111;
			// PEs: 2 -> 56
			// srcs: (241, 101)(805) -9 --> (805) -9:PEGB2, pass, PUGB7
			8'd101 : rdata = 44'b11000111000001000000000000000000000000001111;
			// PEs: 2 -> 56
			// srcs: (242, 102)(805) -9 --> (805) -9:PEGB2, pass, PUGB7
			8'd102 : rdata = 44'b11000111000001000000000000000000000000001111;
			// PEs: 2 -> 56
			// srcs: (243, 103)(805) -9 --> (805) -9:PEGB2, pass, PUGB7
			8'd103 : rdata = 44'b11000111000001000000000000000000000000001111;
			// PEs: 2 -> 56
			// srcs: (244, 104)(805) -9 --> (805) -9:PEGB2, pass, PUGB7
			8'd104 : rdata = 44'b11000111000001000000000000000000000000001111;
			// PEs: 2 -> 56
			// srcs: (245, 105)(805) -9 --> (805) -9:PEGB2, pass, PUGB7
			8'd105 : rdata = 44'b11000111000001000000000000000000000000001111;
			// PEs: 2 -> 56
			// srcs: (250, 106)(805) -9 --> (805) -9:PEGB2, pass, PUGB7
			8'd106 : rdata = 44'b11000111000001000000000000000000000000001111;
			// PEs: 2 -> 56
			// srcs: (253, 107)(805) -9 --> (805) -9:PEGB2, pass, PUGB7
			8'd107 : rdata = 44'b11000111000001000000000000000000000000001111;
			// PEs: 2 -> 8
			// srcs: (255, 108)(805) -9 --> (805) -9:PEGB2, pass, PUNB
			8'd108 : rdata = 44'b11000111000001000000000000000000001000000000;
			// PEs: 2 -> 56
			// srcs: (256, 109)(805) -9 --> (805) -9:PEGB2, pass, PUGB7
			8'd109 : rdata = 44'b11000111000001000000000000000000000000001111;
			// PEs: 2 -> 8
			// srcs: (257, 110)(805) -9 --> (805) -9:PEGB2, pass, PUNB
			8'd110 : rdata = 44'b11000111000001000000000000000000001000000000;
			// PEs: 2 -> 8
			// srcs: (258, 111)(805) -9 --> (805) -9:PEGB2, pass, PUNB
			8'd111 : rdata = 44'b11000111000001000000000000000000001000000000;
			// PEs: 2 -> 8
			// srcs: (260, 112)(805) -9 --> (805) -9:PEGB2, pass, PUNB
			8'd112 : rdata = 44'b11000111000001000000000000000000001000000000;
			// PEs: 2 -> 8
			// srcs: (261, 113)(805) -9 --> (805) -9:PEGB2, pass, PUNB
			8'd113 : rdata = 44'b11000111000001000000000000000000001000000000;
			// PEs: 2 -> 8
			// srcs: (263, 114)(805) -9 --> (805) -9:PEGB2, pass, PUNB
			8'd114 : rdata = 44'b11000111000001000000000000000000001000000000;
			// PEs: 2 -> 8
			// srcs: (264, 115)(805) -9 --> (805) -9:PEGB2, pass, PUNB
			8'd115 : rdata = 44'b11000111000001000000000000000000001000000000;
			// PEs: 2 -> 16
			// srcs: (266, 116)(805) -9 --> (805) -9:PEGB2, pass, PUGB2
			8'd116 : rdata = 44'b11000111000001000000000000000000000000001010;
			// PEs: 2 -> 16
			// srcs: (267, 117)(805) -9 --> (805) -9:PEGB2, pass, PUGB2
			8'd117 : rdata = 44'b11000111000001000000000000000000000000001010;
			// PEs: 2 -> 16
			// srcs: (269, 118)(805) -9 --> (805) -9:PEGB2, pass, PUGB2
			8'd118 : rdata = 44'b11000111000001000000000000000000000000001010;
			// PEs: 2 -> 16
			// srcs: (270, 119)(805) -9 --> (805) -9:PEGB2, pass, PUGB2
			8'd119 : rdata = 44'b11000111000001000000000000000000000000001010;
			// PEs: 2 -> 16
			// srcs: (271, 120)(805) -9 --> (805) -9:PEGB2, pass, PUGB2
			8'd120 : rdata = 44'b11000111000001000000000000000000000000001010;
			// PEs: 2 -> 16
			// srcs: (272, 121)(805) -9 --> (805) -9:PEGB2, pass, PUGB2
			8'd121 : rdata = 44'b11000111000001000000000000000000000000001010;
			// PEs: 2 -> 16
			// srcs: (273, 122)(805) -9 --> (805) -9:PEGB2, pass, PUGB2
			8'd122 : rdata = 44'b11000111000001000000000000000000000000001010;
			// PEs: 2 -> 24
			// srcs: (274, 123)(805) -9 --> (805) -9:PEGB2, pass, PUGB3
			8'd123 : rdata = 44'b11000111000001000000000000000000000000001011;
			// PEs: 2 -> 24
			// srcs: (276, 124)(805) -9 --> (805) -9:PEGB2, pass, PUGB3
			8'd124 : rdata = 44'b11000111000001000000000000000000000000001011;
			// PEs: 2 -> 24
			// srcs: (277, 125)(805) -9 --> (805) -9:PEGB2, pass, PUGB3
			8'd125 : rdata = 44'b11000111000001000000000000000000000000001011;
			// PEs: 2 -> 24
			// srcs: (279, 126)(805) -9 --> (805) -9:PEGB2, pass, PUGB3
			8'd126 : rdata = 44'b11000111000001000000000000000000000000001011;
			// PEs: 2 -> 24
			// srcs: (280, 127)(805) -9 --> (805) -9:PEGB2, pass, PUGB3
			8'd127 : rdata = 44'b11000111000001000000000000000000000000001011;
			// PEs: 2 -> 24
			// srcs: (282, 128)(805) -9 --> (805) -9:PEGB2, pass, PUGB3
			8'd128 : rdata = 44'b11000111000001000000000000000000000000001011;
			// PEs: 2 -> 24
			// srcs: (283, 129)(805) -9 --> (805) -9:PEGB2, pass, PUGB3
			8'd129 : rdata = 44'b11000111000001000000000000000000000000001011;
			// PEs: 2 -> 8
			// srcs: (284, 130)(805) -9 --> (805) -9:PEGB2, pass, PUNB
			8'd130 : rdata = 44'b11000111000001000000000000000000001000000000;
			// PEs: 2 -> 32
			// srcs: (285, 131)(805) -9 --> (805) -9:PEGB2, pass, PUGB4
			8'd131 : rdata = 44'b11000111000001000000000000000000000000001100;
			// PEs: 2 -> 32
			// srcs: (286, 132)(805) -9 --> (805) -9:PEGB2, pass, PUGB4
			8'd132 : rdata = 44'b11000111000001000000000000000000000000001100;
			// PEs: 2 -> 8
			// srcs: (287, 133)(805) -9 --> (805) -9:PEGB2, pass, PUNB
			8'd133 : rdata = 44'b11000111000001000000000000000000001000000000;
			// PEs: 2 -> 32
			// srcs: (288, 134)(805) -9 --> (805) -9:PEGB2, pass, PUGB4
			8'd134 : rdata = 44'b11000111000001000000000000000000000000001100;
			// PEs: 2 -> 32
			// srcs: (289, 135)(805) -9 --> (805) -9:PEGB2, pass, PUGB4
			8'd135 : rdata = 44'b11000111000001000000000000000000000000001100;
			// PEs: 2 -> 8
			// srcs: (290, 136)(805) -9 --> (805) -9:PEGB2, pass, PUNB
			8'd136 : rdata = 44'b11000111000001000000000000000000001000000000;
			// PEs: 2 -> 32
			// srcs: (291, 137)(805) -9 --> (805) -9:PEGB2, pass, PUGB4
			8'd137 : rdata = 44'b11000111000001000000000000000000000000001100;
			// PEs: 2 -> 32
			// srcs: (292, 138)(805) -9 --> (805) -9:PEGB2, pass, PUGB4
			8'd138 : rdata = 44'b11000111000001000000000000000000000000001100;
			// PEs: 2 -> 8
			// srcs: (293, 139)(805) -9 --> (805) -9:PEGB2, pass, PUNB
			8'd139 : rdata = 44'b11000111000001000000000000000000001000000000;
			// PEs: 2 -> 32
			// srcs: (294, 140)(805) -9 --> (805) -9:PEGB2, pass, PUGB4
			8'd140 : rdata = 44'b11000111000001000000000000000000000000001100;
			// PEs: 2 -> 40
			// srcs: (295, 141)(805) -9 --> (805) -9:PEGB2, pass, PUGB5
			8'd141 : rdata = 44'b11000111000001000000000000000000000000001101;
			// PEs: 2 -> 40
			// srcs: (296, 142)(805) -9 --> (805) -9:PEGB2, pass, PUGB5
			8'd142 : rdata = 44'b11000111000001000000000000000000000000001101;
			// PEs: 2 -> 40
			// srcs: (297, 143)(805) -9 --> (805) -9:PEGB2, pass, PUGB5
			8'd143 : rdata = 44'b11000111000001000000000000000000000000001101;
			// PEs: 2 -> 40
			// srcs: (298, 144)(805) -9 --> (805) -9:PEGB2, pass, PUGB5
			8'd144 : rdata = 44'b11000111000001000000000000000000000000001101;
			// PEs: 2 -> 40
			// srcs: (299, 145)(805) -9 --> (805) -9:PEGB2, pass, PUGB5
			8'd145 : rdata = 44'b11000111000001000000000000000000000000001101;
			// PEs: 2 -> 8
			// srcs: (300, 146)(805) -9 --> (805) -9:PEGB2, pass, PUNB
			8'd146 : rdata = 44'b11000111000001000000000000000000001000000000;
			// PEs: 2 -> 40
			// srcs: (301, 147)(805) -9 --> (805) -9:PEGB2, pass, PUGB5
			8'd147 : rdata = 44'b11000111000001000000000000000000000000001101;
			// PEs: 2 -> 40
			// srcs: (302, 148)(805) -9 --> (805) -9:PEGB2, pass, PUGB5
			8'd148 : rdata = 44'b11000111000001000000000000000000000000001101;
			// PEs: 2 -> 8
			// srcs: (303, 149)(805) -9 --> (805) -9:PEGB2, pass, PUNB
			8'd149 : rdata = 44'b11000111000001000000000000000000001000000000;
			// PEs: 2 -> 48
			// srcs: (304, 150)(805) -9 --> (805) -9:PEGB2, pass, PUGB6
			8'd150 : rdata = 44'b11000111000001000000000000000000000000001110;
			// PEs: 2 -> 48
			// srcs: (305, 151)(805) -9 --> (805) -9:PEGB2, pass, PUGB6
			8'd151 : rdata = 44'b11000111000001000000000000000000000000001110;
			// PEs: 2 -> 8
			// srcs: (306, 152)(805) -9 --> (805) -9:PEGB2, pass, PUNB
			8'd152 : rdata = 44'b11000111000001000000000000000000001000000000;
			// PEs: 2 -> 48
			// srcs: (307, 153)(805) -9 --> (805) -9:PEGB2, pass, PUGB6
			8'd153 : rdata = 44'b11000111000001000000000000000000000000001110;
			// PEs: 2 -> 48
			// srcs: (308, 154)(805) -9 --> (805) -9:PEGB2, pass, PUGB6
			8'd154 : rdata = 44'b11000111000001000000000000000000000000001110;
			// PEs: 2 -> 16
			// srcs: (309, 155)(805) -9 --> (805) -9:PEGB2, pass, PUGB2
			8'd155 : rdata = 44'b11000111000001000000000000000000000000001010;
			// PEs: 2 -> 48
			// srcs: (310, 156)(805) -9 --> (805) -9:PEGB2, pass, PUGB6
			8'd156 : rdata = 44'b11000111000001000000000000000000000000001110;
			// PEs: 2 -> 48
			// srcs: (311, 157)(805) -9 --> (805) -9:PEGB2, pass, PUGB6
			8'd157 : rdata = 44'b11000111000001000000000000000000000000001110;
			// PEs: 2 -> 16
			// srcs: (312, 158)(805) -9 --> (805) -9:PEGB2, pass, PUGB2
			8'd158 : rdata = 44'b11000111000001000000000000000000000000001010;
			// PEs: 2 -> 48
			// srcs: (313, 159)(805) -9 --> (805) -9:PEGB2, pass, PUGB6
			8'd159 : rdata = 44'b11000111000001000000000000000000000000001110;
			// PEs: 2 -> 56
			// srcs: (314, 160)(805) -9 --> (805) -9:PEGB2, pass, PUGB7
			8'd160 : rdata = 44'b11000111000001000000000000000000000000001111;
			// PEs: 2 -> 16
			// srcs: (315, 161)(805) -9 --> (805) -9:PEGB2, pass, PUGB2
			8'd161 : rdata = 44'b11000111000001000000000000000000000000001010;
			// PEs: 2 -> 56
			// srcs: (316, 162)(805) -9 --> (805) -9:PEGB2, pass, PUGB7
			8'd162 : rdata = 44'b11000111000001000000000000000000000000001111;
			// PEs: 2 -> 56
			// srcs: (317, 163)(805) -9 --> (805) -9:PEGB2, pass, PUGB7
			8'd163 : rdata = 44'b11000111000001000000000000000000000000001111;
			// PEs: 2 -> 16
			// srcs: (318, 164)(805) -9 --> (805) -9:PEGB2, pass, PUGB2
			8'd164 : rdata = 44'b11000111000001000000000000000000000000001010;
			// PEs: 2 -> 56
			// srcs: (319, 165)(805) -9 --> (805) -9:PEGB2, pass, PUGB7
			8'd165 : rdata = 44'b11000111000001000000000000000000000000001111;
			// PEs: 2 -> 56
			// srcs: (320, 166)(805) -9 --> (805) -9:PEGB2, pass, PUGB7
			8'd166 : rdata = 44'b11000111000001000000000000000000000000001111;
			// PEs: 2 -> 56
			// srcs: (321, 167)(805) -9 --> (805) -9:PEGB2, pass, PUGB7
			8'd167 : rdata = 44'b11000111000001000000000000000000000000001111;
			// PEs: 2 -> 56
			// srcs: (322, 168)(805) -9 --> (805) -9:PEGB2, pass, PUGB7
			8'd168 : rdata = 44'b11000111000001000000000000000000000000001111;
			// PEs: 2 -> 16
			// srcs: (325, 169)(805) -9 --> (805) -9:PEGB2, pass, PUGB2
			8'd169 : rdata = 44'b11000111000001000000000000000000000000001010;
			// PEs: 2 -> 16
			// srcs: (328, 170)(805) -9 --> (805) -9:PEGB2, pass, PUGB2
			8'd170 : rdata = 44'b11000111000001000000000000000000000000001010;
			// PEs: 2 -> 16
			// srcs: (331, 171)(805) -9 --> (805) -9:PEGB2, pass, PUGB2
			8'd171 : rdata = 44'b11000111000001000000000000000000000000001010;
			// PEs: 2 -> 8
			// srcs: (333, 172)(805) -9 --> (805) -9:PEGB2, pass, PUNB
			8'd172 : rdata = 44'b11000111000001000000000000000000001000000000;
			// PEs: 2 -> 24
			// srcs: (334, 173)(805) -9 --> (805) -9:PEGB2, pass, PUGB3
			8'd173 : rdata = 44'b11000111000001000000000000000000000000001011;
			// PEs: 2 -> 8
			// srcs: (335, 174)(805) -9 --> (805) -9:PEGB2, pass, PUNB
			8'd174 : rdata = 44'b11000111000001000000000000000000001000000000;
			// PEs: 2 -> 8
			// srcs: (336, 175)(805) -9 --> (805) -9:PEGB2, pass, PUNB
			8'd175 : rdata = 44'b11000111000001000000000000000000001000000000;
			// PEs: 2 -> 24
			// srcs: (337, 176)(805) -9 --> (805) -9:PEGB2, pass, PUGB3
			8'd176 : rdata = 44'b11000111000001000000000000000000000000001011;
			// PEs: 2 -> 8
			// srcs: (338, 177)(805) -9 --> (805) -9:PEGB2, pass, PUNB
			8'd177 : rdata = 44'b11000111000001000000000000000000001000000000;
			// PEs: 2 -> 8
			// srcs: (339, 178)(805) -9 --> (805) -9:PEGB2, pass, PUNB
			8'd178 : rdata = 44'b11000111000001000000000000000000001000000000;
			// PEs: 2 -> 24
			// srcs: (340, 179)(805) -9 --> (805) -9:PEGB2, pass, PUGB3
			8'd179 : rdata = 44'b11000111000001000000000000000000000000001011;
			// PEs: 2 -> 8
			// srcs: (341, 180)(805) -9 --> (805) -9:PEGB2, pass, PUNB
			8'd180 : rdata = 44'b11000111000001000000000000000000001000000000;
			// PEs: 2 -> 8
			// srcs: (342, 181)(805) -9 --> (805) -9:PEGB2, pass, PUNB
			8'd181 : rdata = 44'b11000111000001000000000000000000001000000000;
			// PEs: 2 -> 24
			// srcs: (343, 182)(805) -9 --> (805) -9:PEGB2, pass, PUGB3
			8'd182 : rdata = 44'b11000111000001000000000000000000000000001011;
			// PEs: 2 -> 16
			// srcs: (344, 183)(805) -9 --> (805) -9:PEGB2, pass, PUGB2
			8'd183 : rdata = 44'b11000111000001000000000000000000000000001010;
			// PEs: 2 -> 16
			// srcs: (345, 184)(805) -9 --> (805) -9:PEGB2, pass, PUGB2
			8'd184 : rdata = 44'b11000111000001000000000000000000000000001010;
			// PEs: 2 -> 16
			// srcs: (346, 185)(805) -9 --> (805) -9:PEGB2, pass, PUGB2
			8'd185 : rdata = 44'b11000111000001000000000000000000000000001010;
			// PEs: 2 -> 16
			// srcs: (347, 186)(805) -9 --> (805) -9:PEGB2, pass, PUGB2
			8'd186 : rdata = 44'b11000111000001000000000000000000000000001010;
			// PEs: 2 -> 16
			// srcs: (348, 187)(805) -9 --> (805) -9:PEGB2, pass, PUGB2
			8'd187 : rdata = 44'b11000111000001000000000000000000000000001010;
			// PEs: 2 -> 16
			// srcs: (349, 188)(805) -9 --> (805) -9:PEGB2, pass, PUGB2
			8'd188 : rdata = 44'b11000111000001000000000000000000000000001010;
			// PEs: 2 -> 24
			// srcs: (350, 189)(805) -9 --> (805) -9:PEGB2, pass, PUGB3
			8'd189 : rdata = 44'b11000111000001000000000000000000000000001011;
			// PEs: 2 -> 16
			// srcs: (351, 190)(805) -9 --> (805) -9:PEGB2, pass, PUGB2
			8'd190 : rdata = 44'b11000111000001000000000000000000000000001010;
			// PEs: 2 -> 24
			// srcs: (352, 191)(805) -9 --> (805) -9:PEGB2, pass, PUGB3
			8'd191 : rdata = 44'b11000111000001000000000000000000000000001011;
			// PEs: 2 -> 24
			// srcs: (353, 192)(805) -9 --> (805) -9:PEGB2, pass, PUGB3
			8'd192 : rdata = 44'b11000111000001000000000000000000000000001011;
			// PEs: 2 -> 24
			// srcs: (354, 193)(805) -9 --> (805) -9:PEGB2, pass, PUGB3
			8'd193 : rdata = 44'b11000111000001000000000000000000000000001011;
			// PEs: 2 -> 24
			// srcs: (355, 194)(805) -9 --> (805) -9:PEGB2, pass, PUGB3
			8'd194 : rdata = 44'b11000111000001000000000000000000000000001011;
			// PEs: 2 -> 24
			// srcs: (356, 195)(805) -9 --> (805) -9:PEGB2, pass, PUGB3
			8'd195 : rdata = 44'b11000111000001000000000000000000000000001011;
			// PEs: 2 -> 24
			// srcs: (357, 196)(805) -9 --> (805) -9:PEGB2, pass, PUGB3
			8'd196 : rdata = 44'b11000111000001000000000000000000000000001011;
			// PEs: 2 -> 24
			// srcs: (358, 197)(805) -9 --> (805) -9:PEGB2, pass, PUGB3
			8'd197 : rdata = 44'b11000111000001000000000000000000000000001011;
			// PEs: 2 -> 32
			// srcs: (359, 198)(805) -9 --> (805) -9:PEGB2, pass, PUGB4
			8'd198 : rdata = 44'b11000111000001000000000000000000000000001100;
			// PEs: 2 -> 24
			// srcs: (360, 199)(805) -9 --> (805) -9:PEGB2, pass, PUGB3
			8'd199 : rdata = 44'b11000111000001000000000000000000000000001011;
			// PEs: 2 -> 24
			// srcs: (361, 200)(805) -9 --> (805) -9:PEGB2, pass, PUGB3
			8'd200 : rdata = 44'b11000111000001000000000000000000000000001011;
			// PEs: 2 -> 32
			// srcs: (362, 201)(805) -9 --> (805) -9:PEGB2, pass, PUGB4
			8'd201 : rdata = 44'b11000111000001000000000000000000000000001100;
			// PEs: 2 -> 32
			// srcs: (363, 202)(805) -9 --> (805) -9:PEGB2, pass, PUGB4
			8'd202 : rdata = 44'b11000111000001000000000000000000000000001100;
			// PEs: 2 -> 32
			// srcs: (364, 203)(805) -9 --> (805) -9:PEGB2, pass, PUGB4
			8'd203 : rdata = 44'b11000111000001000000000000000000000000001100;
			// PEs: 2 -> 32
			// srcs: (365, 204)(805) -9 --> (805) -9:PEGB2, pass, PUGB4
			8'd204 : rdata = 44'b11000111000001000000000000000000000000001100;
			// PEs: 2 -> 32
			// srcs: (366, 205)(805) -9 --> (805) -9:PEGB2, pass, PUGB4
			8'd205 : rdata = 44'b11000111000001000000000000000000000000001100;
			// PEs: 2 -> 32
			// srcs: (367, 206)(805) -9 --> (805) -9:PEGB2, pass, PUGB4
			8'd206 : rdata = 44'b11000111000001000000000000000000000000001100;
			// PEs: 2 -> 32
			// srcs: (368, 207)(805) -9 --> (805) -9:PEGB2, pass, PUGB4
			8'd207 : rdata = 44'b11000111000001000000000000000000000000001100;
			default : rdata = 44'b00000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 1) begin
	always @(*) begin
		case(address)
			// PEs: 1, 1 -> 3
			// srcs: (1, 0)(4) 2, (205) 3 --> (405) 6:ND0, NW0, *, PEGB3
			8'd0 : rdata = 44'b00011011000000000100000000000000000010110000;
			// PEs: 1, 1 -> 2
			// srcs: (2, 1)(81) 6, (282) 8 --> (482) 48:ND1, NW1, *, PENB
			8'd1 : rdata = 44'b00011011000000010100000000100000000100000000;
			// PEs: 1, 1 -> 2
			// srcs: (3, 2)(158) 1, (359) 9 --> (559) 9:ND2, NW2, *, PENB
			8'd2 : rdata = 44'b00011011000000100100000001000000000100000000;
			// PEs: 1, 1 -> 0
			// srcs: (4, 3)(94) 1, (295) 4 --> (495) 4:ND3, NW3, *, PEGB0
			8'd3 : rdata = 44'b00011011000000110100000001100000000010000000;
			// PEs: 6 -> 
			// srcs: (6, 4)(410) 0 --> (410) 0:PEGB6, pass, 
			8'd4 : rdata = 44'b11000111000011000000000000000000000000000000;
			// PEs: 5, 1 -> 0
			// srcs: (9, 5)(409) 0, (410) 0 --> (608) 0:PEGB5, ALU, +, PEGB0
			8'd5 : rdata = 44'b00001111000010100011111111100000000010000000;
			// PEs: 0 -> 
			// srcs: (21, 6)(632) 75 --> (632) 75:PENB, pass, 
			8'd6 : rdata = 44'b11000110111111100000000000000000000000000000;
			// PEs: 1, 0 -> 0
			// srcs: (28, 7)(632) 75, (436) 9 --> (633) 84:ALU, PENB, +, PEGB0
			8'd7 : rdata = 44'b00001001111111111101111111000000000010000000;
			// PEs: 0, 2 -> 1
			// srcs: (29, 8)(678) 62, (679) 66 --> (680) 128:PENB, PEGB2, +, NI0
			8'd8 : rdata = 44'b00001110111111101110000010010000000000000000;
			// PEs: 4, 0 -> 2
			// srcs: (30, 9)(681) 97, (486) 72 --> (682) 169:PEGB4, PENB, +, PENB
			8'd9 : rdata = 44'b00001111000010001101111111000000000100000000;
			// PEs: 6, 0 -> 0
			// srcs: (31, 10)(684) 26, (489) 32 --> (685) 58:PEGB6, PENB, +, PEGB0
			8'd10 : rdata = 44'b00001111000011001101111111000000000010000000;
			// PEs: 0, 3 -> 0
			// srcs: (32, 11)(695) 65, (501) 12 --> (696) 77:PENB, PEGB3, +, PEGB0
			8'd11 : rdata = 44'b00001110111111101110000011000000000010000000;
			// PEs: 2, 0 -> 1
			// srcs: (33, 12)(756) 12, (561) 18 --> (757) 30:PEGB2, PENB, +, NI1
			8'd12 : rdata = 44'b00001111000001001101111111010100000000000000;
			// PEs: 1 -> 2
			// srcs: (37, 16)(680) 128 --> (680) 128:NI0, pass, PENB
			8'd13 : rdata = 44'b11000101000000000000000000000000000100000000;
			// PEs: 6, 0 -> 1
			// srcs: (49, 13)(761) 34, (567) 7 --> (762) 41:PEGB6, PENB, +, NI0
			8'd14 : rdata = 44'b00001111000011001101111111010000000000000000;
			// PEs: 0 -> 
			// srcs: (51, 14)(644) 99 --> (644) 99:PENB, pass, 
			8'd15 : rdata = 44'b11000110111111100000000000000000000000000000;
			// PEs: 0, 1 -> 0
			// srcs: (57, 15)(642) 81, (644) 99 --> (645) 180:PENB, ALU, +, PEGB0
			8'd16 : rdata = 44'b00001110111111100011111111100000000010000000;
			// PEs: 0, 1 -> 1
			// srcs: (58, 17)(755) 48, (757) 30 --> (758) 78:PENB, NI1, +, NI2
			8'd17 : rdata = 44'b00001110111111101010000000111000000000000000;
			// PEs: 0, 1 -> 2
			// srcs: (68, 18)(760) 57, (762) 41 --> (763) 98:PENB, NI0, +, PENB
			8'd18 : rdata = 44'b00001110111111101010000000000000000100000000;
			// PEs: 1 -> 2
			// srcs: (75, 19)(758) 78 --> (758) 78:NI2, pass, PENB
			8'd19 : rdata = 44'b11000101000000100000000000000000000100000000;
			// PEs: 2, 0 -> 0
			// srcs: (109, 20)(764) 176, (775) 272 --> (776) 448:PEGB2, PENB, +, PEGB0
			8'd20 : rdata = 44'b00001111000001001101111111000000000010000000;
			// PEs: 0 -> 
			// srcs: (151, 21)(802) 2056 --> (802) 2056:PENB, pass, 
			8'd21 : rdata = 44'b11000110111111100000000000000000000000000000;
			// PEs: 0, 1 -> 
			// srcs: (158, 22)(703) 2052, (802) 2056 --> (803) 4108:PENB, ALU, +, ALU
			8'd22 : rdata = 44'b00001110111111100011111111100000000000000000;
			// PEs: 1 -> 2
			// srcs: (159, 23)(803) 4108 --> (804) 0:ALU, sigmoid, PENB
			8'd23 : rdata = 44'b10000001111111110000000000000000000100000000;
			// PEs: 2, 1 -> 
			// srcs: (168, 24)(805) -9, (4) 2 --> (806) -18:PEGB2, ND0, *, 
			8'd24 : rdata = 44'b00011111000001000110000000000000000000000000;
			// PEs: 1, 1 -> 
			// srcs: (171, 28)(3) 1, (806) -18 --> (1006) -18:NM0, ALU, *, 
			8'd25 : rdata = 44'b00011100000000000011111111100000000000000000;
			// PEs: 1, 1 -> 1
			// srcs: (174, 32)(205) 3, (1006) -18 --> (1206) 21:NW0, ALU, -, NW0
			8'd26 : rdata = 44'b00010010000000000011111111100010000000000000;
			// PEs: 2, 1 -> 
			// srcs: (246, 25)(805) -9, (81) 6 --> (883) -54:PEGB2, ND1, *, 
			8'd27 : rdata = 44'b00011111000001000110000000100000000000000000;
			// PEs: 1, 1 -> 
			// srcs: (249, 29)(3) 1, (883) -54 --> (1083) -54:NM0, ALU, *, 
			8'd28 : rdata = 44'b00011100000000000011111111100000000000000000;
			// PEs: 1, 1 -> 1
			// srcs: (252, 33)(282) 8, (1083) -54 --> (1283) 62:NW1, ALU, -, NW1
			8'd29 : rdata = 44'b00010010000000010011111111100010010000000000;
			// PEs: 2, 1 -> 
			// srcs: (259, 26)(805) -9, (94) 1 --> (896) -9:PEGB2, ND3, *, 
			8'd30 : rdata = 44'b00011111000001000110000001100000000000000000;
			// PEs: 1, 1 -> 
			// srcs: (262, 30)(3) 1, (896) -9 --> (1096) -9:NM0, ALU, *, 
			8'd31 : rdata = 44'b00011100000000000011111111100000000000000000;
			// PEs: 1, 1 -> 1
			// srcs: (265, 34)(295) 4, (1096) -9 --> (1296) 13:NW3, ALU, -, NW3
			8'd32 : rdata = 44'b00010010000000110011111111100010110000000000;
			// PEs: 2, 1 -> 
			// srcs: (323, 27)(805) -9, (158) 1 --> (960) -9:PEGB2, ND2, *, 
			8'd33 : rdata = 44'b00011111000001000110000001000000000000000000;
			// PEs: 1, 1 -> 
			// srcs: (326, 31)(3) 1, (960) -9 --> (1160) -9:NM0, ALU, *, 
			8'd34 : rdata = 44'b00011100000000000011111111100000000000000000;
			// PEs: 1, 1 -> 1
			// srcs: (329, 35)(359) 9, (1160) -9 --> (1360) 18:NW2, ALU, -, NW2
			8'd35 : rdata = 44'b00010010000000100011111111100010100000000000;
			default : rdata = 44'b00000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 2) begin
	always @(*) begin
		case(address)
			// PEs: 2, 2 -> 3
			// srcs: (1, 0)(5) 2, (206) 6 --> (406) 12:ND0, NW0, *, PENB
			8'd0 : rdata = 44'b00011011000000000100000000000000000100000000;
			// PEs: 2, 2 -> 2
			// srcs: (2, 1)(82) 2, (283) 9 --> (483) 18:ND1, NW1, *, NI0
			8'd1 : rdata = 44'b00011011000000010100000000110000000000000000;
			// PEs: 2, 2 -> 2
			// srcs: (3, 2)(159) 1, (360) 3 --> (560) 3:ND2, NW2, *, NI1
			8'd2 : rdata = 44'b00011011000000100100000001010100000000000000;
			// PEs: 2, 2 -> 0
			// srcs: (4, 3)(97) 8, (298) 5 --> (498) 40:ND3, NW3, *, PEGB0
			8'd3 : rdata = 44'b00011011000000110100000001100000000010000000;
			// PEs: 1, 2 -> 1
			// srcs: (5, 5)(482) 48, (483) 18 --> (679) 66:PENB, NI0, +, PEGB1
			8'd4 : rdata = 44'b00001110111111101010000000000000000010010000;
			// PEs: 1, 2 -> 1
			// srcs: (6, 4)(559) 9, (560) 3 --> (756) 12:PENB, NI1, +, PEGB1
			8'd5 : rdata = 44'b00001110111111101010000000100000000010010000;
			// PEs: 1 -> 
			// srcs: (32, 6)(682) 169 --> (682) 169:PENB, pass, 
			8'd6 : rdata = 44'b11000110111111100000000000000000000000000000;
			// PEs: 1, 2 -> 0
			// srcs: (39, 7)(680) 128, (682) 169 --> (683) 297:PENB, ALU, +, PEGB0
			8'd7 : rdata = 44'b00001110111111100011111111100000000010000000;
			// PEs: 1 -> 
			// srcs: (70, 8)(763) 98 --> (763) 98:PENB, pass, 
			8'd8 : rdata = 44'b11000110111111100000000000000000000000000000;
			// PEs: 1, 2 -> 1
			// srcs: (77, 9)(758) 78, (763) 98 --> (764) 176:PENB, ALU, +, PEGB1
			8'd9 : rdata = 44'b00001110111111100011111111100000000010010000;
			// PEs: 1, 2 -> 3, 1, 2
			// srcs: (162, 10)(804) 0, (204) 9 --> (805) -9:PENB, ND4, -, NI0, PENB, PEGB1
			8'd10 : rdata = 44'b00010110111111100110000010010000000110010000;
			// PEs: 2 -> 4
			// srcs: (164, 12)(805) 0 --> (805) -9:ALU, pass, PEGB4
			8'd11 : rdata = 44'b11000001111111110000000000000000000011000000;
			// PEs: 2, 2 -> 3
			// srcs: (165, 11)(805) -9, (5) 2 --> (807) -18:NI0, ND0, *, PENB
			8'd12 : rdata = 44'b00011101000000000110000000000000000100000000;
			// PEs: 2 -> 5
			// srcs: (166, 13)(805) -9 --> (805) -9:NI0, pass, PEGB5
			8'd13 : rdata = 44'b11000101000000000000000000000000000011010000;
			// PEs: 2 -> 6
			// srcs: (167, 14)(805) -9 --> (805) -9:NI0, pass, PEGB6
			8'd14 : rdata = 44'b11000101000000000000000000000000000011100000;
			// PEs: 2 -> 0
			// srcs: (168, 15)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd15 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 7
			// srcs: (169, 16)(805) -9 --> (805) -9:NI0, pass, PEGB7
			8'd16 : rdata = 44'b11000101000000000000000000000000000011110000;
			// PEs: 2 -> 0
			// srcs: (170, 17)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd17 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (171, 18)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd18 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (172, 19)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd19 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (173, 20)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd20 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (174, 21)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd21 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (175, 22)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd22 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (176, 23)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd23 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (177, 24)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd24 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (178, 25)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd25 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (179, 26)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd26 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (180, 27)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd27 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (181, 28)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd28 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (182, 29)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd29 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (183, 30)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd30 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (184, 31)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd31 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (185, 32)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd32 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (186, 33)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd33 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (187, 34)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd34 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (188, 35)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd35 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (189, 36)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd36 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (190, 37)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd37 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (191, 38)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd38 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (192, 39)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd39 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (193, 40)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd40 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (194, 41)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd41 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (195, 42)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd42 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (196, 43)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd43 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (197, 44)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd44 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (198, 45)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd45 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (199, 46)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd46 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (200, 47)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd47 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (201, 48)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd48 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (202, 49)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd49 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (203, 50)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd50 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (204, 51)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd51 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (205, 52)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd52 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (206, 53)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd53 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (207, 54)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd54 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (208, 55)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd55 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (209, 56)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd56 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (210, 57)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd57 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (211, 58)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd58 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (212, 59)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd59 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (213, 60)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd60 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (214, 61)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd61 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (215, 62)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd62 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (216, 63)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd63 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (217, 64)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd64 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (218, 65)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd65 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (219, 66)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd66 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (220, 67)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd67 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (221, 68)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd68 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (222, 69)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd69 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (223, 70)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd70 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (224, 71)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd71 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (225, 72)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd72 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (226, 73)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd73 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (227, 74)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd74 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (228, 75)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd75 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (229, 76)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd76 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (230, 77)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd77 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (231, 78)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd78 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (232, 79)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd79 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (233, 80)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd80 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (234, 81)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd81 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (235, 82)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd82 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (236, 83)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd83 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (237, 84)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd84 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (238, 85)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd85 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 1
			// srcs: (239, 86)(805) -9 --> (805) -9:NI0, pass, PEGB1
			8'd86 : rdata = 44'b11000101000000000000000000000000000010010000;
			// PEs: 2, 2 -> 3
			// srcs: (240, 87)(805) -9, (82) 2 --> (884) -18:NI0, ND1, *, PENB
			8'd87 : rdata = 44'b00011101000000000110000000100000000100000000;
			// PEs: 2 -> 3
			// srcs: (241, 88)(805) -9 --> (805) -9:NI0, pass, PENB
			8'd88 : rdata = 44'b11000101000000000000000000000000000100000000;
			// PEs: 2 -> 4
			// srcs: (242, 89)(805) -9 --> (805) -9:NI0, pass, PEGB4
			8'd89 : rdata = 44'b11000101000000000000000000000000000011000000;
			// PEs: 2 -> 0
			// srcs: (243, 90)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd90 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 5
			// srcs: (244, 91)(805) -9 --> (805) -9:NI0, pass, PEGB5
			8'd91 : rdata = 44'b11000101000000000000000000000000000011010000;
			// PEs: 2 -> 6
			// srcs: (245, 92)(805) -9 --> (805) -9:NI0, pass, PEGB6
			8'd92 : rdata = 44'b11000101000000000000000000000000000011100000;
			// PEs: 2 -> 0
			// srcs: (246, 93)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd93 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 7
			// srcs: (247, 94)(805) -9 --> (805) -9:NI0, pass, PEGB7
			8'd94 : rdata = 44'b11000101000000000000000000000000000011110000;
			// PEs: 2 -> 0
			// srcs: (248, 95)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd95 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (249, 96)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd96 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (250, 97)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd97 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (251, 98)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd98 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 1
			// srcs: (252, 99)(805) -9 --> (805) -9:NI0, pass, PEGB1
			8'd99 : rdata = 44'b11000101000000000000000000000000000010010000;
			// PEs: 2 -> 0
			// srcs: (253, 100)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd100 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (254, 101)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd101 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2, 2 -> 3
			// srcs: (255, 102)(805) -9, (97) 8 --> (899) -72:NI0, ND3, *, PENB
			8'd102 : rdata = 44'b00011101000000000110000001100000000100000000;
			// PEs: 2 -> 0
			// srcs: (256, 103)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd103 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (257, 104)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd104 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 3
			// srcs: (258, 105)(805) -9 --> (805) -9:NI0, pass, PENB
			8'd105 : rdata = 44'b11000101000000000000000000000000000100000000;
			// PEs: 2 -> 0
			// srcs: (259, 106)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd106 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (260, 107)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd107 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 4
			// srcs: (261, 108)(805) -9 --> (805) -9:NI0, pass, PEGB4
			8'd108 : rdata = 44'b11000101000000000000000000000000000011000000;
			// PEs: 2 -> 0
			// srcs: (262, 109)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd109 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (263, 110)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd110 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (264, 111)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd111 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (265, 112)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd112 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (266, 113)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd113 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (267, 114)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd114 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 5
			// srcs: (268, 115)(805) -9 --> (805) -9:NI0, pass, PEGB5
			8'd115 : rdata = 44'b11000101000000000000000000000000000011010000;
			// PEs: 2 -> 0
			// srcs: (269, 116)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd116 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (270, 117)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd117 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 6
			// srcs: (271, 118)(805) -9 --> (805) -9:NI0, pass, PEGB6
			8'd118 : rdata = 44'b11000101000000000000000000000000000011100000;
			// PEs: 2 -> 0
			// srcs: (272, 119)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd119 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (273, 120)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd120 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 7
			// srcs: (274, 121)(805) -9 --> (805) -9:NI0, pass, PEGB7
			8'd121 : rdata = 44'b11000101000000000000000000000000000011110000;
			// PEs: 2 -> 0
			// srcs: (275, 122)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd122 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (276, 123)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd123 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (277, 124)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd124 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (278, 125)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd125 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (279, 126)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd126 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (280, 127)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd127 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (281, 128)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd128 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (282, 129)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd129 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (283, 130)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd130 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (284, 131)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd131 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (285, 132)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd132 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (286, 133)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd133 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (287, 134)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd134 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (288, 135)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd135 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (289, 136)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd136 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (290, 137)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd137 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (291, 138)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd138 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (292, 139)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd139 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (293, 140)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd140 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (294, 141)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd141 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (295, 142)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd142 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (296, 143)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd143 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (297, 144)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd144 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (298, 145)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd145 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (299, 146)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd146 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (300, 147)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd147 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (301, 148)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd148 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (302, 149)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd149 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (303, 150)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd150 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (304, 151)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd151 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (305, 152)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd152 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (306, 153)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd153 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (307, 154)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd154 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (308, 155)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd155 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (309, 156)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd156 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (310, 157)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd157 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (311, 158)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd158 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (312, 159)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd159 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (313, 160)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd160 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (314, 161)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd161 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (315, 162)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd162 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 1
			// srcs: (316, 163)(805) -9 --> (805) -9:NI0, pass, PEGB1
			8'd163 : rdata = 44'b11000101000000000000000000000000000010010000;
			// PEs: 2, 2 -> 3
			// srcs: (317, 164)(805) -9, (159) 1 --> (961) -9:NI0, ND2, *, PENB
			8'd164 : rdata = 44'b00011101000000000110000001000000000100000000;
			// PEs: 2 -> 0
			// srcs: (318, 165)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd165 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 3
			// srcs: (319, 166)(805) -9 --> (805) -9:NI0, pass, PENB
			8'd166 : rdata = 44'b11000101000000000000000000000000000100000000;
			// PEs: 2 -> 4
			// srcs: (320, 167)(805) -9 --> (805) -9:NI0, pass, PEGB4
			8'd167 : rdata = 44'b11000101000000000000000000000000000011000000;
			// PEs: 2 -> 0
			// srcs: (321, 168)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd168 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 5
			// srcs: (322, 169)(805) -9 --> (805) -9:NI0, pass, PEGB5
			8'd169 : rdata = 44'b11000101000000000000000000000000000011010000;
			// PEs: 2 -> 6
			// srcs: (323, 170)(805) -9 --> (805) -9:NI0, pass, PEGB6
			8'd170 : rdata = 44'b11000101000000000000000000000000000011100000;
			// PEs: 2 -> 0
			// srcs: (324, 171)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd171 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 7
			// srcs: (325, 172)(805) -9 --> (805) -9:NI0, pass, PEGB7
			8'd172 : rdata = 44'b11000101000000000000000000000000000011110000;
			// PEs: 2 -> 0
			// srcs: (326, 173)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd173 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (327, 174)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd174 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (328, 175)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd175 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (329, 176)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd176 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (330, 177)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd177 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (331, 178)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd178 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (332, 179)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd179 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (333, 180)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd180 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (334, 181)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd181 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (335, 182)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd182 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (336, 183)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd183 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (337, 184)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd184 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (338, 185)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd185 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (339, 186)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd186 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (340, 187)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd187 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (341, 188)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd188 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (342, 189)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd189 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (343, 190)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd190 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (344, 191)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd191 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (345, 192)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd192 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (346, 193)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd193 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (347, 194)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd194 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (348, 195)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd195 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (349, 196)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd196 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (350, 197)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd197 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (351, 198)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd198 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (352, 199)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd199 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (353, 200)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd200 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (354, 201)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd201 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (355, 202)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd202 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (356, 203)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd203 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (357, 204)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd204 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (358, 205)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd205 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (359, 206)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd206 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (360, 207)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd207 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (361, 208)(805) -9 --> (805) -9:NI0, pass, PEGB0
			8'd208 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 2, 3 -> 2
			// srcs: (362, 209)(206) 6, (1007) -18 --> (1207) 24:NW0, PEGB3, -, NW0
			8'd209 : rdata = 44'b00010010000000001110000011000010000000000000;
			// PEs: 2, 3 -> 2
			// srcs: (363, 210)(283) 9, (1084) -18 --> (1284) 27:NW1, PEGB3, -, NW1
			8'd210 : rdata = 44'b00010010000000011110000011000010010000000000;
			// PEs: 2, 3 -> 2
			// srcs: (364, 211)(298) 5, (1099) -72 --> (1299) 77:NW3, PEGB3, -, NW3
			8'd211 : rdata = 44'b00010010000000111110000011000010110000000000;
			// PEs: 2, 3 -> 2
			// srcs: (365, 212)(360) 3, (1161) -9 --> (1361) 12:NW2, PEGB3, -, NW2
			8'd212 : rdata = 44'b00010010000000101110000011000010100000000000;
			default : rdata = 44'b00000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 3) begin
	always @(*) begin
		case(address)
			// PEs: 3, 3 -> 5
			// srcs: (1, 0)(6) 2, (207) 4 --> (407) 8:ND0, NW0, *, PEGB5
			8'd0 : rdata = 44'b00011011000000000100000000000000000011010000;
			// PEs: 3, 3 -> 4
			// srcs: (2, 1)(83) 6, (284) 8 --> (484) 48:ND1, NW1, *, PENB
			8'd1 : rdata = 44'b00011011000000010100000000100000000100000000;
			// PEs: 3, 3 -> 4
			// srcs: (3, 2)(161) 3, (362) 7 --> (562) 21:ND2, NW2, *, PENB
			8'd2 : rdata = 44'b00011011000000100100000001000000000100000000;
			// PEs: 3, 3 -> 1
			// srcs: (4, 3)(100) 3, (301) 4 --> (501) 12:ND3, NW3, *, PEGB1
			8'd3 : rdata = 44'b00011011000000110100000001100000000010010000;
			// PEs: 1, 2 -> 7
			// srcs: (7, 4)(405) 6, (406) 12 --> (605) 18:PEGB1, PENB, +, PEGB7
			8'd4 : rdata = 44'b00001111000000101101111111000000000011110000;
			// PEs: 2, 3 -> 4
			// srcs: (165, 5)(805) -9, (6) 2 --> (808) -18:PENB, ND0, *, PENB
			8'd5 : rdata = 44'b00011110111111100110000000000000000100000000;
			// PEs: 3, 2 -> 2
			// srcs: (168, 9)(3) 1, (807) -18 --> (1007) -18:NM0, PENB, *, PEGB2
			8'd6 : rdata = 44'b00011100000000001101111111000000000010100000;
			// PEs: 3, 4 -> 3
			// srcs: (174, 14)(207) 4, (1008) -18 --> (1208) 22:NW0, PEGB4, -, NW0
			8'd7 : rdata = 44'b00010010000000001110000100000010000000000000;
			// PEs: 3, 2 -> 2
			// srcs: (243, 10)(3) 1, (884) -18 --> (1084) -18:NM0, PENB, *, PEGB2
			8'd8 : rdata = 44'b00011100000000001101111111000000000010100000;
			// PEs: 2, 3 -> 
			// srcs: (245, 6)(805) -9, (83) 6 --> (885) -54:PENB, ND1, *, 
			8'd9 : rdata = 44'b00011110111111100110000000100000000000000000;
			// PEs: 3, 3 -> 
			// srcs: (248, 11)(3) 1, (885) -54 --> (1085) -54:NM0, ALU, *, 
			8'd10 : rdata = 44'b00011100000000000011111111100000000000000000;
			// PEs: 3, 3 -> 3
			// srcs: (251, 15)(284) 8, (1085) -54 --> (1285) 62:NW1, ALU, -, NW1
			8'd11 : rdata = 44'b00010010000000010011111111100010010000000000;
			// PEs: 3, 2 -> 2
			// srcs: (258, 12)(3) 1, (899) -72 --> (1099) -72:NM0, PENB, *, PEGB2
			8'd12 : rdata = 44'b00011100000000001101111111000000000010100000;
			// PEs: 2, 3 -> 4
			// srcs: (262, 7)(805) -9, (100) 3 --> (902) -27:PENB, ND3, *, PENB
			8'd13 : rdata = 44'b00011110111111100110000001100000000100000000;
			// PEs: 3, 4 -> 3
			// srcs: (271, 16)(301) 4, (1102) -27 --> (1302) 31:NW3, PEGB4, -, NW3
			8'd14 : rdata = 44'b00010010000000111110000100000010110000000000;
			// PEs: 3, 2 -> 2
			// srcs: (320, 13)(3) 1, (961) -9 --> (1161) -9:NM0, PENB, *, PEGB2
			8'd15 : rdata = 44'b00011100000000001101111111000000000010100000;
			// PEs: 2, 3 -> 4
			// srcs: (323, 8)(805) -9, (161) 3 --> (963) -27:PENB, ND2, *, PENB
			8'd16 : rdata = 44'b00011110111111100110000001000000000100000000;
			// PEs: 3, 4 -> 3
			// srcs: (332, 17)(362) 7, (1163) -27 --> (1363) 34:NW2, PEGB4, -, NW2
			8'd17 : rdata = 44'b00010010000000101110000100000010100000000000;
			default : rdata = 44'b00000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 4) begin
	always @(*) begin
		case(address)
			// PEs: 4, 4 -> 5
			// srcs: (1, 0)(7) 8, (208) 6 --> (408) 48:ND0, NW0, *, PENB
			8'd0 : rdata = 44'b00011011000000000100000000000000000100000000;
			// PEs: 4, 4 -> 4
			// srcs: (2, 1)(84) 7, (285) 7 --> (485) 49:ND1, NW1, *, NI0
			8'd1 : rdata = 44'b00011011000000010100000000110000000000000000;
			// PEs: 4, 4 -> 4
			// srcs: (3, 2)(162) 9, (363) 4 --> (563) 36:ND2, NW2, *, NI1
			8'd2 : rdata = 44'b00011011000000100100000001010100000000000000;
			// PEs: 4, 4 -> 0
			// srcs: (4, 3)(103) 1, (304) 5 --> (504) 5:ND3, NW3, *, PEGB0
			8'd3 : rdata = 44'b00011011000000110100000001100000000010000000;
			// PEs: 3, 4 -> 1
			// srcs: (5, 4)(484) 48, (485) 49 --> (681) 97:PENB, NI0, +, PEGB1
			8'd4 : rdata = 44'b00001110111111101010000000000000000010010000;
			// PEs: 3, 4 -> 0
			// srcs: (6, 5)(562) 21, (563) 36 --> (759) 57:PENB, NI1, +, PEGB0
			8'd5 : rdata = 44'b00001110111111101010000000100000000010000000;
			// PEs: 4, 3 -> 3
			// srcs: (168, 10)(3) 1, (808) -18 --> (1008) -18:NM0, PENB, *, PEGB3
			8'd6 : rdata = 44'b00011100000000001101111111000000000010110000;
			// PEs: 2, 4 -> 5
			// srcs: (171, 6)(805) -9, (7) 8 --> (809) -72:PEGB2, ND0, *, PENB
			8'd7 : rdata = 44'b00011111000001000110000000000000000100000000;
			// PEs: 4, 5 -> 4
			// srcs: (180, 15)(208) 6, (1009) -72 --> (1209) 78:NW0, PEGB5, -, NW0
			8'd8 : rdata = 44'b00010010000000001110000101000010000000000000;
			// PEs: 2, 4 -> 
			// srcs: (249, 7)(805) -9, (84) 7 --> (886) -63:PEGB2, ND1, *, 
			8'd9 : rdata = 44'b00011111000001000110000000100000000000000000;
			// PEs: 4, 4 -> 
			// srcs: (252, 11)(3) 1, (886) -63 --> (1086) -63:NM0, ALU, *, 
			8'd10 : rdata = 44'b00011100000000000011111111100000000000000000;
			// PEs: 4, 4 -> 4
			// srcs: (255, 16)(285) 7, (1086) -63 --> (1286) 70:NW1, ALU, -, NW1
			8'd11 : rdata = 44'b00010010000000010011111111100010010000000000;
			// PEs: 4, 3 -> 3
			// srcs: (265, 12)(3) 1, (902) -27 --> (1102) -27:NM0, PENB, *, PEGB3
			8'd12 : rdata = 44'b00011100000000001101111111000000000010110000;
			// PEs: 2, 4 -> 5
			// srcs: (268, 8)(805) -9, (103) 1 --> (905) -9:PEGB2, ND3, *, PENB
			8'd13 : rdata = 44'b00011111000001000110000001100000000100000000;
			// PEs: 4, 5 -> 4
			// srcs: (277, 17)(304) 5, (1105) -9 --> (1305) 14:NW3, PEGB5, -, NW3
			8'd14 : rdata = 44'b00010010000000111110000101000010110000000000;
			// PEs: 4, 3 -> 3
			// srcs: (326, 13)(3) 1, (963) -27 --> (1163) -27:NM0, PENB, *, PEGB3
			8'd15 : rdata = 44'b00011100000000001101111111000000000010110000;
			// PEs: 2, 4 -> 
			// srcs: (327, 9)(805) -9, (162) 9 --> (964) -81:PEGB2, ND2, *, 
			8'd16 : rdata = 44'b00011111000001000110000001000000000000000000;
			// PEs: 4, 4 -> 
			// srcs: (330, 14)(3) 1, (964) -81 --> (1164) -81:NM0, ALU, *, 
			8'd17 : rdata = 44'b00011100000000000011111111100000000000000000;
			// PEs: 4, 4 -> 4
			// srcs: (333, 18)(363) 4, (1164) -81 --> (1364) 85:NW2, ALU, -, NW2
			8'd18 : rdata = 44'b00010010000000100011111111100010100000000000;
			default : rdata = 44'b00000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 5) begin
	always @(*) begin
		case(address)
			// PEs: 5, 5 -> 1
			// srcs: (1, 0)(8) 0, (209) 5 --> (409) 0:ND0, NW0, *, PEGB1
			8'd0 : rdata = 44'b00011011000000000100000000000000000010010000;
			// PEs: 5, 5 -> 6
			// srcs: (2, 1)(86) 8, (287) 2 --> (487) 16:ND1, NW1, *, PENB
			8'd1 : rdata = 44'b00011011000000010100000000100000000100000000;
			// PEs: 5, 5 -> 6
			// srcs: (3, 2)(164) 3, (365) 3 --> (565) 9:ND2, NW2, *, PENB
			8'd2 : rdata = 44'b00011011000000100100000001000000000100000000;
			// PEs: 5, 5 -> 0
			// srcs: (4, 3)(110) 7, (311) 2 --> (511) 14:ND3, NW3, *, PEGB0
			8'd3 : rdata = 44'b00011011000000110100000001100000000010000000;
			// PEs: 3, 4 -> 7
			// srcs: (7, 4)(407) 8, (408) 48 --> (606) 56:PEGB3, PENB, +, PEGB7
			8'd4 : rdata = 44'b00001111000001101101111111000000000011110000;
			// PEs: 2, 5 -> 5
			// srcs: (173, 5)(805) -9, (8) 0 --> (810) 0:PEGB2, ND0, *, NI0
			8'd5 : rdata = 44'b00011111000001000110000000010000000000000000;
			// PEs: 5, 4 -> 4
			// srcs: (174, 9)(3) 1, (809) -72 --> (1009) -72:NM0, PENB, *, PEGB4
			8'd6 : rdata = 44'b00011100000000001101111111000000000011000000;
			// PEs: 5, 5 -> 
			// srcs: (176, 10)(3) 1, (810) 0 --> (1010) 0:NM0, NI0, *, 
			8'd7 : rdata = 44'b00011100000000001010000000000000000000000000;
			// PEs: 5, 5 -> 5
			// srcs: (179, 14)(209) 5, (1010) 0 --> (1210) 5:NW0, ALU, -, NW0
			8'd8 : rdata = 44'b00010010000000000011111111100010000000000000;
			// PEs: 2, 5 -> 
			// srcs: (251, 6)(805) -9, (86) 8 --> (888) -72:PEGB2, ND1, *, 
			8'd9 : rdata = 44'b00011111000001000110000000100000000000000000;
			// PEs: 5, 5 -> 
			// srcs: (254, 11)(3) 1, (888) -72 --> (1088) -72:NM0, ALU, *, 
			8'd10 : rdata = 44'b00011100000000000011111111100000000000000000;
			// PEs: 5, 5 -> 5
			// srcs: (257, 15)(287) 2, (1088) -72 --> (1288) 74:NW1, ALU, -, NW1
			8'd11 : rdata = 44'b00010010000000010011111111100010010000000000;
			// PEs: 5, 4 -> 4
			// srcs: (271, 12)(3) 1, (905) -9 --> (1105) -9:NM0, PENB, *, PEGB4
			8'd12 : rdata = 44'b00011100000000001101111111000000000011000000;
			// PEs: 2, 5 -> 
			// srcs: (275, 7)(805) -9, (110) 7 --> (912) -63:PEGB2, ND3, *, 
			8'd13 : rdata = 44'b00011111000001000110000001100000000000000000;
			// PEs: 5, 5 -> 
			// srcs: (278, 13)(3) 1, (912) -63 --> (1112) -63:NM0, ALU, *, 
			8'd14 : rdata = 44'b00011100000000000011111111100000000000000000;
			// PEs: 5, 5 -> 5
			// srcs: (281, 16)(311) 2, (1112) -63 --> (1312) 65:NW3, ALU, -, NW3
			8'd15 : rdata = 44'b00010010000000110011111111100010110000000000;
			// PEs: 2, 5 -> 6
			// srcs: (329, 8)(805) -9, (164) 3 --> (966) -27:PEGB2, ND2, *, PENB
			8'd16 : rdata = 44'b00011111000001000110000001000000000100000000;
			// PEs: 5, 6 -> 5
			// srcs: (338, 17)(365) 3, (1166) -27 --> (1366) 30:NW2, PEGB6, -, NW2
			8'd17 : rdata = 44'b00010010000000101110000110000010100000000000;
			default : rdata = 44'b00000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 6) begin
	always @(*) begin
		case(address)
			// PEs: 6, 6 -> 1
			// srcs: (1, 0)(9) 0, (210) 3 --> (410) 0:ND0, NW0, *, PEGB1
			8'd0 : rdata = 44'b00011011000000000100000000000000000010010000;
			// PEs: 6, 6 -> 6
			// srcs: (2, 1)(87) 5, (288) 2 --> (488) 10:ND1, NW1, *, NI0
			8'd1 : rdata = 44'b00011011000000010100000000110000000000000000;
			// PEs: 6, 6 -> 6
			// srcs: (3, 2)(165) 5, (366) 5 --> (566) 25:ND2, NW2, *, NI1
			8'd2 : rdata = 44'b00011011000000100100000001010100000000000000;
			// PEs: 6, 6 -> 0
			// srcs: (4, 3)(113) 4, (314) 5 --> (514) 20:ND3, NW3, *, PEGB0
			8'd3 : rdata = 44'b00011011000000110100000001100000000010000000;
			// PEs: 5, 6 -> 1
			// srcs: (5, 4)(487) 16, (488) 10 --> (684) 26:PENB, NI0, +, PEGB1
			8'd4 : rdata = 44'b00001110111111101010000000000000000010010000;
			// PEs: 5, 6 -> 1
			// srcs: (6, 5)(565) 9, (566) 25 --> (761) 34:PENB, NI1, +, PEGB1
			8'd5 : rdata = 44'b00001110111111101010000000100000000010010000;
			// PEs: 2, 6 -> 
			// srcs: (174, 6)(805) -9, (9) 0 --> (811) 0:PEGB2, ND0, *, 
			8'd6 : rdata = 44'b00011111000001000110000000000000000000000000;
			// PEs: 6, 6 -> 
			// srcs: (177, 10)(3) 1, (811) 0 --> (1011) 0:NM0, ALU, *, 
			8'd7 : rdata = 44'b00011100000000000011111111100000000000000000;
			// PEs: 6, 6 -> 6
			// srcs: (180, 14)(210) 3, (1011) 0 --> (1211) 3:NW0, ALU, -, NW0
			8'd8 : rdata = 44'b00010010000000000011111111100010000000000000;
			// PEs: 2, 6 -> 
			// srcs: (252, 7)(805) -9, (87) 5 --> (889) -45:PEGB2, ND1, *, 
			8'd9 : rdata = 44'b00011111000001000110000000100000000000000000;
			// PEs: 6, 6 -> 
			// srcs: (255, 11)(3) 1, (889) -45 --> (1089) -45:NM0, ALU, *, 
			8'd10 : rdata = 44'b00011100000000000011111111100000000000000000;
			// PEs: 6, 6 -> 6
			// srcs: (258, 15)(288) 2, (1089) -45 --> (1289) 47:NW1, ALU, -, NW1
			8'd11 : rdata = 44'b00010010000000010011111111100010010000000000;
			// PEs: 2, 6 -> 
			// srcs: (278, 8)(805) -9, (113) 4 --> (915) -36:PEGB2, ND3, *, 
			8'd12 : rdata = 44'b00011111000001000110000001100000000000000000;
			// PEs: 6, 6 -> 
			// srcs: (281, 12)(3) 1, (915) -36 --> (1115) -36:NM0, ALU, *, 
			8'd13 : rdata = 44'b00011100000000000011111111100000000000000000;
			// PEs: 6, 6 -> 6
			// srcs: (284, 16)(314) 5, (1115) -36 --> (1315) 41:NW3, ALU, -, NW3
			8'd14 : rdata = 44'b00010010000000110011111111100010110000000000;
			// PEs: 2, 6 -> 7
			// srcs: (330, 9)(805) -9, (165) 5 --> (967) -45:PEGB2, ND2, *, PENB
			8'd15 : rdata = 44'b00011111000001000110000001000000000100000000;
			// PEs: 6, 5 -> 5
			// srcs: (332, 13)(3) 1, (966) -27 --> (1166) -27:NM0, PENB, *, PEGB5
			8'd16 : rdata = 44'b00011100000000001101111111000000000011010000;
			// PEs: 6, 7 -> 6
			// srcs: (339, 17)(366) 5, (1167) -45 --> (1367) 50:NW2, PEGB7, -, NW2
			8'd17 : rdata = 44'b00010010000000101110000111000010100000000000;
			default : rdata = 44'b00000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 7) begin
	always @(*) begin
		case(address)
			// PEs: 7, 7 -> 0
			// srcs: (1, 0)(11) 2, (212) 7 --> (412) 14:ND0, NW0, *, PENB
			8'd0 : rdata = 44'b00011011000000000100000000000000000100000000;
			// PEs: 7, 7 -> 0
			// srcs: (2, 1)(89) 4, (290) 9 --> (490) 36:ND1, NW1, *, PENB
			8'd1 : rdata = 44'b00011011000000010100000000100000000100000000;
			// PEs: 7, 7 -> 0
			// srcs: (3, 2)(167) 2, (368) 1 --> (568) 2:ND2, NW2, *, PENB
			8'd2 : rdata = 44'b00011011000000100100000001000000000100000000;
			// PEs: 7, 7 -> 0
			// srcs: (4, 3)(116) 6, (317) 0 --> (517) 0:ND3, NW3, *, PENB
			8'd3 : rdata = 44'b00011011000000110100000001100000000100000000;
			// PEs: 5 -> 
			// srcs: (12, 4)(606) 56 --> (606) 56:PEGB5, pass, 
			8'd4 : rdata = 44'b11000111000010100000000000000000000000000000;
			// PEs: 3, 7 -> 0
			// srcs: (15, 5)(605) 18, (606) 56 --> (607) 74:PEGB3, ALU, +, PENB
			8'd5 : rdata = 44'b00001111000001100011111111100000000100000000;
			// PEs: 2, 7 -> 
			// srcs: (176, 6)(805) -9, (11) 2 --> (813) -18:PEGB2, ND0, *, 
			8'd6 : rdata = 44'b00011111000001000110000000000000000000000000;
			// PEs: 7, 7 -> 
			// srcs: (179, 10)(3) 1, (813) -18 --> (1013) -18:NM0, ALU, *, 
			8'd7 : rdata = 44'b00011100000000000011111111100000000000000000;
			// PEs: 7, 7 -> 7
			// srcs: (182, 15)(212) 7, (1013) -18 --> (1213) 25:NW0, ALU, -, NW0
			8'd8 : rdata = 44'b00010010000000000011111111100010000000000000;
			// PEs: 2, 7 -> 
			// srcs: (254, 7)(805) -9, (89) 4 --> (891) -36:PEGB2, ND1, *, 
			8'd9 : rdata = 44'b00011111000001000110000000100000000000000000;
			// PEs: 7, 7 -> 
			// srcs: (257, 11)(3) 1, (891) -36 --> (1091) -36:NM0, ALU, *, 
			8'd10 : rdata = 44'b00011100000000000011111111100000000000000000;
			// PEs: 7, 7 -> 7
			// srcs: (260, 16)(290) 9, (1091) -36 --> (1291) 45:NW1, ALU, -, NW1
			8'd11 : rdata = 44'b00010010000000010011111111100010010000000000;
			// PEs: 2, 7 -> 
			// srcs: (281, 8)(805) -9, (116) 6 --> (918) -54:PEGB2, ND3, *, 
			8'd12 : rdata = 44'b00011111000001000110000001100000000000000000;
			// PEs: 7, 7 -> 
			// srcs: (284, 12)(3) 1, (918) -54 --> (1118) -54:NM0, ALU, *, 
			8'd13 : rdata = 44'b00011100000000000011111111100000000000000000;
			// PEs: 7, 7 -> 7
			// srcs: (287, 17)(317) 0, (1118) -54 --> (1318) 54:NW3, ALU, -, NW3
			8'd14 : rdata = 44'b00010010000000110011111111100010110000000000;
			// PEs: 2, 7 -> 7
			// srcs: (332, 9)(805) -9, (167) 2 --> (969) -18:PEGB2, ND2, *, NI0
			8'd15 : rdata = 44'b00011111000001000110000001010000000000000000;
			// PEs: 7, 6 -> 6
			// srcs: (333, 13)(3) 1, (967) -45 --> (1167) -45:NM0, PENB, *, PEGB6
			8'd16 : rdata = 44'b00011100000000001101111111000000000011100000;
			// PEs: 7, 7 -> 
			// srcs: (335, 14)(3) 1, (969) -18 --> (1169) -18:NM0, NI0, *, 
			8'd17 : rdata = 44'b00011100000000001010000000000000000000000000;
			// PEs: 7, 7 -> 7
			// srcs: (338, 18)(368) 1, (1169) -18 --> (1369) 19:NW2, ALU, -, NW2
			8'd18 : rdata = 44'b00010010000000100011111111100010100000000000;
			default : rdata = 44'b00000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 8) begin
	always @(*) begin
		case(address)
			// PEs: 0 -> 9
			// srcs: (5, 0)(412) 14 --> (412) 14:PUNB, pass, PENB
			8'd0 : rdata = 44'b11000110111111110000000000000000000100000000;
			// PEs: 0 -> 9
			// srcs: (6, 1)(490) 36 --> (490) 36:PUNB, pass, PENB
			8'd1 : rdata = 44'b11000110111111110000000000000000000100000000;
			// PEs: 0 -> 9
			// srcs: (7, 2)(568) 2 --> (568) 2:PUNB, pass, PENB
			8'd2 : rdata = 44'b11000110111111110000000000000000000100000000;
			// PEs: 15 -> 0
			// srcs: (8, 13)(695) 65 --> (695) 65:PENB, pass, PUGB0
			8'd3 : rdata = 44'b11000110111111100000000000000000000000001000;
			// PEs: 11 -> 24
			// srcs: (9, 16)(526) 0 --> (526) 0:PEGB3, pass, PUGB3
			8'd4 : rdata = 44'b11000111000001100000000000000000000000001011;
			// PEs: 10 -> 16
			// srcs: (12, 4)(613) 60 --> (613) 60:PEGB2, pass, PUNB
			8'd5 : rdata = 44'b11000111000001000000000000000000001000000000;
			// PEs: 9 -> 32
			// srcs: (13, 3)(611) 22 --> (611) 22:PEGB1, pass, PUGB4
			8'd6 : rdata = 44'b11000111000000100000000000000000000000001100;
			// PEs: 11 -> 32
			// srcs: (14, 5)(617) 112 --> (617) 112:PEGB3, pass, PUGB4
			8'd7 : rdata = 44'b11000111000001100000000000000000000000001100;
			// PEs: 12 -> 40
			// srcs: (15, 6)(619) 91 --> (619) 91:PEGB4, pass, PUGB5
			8'd8 : rdata = 44'b11000111000010000000000000000000000000001101;
			// PEs: 13 -> 40
			// srcs: (16, 18)(536) 9 --> (536) 9:PEGB5, pass, PUGB5
			8'd9 : rdata = 44'b11000111000010100000000000000000000000001101;
			// PEs: 15 -> 48
			// srcs: (17, 20)(542) 72 --> (542) 72:PENB, pass, PUGB6
			8'd10 : rdata = 44'b11000110111111100000000000000000000000001110;
			// PEs: 9 -> 24
			// srcs: (18, 21)(765) 2 --> (765) 2:PEGB1, pass, PUGB3
			8'd11 : rdata = 44'b11000111000000100000000000000000000000001011;
			// PEs: 14 -> 24
			// srcs: (19, 22)(767) 67 --> (767) 67:PEGB6, pass, PUGB3
			8'd12 : rdata = 44'b11000111000011000000000000000000000000001011;
			// PEs: 24 -> 8
			// srcs: (20, 7)(635) 18 --> (635) 18:PUGB3, pass, NI0
			8'd13 : rdata = 44'b11000111000001110000000000010000000000000000;
			// PEs: 40 -> 9
			// srcs: (21, 8)(439) 18 --> (439) 18:PUGB5, pass, PENB
			8'd14 : rdata = 44'b11000111000010110000000000000000000100000000;
			// PEs: 9 -> 16
			// srcs: (23, 14)(520) 7 --> (520) 7:PEGB1, pass, PUNB
			8'd15 : rdata = 44'b11000111000000100000000000000000001000000000;
			// PEs: 10 -> 32
			// srcs: (24, 15)(523) 18 --> (523) 18:PEGB2, pass, PUGB4
			8'd16 : rdata = 44'b11000111000001000000000000000000000000001100;
			// PEs: 15 -> 24
			// srcs: (26, 24)(772) 48 --> (772) 48:PENB, pass, PUGB3
			8'd17 : rdata = 44'b11000110111111100000000000000000000000001011;
			// PEs: 8 -> 9
			// srcs: (27, 9)(635) 18 --> (635) 18:NI0, pass, PENB
			8'd18 : rdata = 44'b11000101000000000000000000000000000100000000;
			// PEs: 56 -> 9
			// srcs: (28, 10)(492) 0 --> (492) 0:PUGB7, pass, PENB
			8'd19 : rdata = 44'b11000111000011110000000000000000000100000000;
			// PEs: 0 -> 9
			// srcs: (29, 11)(495) 4 --> (495) 4:PUNB, pass, PENB
			8'd20 : rdata = 44'b11000110111111110000000000000000000100000000;
			// PEs: 0 -> 9
			// srcs: (30, 12)(498) 40 --> (498) 40:PUNB, pass, PENB
			8'd21 : rdata = 44'b11000110111111110000000000000000000100000000;
			// PEs: 40 -> 9
			// srcs: (31, 19)(734) 55 --> (734) 55:PUGB5, pass, PENB
			8'd22 : rdata = 44'b11000111000010110000000000000000000100000000;
			// PEs: 12 -> 32
			// srcs: (32, 17)(529) 5 --> (529) 5:PEGB4, pass, PUGB4
			8'd23 : rdata = 44'b11000111000010000000000000000000000000001100;
			// PEs: 13 -> 32
			// srcs: (33, 23)(770) 78 --> (770) 78:PEGB5, pass, PUGB4
			8'd24 : rdata = 44'b11000111000010100000000000000000000000001100;
			// PEs: 9 -> 16
			// srcs: (38, 27)(735) 118 --> (735) 118:PEGB1, pass, PUNB
			8'd25 : rdata = 44'b11000111000000100000000000000000001000000000;
			// PEs: 10 -> 16
			// srcs: (46, 30)(694) 85 --> (694) 85:PEGB2, pass, PUNB
			8'd26 : rdata = 44'b11000111000001000000000000000000001000000000;
			// PEs: 32 -> 9
			// srcs: (47, 25)(638) 30 --> (638) 30:PUGB4, pass, PENB
			8'd27 : rdata = 44'b11000111000010010000000000000000000100000000;
			// PEs: 0 -> 9
			// srcs: (48, 26)(685) 58 --> (685) 58:PUNB, pass, PENB
			8'd28 : rdata = 44'b11000110111111110000000000000000000100000000;
			// PEs: 48 -> 9
			// srcs: (69, 28)(634) 183 --> (634) 183:PUGB6, pass, PENB
			8'd29 : rdata = 44'b11000111000011010000000000000000000100000000;
			// PEs: 0 -> 9
			// srcs: (70, 29)(683) 297 --> (683) 297:PUNB, pass, PENB
			8'd30 : rdata = 44'b11000110111111110000000000000000000100000000;
			// PEs: 40 -> 8
			// srcs: (77, 31)(616) 207 --> (616) 207:PUGB5, pass, NI0
			8'd31 : rdata = 44'b11000111000010110000000000010000000000000000;
			// PEs: 9 -> 16
			// srcs: (78, 34)(640) 249 --> (640) 249:PEGB1, pass, PUNB
			8'd32 : rdata = 44'b11000111000000100000000000000000001000000000;
			// PEs: 9 -> 16
			// srcs: (79, 35)(689) 409 --> (689) 409:PEGB1, pass, PUNB
			8'd33 : rdata = 44'b11000111000000100000000000000000001000000000;
			// PEs: 56 -> 9
			// srcs: (82, 32)(627) 316 --> (627) 316:PUGB7, pass, PENB
			8'd34 : rdata = 44'b11000111000011110000000000000000000100000000;
			// PEs: 8 -> 9
			// srcs: (89, 33)(616) 207 --> (616) 207:NI0, pass, PENB
			8'd35 : rdata = 44'b11000101000000000000000000000000000100000000;
			// PEs: 9 -> 16
			// srcs: (96, 36)(628) 523 --> (628) 523:PEGB1, pass, PUNB
			8'd36 : rdata = 44'b11000111000000100000000000000000001000000000;
			// PEs: 0 -> 9
			// srcs: (179, 37)(805) -9 --> (805) -9:PUNB, pass, PENB
			8'd37 : rdata = 44'b11000110111111110000000000000000000100000000;
			// PEs: 0 -> 10
			// srcs: (181, 38)(805) -9 --> (805) -9:PUNB, pass, PEGB2
			8'd38 : rdata = 44'b11000110111111110000000000000000000010100000;
			// PEs: 0 -> 11
			// srcs: (182, 39)(805) -9 --> (805) -9:PUNB, pass, PEGB3
			8'd39 : rdata = 44'b11000110111111110000000000000000000010110000;
			// PEs: 0 -> 12
			// srcs: (184, 40)(805) -9 --> (805) -9:PUNB, pass, PEGB4
			8'd40 : rdata = 44'b11000110111111110000000000000000000011000000;
			// PEs: 0 -> 13
			// srcs: (185, 41)(805) -9 --> (805) -9:PUNB, pass, PEGB5
			8'd41 : rdata = 44'b11000110111111110000000000000000000011010000;
			// PEs: 0 -> 14
			// srcs: (187, 42)(805) -9 --> (805) -9:PUNB, pass, PEGB6
			8'd42 : rdata = 44'b11000110111111110000000000000000000011100000;
			// PEs: 0 -> 15
			// srcs: (188, 43)(805) -9 --> (805) -9:PUNB, pass, PEGB7
			8'd43 : rdata = 44'b11000110111111110000000000000000000011110000;
			// PEs: 0 -> 9
			// srcs: (257, 44)(805) -9 --> (805) -9:PUNB, pass, PENB
			8'd44 : rdata = 44'b11000110111111110000000000000000000100000000;
			// PEs: 0 -> 10
			// srcs: (259, 45)(805) -9 --> (805) -9:PUNB, pass, PEGB2
			8'd45 : rdata = 44'b11000110111111110000000000000000000010100000;
			// PEs: 0 -> 11
			// srcs: (260, 46)(805) -9 --> (805) -9:PUNB, pass, PEGB3
			8'd46 : rdata = 44'b11000110111111110000000000000000000010110000;
			// PEs: 0 -> 12
			// srcs: (262, 47)(805) -9 --> (805) -9:PUNB, pass, PEGB4
			8'd47 : rdata = 44'b11000110111111110000000000000000000011000000;
			// PEs: 0 -> 13
			// srcs: (263, 48)(805) -9 --> (805) -9:PUNB, pass, PEGB5
			8'd48 : rdata = 44'b11000110111111110000000000000000000011010000;
			// PEs: 0 -> 14
			// srcs: (265, 49)(805) -9 --> (805) -9:PUNB, pass, PEGB6
			8'd49 : rdata = 44'b11000110111111110000000000000000000011100000;
			// PEs: 0 -> 15
			// srcs: (266, 50)(805) -9 --> (805) -9:PUNB, pass, PEGB7
			8'd50 : rdata = 44'b11000110111111110000000000000000000011110000;
			// PEs: 0 -> 9
			// srcs: (286, 51)(805) -9 --> (805) -9:PUNB, pass, PENB
			8'd51 : rdata = 44'b11000110111111110000000000000000000100000000;
			// PEs: 0 -> 10
			// srcs: (289, 52)(805) -9 --> (805) -9:PUNB, pass, PEGB2
			8'd52 : rdata = 44'b11000110111111110000000000000000000010100000;
			// PEs: 0 -> 11
			// srcs: (292, 53)(805) -9 --> (805) -9:PUNB, pass, PEGB3
			8'd53 : rdata = 44'b11000110111111110000000000000000000010110000;
			// PEs: 0 -> 12
			// srcs: (295, 54)(805) -9 --> (805) -9:PUNB, pass, PEGB4
			8'd54 : rdata = 44'b11000110111111110000000000000000000011000000;
			// PEs: 0 -> 13
			// srcs: (302, 55)(805) -9 --> (805) -9:PUNB, pass, PEGB5
			8'd55 : rdata = 44'b11000110111111110000000000000000000011010000;
			// PEs: 0 -> 14
			// srcs: (305, 56)(805) -9 --> (805) -9:PUNB, pass, PEGB6
			8'd56 : rdata = 44'b11000110111111110000000000000000000011100000;
			// PEs: 0 -> 15
			// srcs: (308, 57)(805) -9 --> (805) -9:PUNB, pass, PEGB7
			8'd57 : rdata = 44'b11000110111111110000000000000000000011110000;
			// PEs: 0 -> 9
			// srcs: (335, 58)(805) -9 --> (805) -9:PUNB, pass, PENB
			8'd58 : rdata = 44'b11000110111111110000000000000000000100000000;
			// PEs: 0 -> 10
			// srcs: (337, 59)(805) -9 --> (805) -9:PUNB, pass, PEGB2
			8'd59 : rdata = 44'b11000110111111110000000000000000000010100000;
			// PEs: 0 -> 11
			// srcs: (338, 60)(805) -9 --> (805) -9:PUNB, pass, PEGB3
			8'd60 : rdata = 44'b11000110111111110000000000000000000010110000;
			// PEs: 0 -> 12
			// srcs: (340, 61)(805) -9 --> (805) -9:PUNB, pass, PEGB4
			8'd61 : rdata = 44'b11000110111111110000000000000000000011000000;
			// PEs: 0 -> 13
			// srcs: (341, 62)(805) -9 --> (805) -9:PUNB, pass, PEGB5
			8'd62 : rdata = 44'b11000110111111110000000000000000000011010000;
			// PEs: 0 -> 14
			// srcs: (343, 63)(805) -9 --> (805) -9:PUNB, pass, PEGB6
			8'd63 : rdata = 44'b11000110111111110000000000000000000011100000;
			// PEs: 0 -> 15
			// srcs: (344, 64)(805) -9 --> (805) -9:PUNB, pass, PEGB7
			8'd64 : rdata = 44'b11000110111111110000000000000000000011110000;
			default : rdata = 44'b00000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 9) begin
	always @(*) begin
		case(address)
			// PEs: 9, 9 -> 9
			// srcs: (1, 0)(12) 1, (213) 8 --> (413) 8:ND0, NW0, *, NI0
			8'd0 : rdata = 44'b00011011000000000100000000010000000000000000;
			// PEs: 9, 9 -> 9
			// srcs: (2, 1)(90) 2, (291) 9 --> (491) 18:ND1, NW1, *, NI1
			8'd1 : rdata = 44'b00011011000000010100000000110100000000000000;
			// PEs: 9, 9 -> 9
			// srcs: (3, 2)(168) 2, (369) 0 --> (569) 0:ND2, NW2, *, NI2
			8'd2 : rdata = 44'b00011011000000100100000001011000000000000000;
			// PEs: 9, 9 -> 9
			// srcs: (4, 3)(119) 7, (320) 1 --> (520) 7:ND3, NW3, *, NI3
			8'd3 : rdata = 44'b00011011000000110100000001111100000000000000;
			// PEs: 8, 9 -> 8
			// srcs: (8, 4)(412) 14, (413) 8 --> (611) 22:PENB, NI0, +, PEGB0
			8'd4 : rdata = 44'b00001110111111101010000000000000000010000000;
			// PEs: 8, 9 -> 9
			// srcs: (9, 5)(490) 36, (491) 18 --> (686) 54:PENB, NI1, +, NI0
			8'd5 : rdata = 44'b00001110111111101010000000110000000000000000;
			// PEs: 8, 9 -> 8
			// srcs: (10, 6)(568) 2, (569) 0 --> (765) 2:PENB, NI2, +, PEGB0
			8'd6 : rdata = 44'b00001110111111101010000001000000000010000000;
			// PEs: 9 -> 8
			// srcs: (18, 12)(520) 7 --> (520) 7:NI3, pass, PEGB0
			8'd7 : rdata = 44'b11000101000000110000000000000000000010000000;
			// PEs: 8 -> 
			// srcs: (23, 7)(439) 18 --> (439) 18:PENB, pass, 
			8'd8 : rdata = 44'b11000110111111100000000000000000000000000000;
			// PEs: 8, 9 -> 9
			// srcs: (29, 8)(635) 18, (439) 18 --> (636) 36:PENB, ALU, +, NI1
			8'd9 : rdata = 44'b00001110111111100011111111110100000000000000;
			// PEs: 9, 8 -> 9
			// srcs: (30, 9)(686) 54, (492) 0 --> (687) 54:NI0, PENB, +, NI2
			8'd10 : rdata = 44'b00001101000000001101111111011000000000000000;
			// PEs: 11, 8 -> 9
			// srcs: (31, 10)(690) 23, (495) 4 --> (691) 27:PEGB3, PENB, +, NI0
			8'd11 : rdata = 44'b00001111000001101101111111010000000000000000;
			// PEs: 13, 8 -> 10
			// srcs: (32, 11)(692) 18, (498) 40 --> (693) 58:PEGB5, PENB, +, PENB
			8'd12 : rdata = 44'b00001111000010101101111111000000000100000000;
			// PEs: 8, 14 -> 8
			// srcs: (33, 13)(734) 55, (539) 63 --> (735) 118:PENB, PEGB6, +, PEGB0
			8'd13 : rdata = 44'b00001110111111101110000110000000000010000000;
			// PEs: 9 -> 10
			// srcs: (39, 16)(691) 27 --> (691) 27:NI0, pass, PENB
			8'd14 : rdata = 44'b11000101000000000000000000000000000100000000;
			// PEs: 9, 8 -> 9
			// srcs: (49, 14)(636) 36, (638) 30 --> (639) 66:NI1, PENB, +, NI0
			8'd15 : rdata = 44'b00001101000000011101111111010000000000000000;
			// PEs: 8, 9 -> 9
			// srcs: (50, 15)(685) 58, (687) 54 --> (688) 112:PENB, NI2, +, NI1
			8'd16 : rdata = 44'b00001110111111101010000001010100000000000000;
			// PEs: 8, 9 -> 8
			// srcs: (72, 17)(634) 183, (639) 66 --> (640) 249:PENB, NI0, +, PEGB0
			8'd17 : rdata = 44'b00001110111111101010000000000000000010000000;
			// PEs: 8, 9 -> 8
			// srcs: (73, 18)(683) 297, (688) 112 --> (689) 409:PENB, NI1, +, PEGB0
			8'd18 : rdata = 44'b00001110111111101010000000100000000010000000;
			// PEs: 8 -> 
			// srcs: (84, 19)(627) 316 --> (627) 316:PENB, pass, 
			8'd19 : rdata = 44'b11000110111111100000000000000000000000000000;
			// PEs: 8, 9 -> 8
			// srcs: (91, 20)(616) 207, (627) 316 --> (628) 523:PENB, ALU, +, PEGB0
			8'd20 : rdata = 44'b00001110111111100011111111100000000010000000;
			// PEs: 8, 9 -> 10
			// srcs: (181, 21)(805) -9, (12) 1 --> (814) -9:PENB, ND0, *, PENB
			8'd21 : rdata = 44'b00011110111111100110000000000000000100000000;
			// PEs: 9, 10 -> 9
			// srcs: (190, 25)(213) 8, (1014) -9 --> (1214) 17:NW0, PEGB2, -, NW0
			8'd22 : rdata = 44'b00010010000000001110000010000010000000000000;
			// PEs: 8, 9 -> 10
			// srcs: (259, 22)(805) -9, (90) 2 --> (892) -18:PENB, ND1, *, PENB
			8'd23 : rdata = 44'b00011110111111100110000000100000000100000000;
			// PEs: 9, 10 -> 9
			// srcs: (268, 26)(291) 9, (1092) -18 --> (1292) 27:NW1, PEGB2, -, NW1
			8'd24 : rdata = 44'b00010010000000011110000010000010010000000000;
			// PEs: 8, 9 -> 10
			// srcs: (288, 23)(805) -9, (119) 7 --> (921) -63:PENB, ND3, *, PENB
			8'd25 : rdata = 44'b00011110111111100110000001100000000100000000;
			// PEs: 9, 10 -> 9
			// srcs: (297, 27)(320) 1, (1121) -63 --> (1321) 64:NW3, PEGB2, -, NW3
			8'd26 : rdata = 44'b00010010000000111110000010000010110000000000;
			// PEs: 8, 9 -> 10
			// srcs: (337, 24)(805) -9, (168) 2 --> (970) -18:PENB, ND2, *, PENB
			8'd27 : rdata = 44'b00011110111111100110000001000000000100000000;
			// PEs: 9, 10 -> 9
			// srcs: (346, 28)(369) 0, (1170) -18 --> (1370) 18:NW2, PEGB2, -, NW2
			8'd28 : rdata = 44'b00010010000000101110000010000010100000000000;
			default : rdata = 44'b00000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 10) begin
	always @(*) begin
		case(address)
			// PEs: 10, 10 -> 10
			// srcs: (1, 0)(14) 6, (215) 4 --> (415) 24:ND0, NW0, *, NI0
			8'd0 : rdata = 44'b00011011000000000100000000010000000000000000;
			// PEs: 10, 10 -> 11
			// srcs: (2, 1)(92) 7, (293) 1 --> (493) 7:ND1, NW1, *, PENB
			8'd1 : rdata = 44'b00011011000000010100000000100000000100000000;
			// PEs: 10, 10 -> 14
			// srcs: (3, 2)(170) 8, (371) 4 --> (571) 32:ND2, NW2, *, PEGB6
			8'd2 : rdata = 44'b00011011000000100100000001000000000011100000;
			// PEs: 10, 10 -> 10
			// srcs: (4, 3)(122) 3, (323) 6 --> (523) 18:ND3, NW3, *, NI1
			8'd3 : rdata = 44'b00011011000000110100000001110100000000000000;
			// PEs: 10, 11 -> 8
			// srcs: (7, 4)(415) 24, (416) 36 --> (613) 60:NI0, PEGB3, +, PEGB0
			8'd4 : rdata = 44'b00001101000000001110000011000000000010000000;
			// PEs: 10 -> 8
			// srcs: (18, 5)(523) 18 --> (523) 18:NI1, pass, PEGB0
			8'd5 : rdata = 44'b11000101000000010000000000000000000010000000;
			// PEs: 9 -> 
			// srcs: (34, 6)(693) 58 --> (693) 58:PENB, pass, 
			8'd6 : rdata = 44'b11000110111111100000000000000000000000000000;
			// PEs: 9, 10 -> 8
			// srcs: (41, 7)(691) 27, (693) 58 --> (694) 85:PENB, ALU, +, PEGB0
			8'd7 : rdata = 44'b00001110111111100011111111100000000010000000;
			// PEs: 10, 9 -> 9
			// srcs: (184, 12)(3) 1, (814) -9 --> (1014) -9:NM0, PENB, *, PEGB1
			8'd8 : rdata = 44'b00011100000000001101111111000000000010010000;
			// PEs: 8, 10 -> 11
			// srcs: (186, 8)(805) -9, (14) 6 --> (816) -54:PEGB0, ND0, *, PENB
			8'd9 : rdata = 44'b00011111000000000110000000000000000100000000;
			// PEs: 10, 11 -> 10
			// srcs: (195, 17)(215) 4, (1016) -54 --> (1216) 58:NW0, PEGB3, -, NW0
			8'd10 : rdata = 44'b00010010000000001110000011000010000000000000;
			// PEs: 10, 9 -> 9
			// srcs: (262, 13)(3) 1, (892) -18 --> (1092) -18:NM0, PENB, *, PEGB1
			8'd11 : rdata = 44'b00011100000000001101111111000000000010010000;
			// PEs: 8, 10 -> 11
			// srcs: (264, 9)(805) -9, (92) 7 --> (894) -63:PEGB0, ND1, *, PENB
			8'd12 : rdata = 44'b00011111000000000110000000100000000100000000;
			// PEs: 10, 11 -> 10
			// srcs: (273, 18)(293) 1, (1094) -63 --> (1294) 64:NW1, PEGB3, -, NW1
			8'd13 : rdata = 44'b00010010000000011110000011000010010000000000;
			// PEs: 10, 9 -> 9
			// srcs: (291, 14)(3) 1, (921) -63 --> (1121) -63:NM0, PENB, *, PEGB1
			8'd14 : rdata = 44'b00011100000000001101111111000000000010010000;
			// PEs: 8, 10 -> 
			// srcs: (294, 10)(805) -9, (122) 3 --> (924) -27:PEGB0, ND3, *, 
			8'd15 : rdata = 44'b00011111000000000110000001100000000000000000;
			// PEs: 10, 10 -> 
			// srcs: (297, 15)(3) 1, (924) -27 --> (1124) -27:NM0, ALU, *, 
			8'd16 : rdata = 44'b00011100000000000011111111100000000000000000;
			// PEs: 10, 10 -> 10
			// srcs: (300, 19)(323) 6, (1124) -27 --> (1324) 33:NW3, ALU, -, NW3
			8'd17 : rdata = 44'b00010010000000110011111111100010110000000000;
			// PEs: 10, 9 -> 9
			// srcs: (340, 16)(3) 1, (970) -18 --> (1170) -18:NM0, PENB, *, PEGB1
			8'd18 : rdata = 44'b00011100000000001101111111000000000010010000;
			// PEs: 8, 10 -> 11
			// srcs: (342, 11)(805) -9, (170) 8 --> (972) -72:PEGB0, ND2, *, PENB
			8'd19 : rdata = 44'b00011111000000000110000001000000000100000000;
			// PEs: 10, 11 -> 10
			// srcs: (351, 20)(371) 4, (1172) -72 --> (1372) 76:NW2, PEGB3, -, NW2
			8'd20 : rdata = 44'b00010010000000101110000011000010100000000000;
			default : rdata = 44'b00000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 11) begin
	always @(*) begin
		case(address)
			// PEs: 11, 11 -> 10
			// srcs: (1, 0)(15) 4, (216) 9 --> (416) 36:ND0, NW0, *, PEGB2
			8'd0 : rdata = 44'b00011011000000000100000000000000000010100000;
			// PEs: 11, 11 -> 11
			// srcs: (2, 1)(93) 4, (294) 4 --> (494) 16:ND1, NW1, *, NI0
			8'd1 : rdata = 44'b00011011000000010100000000110000000000000000;
			// PEs: 11, 11 -> 14
			// srcs: (3, 2)(171) 7, (372) 5 --> (572) 35:ND2, NW2, *, PEGB6
			8'd2 : rdata = 44'b00011011000000100100000001000000000011100000;
			// PEs: 11, 11 -> 8
			// srcs: (4, 3)(125) 8, (326) 0 --> (526) 0:ND3, NW3, *, PEGB0
			8'd3 : rdata = 44'b00011011000000110100000001100000000010000000;
			// PEs: 10, 11 -> 9
			// srcs: (5, 6)(493) 7, (494) 16 --> (690) 23:PENB, NI0, +, PEGB1
			8'd4 : rdata = 44'b00001110111111101010000000000000000010010000;
			// PEs: 13 -> 
			// srcs: (6, 4)(419) 72 --> (419) 72:PEGB5, pass, 
			8'd5 : rdata = 44'b11000111000010100000000000000000000000000000;
			// PEs: 12, 11 -> 8
			// srcs: (9, 5)(418) 40, (419) 72 --> (617) 112:PEGB4, ALU, +, PEGB0
			8'd6 : rdata = 44'b00001111000010000011111111100000000010000000;
			// PEs: 8, 11 -> 12
			// srcs: (187, 7)(805) -9, (15) 4 --> (817) -36:PEGB0, ND0, *, PENB
			8'd7 : rdata = 44'b00011111000000000110000000000000000100000000;
			// PEs: 11, 10 -> 10
			// srcs: (189, 11)(3) 1, (816) -54 --> (1016) -54:NM0, PENB, *, PEGB2
			8'd8 : rdata = 44'b00011100000000001101111111000000000010100000;
			// PEs: 11, 12 -> 11
			// srcs: (196, 15)(216) 9, (1017) -36 --> (1217) 45:NW0, PEGB4, -, NW0
			8'd9 : rdata = 44'b00010010000000001110000100000010000000000000;
			// PEs: 8, 11 -> 12
			// srcs: (265, 8)(805) -9, (93) 4 --> (895) -36:PEGB0, ND1, *, PENB
			8'd10 : rdata = 44'b00011111000000000110000000100000000100000000;
			// PEs: 11, 10 -> 10
			// srcs: (267, 12)(3) 1, (894) -63 --> (1094) -63:NM0, PENB, *, PEGB2
			8'd11 : rdata = 44'b00011100000000001101111111000000000010100000;
			// PEs: 11, 12 -> 11
			// srcs: (274, 16)(294) 4, (1095) -36 --> (1295) 40:NW1, PEGB4, -, NW1
			8'd12 : rdata = 44'b00010010000000011110000100000010010000000000;
			// PEs: 8, 11 -> 
			// srcs: (297, 9)(805) -9, (125) 8 --> (927) -72:PEGB0, ND3, *, 
			8'd13 : rdata = 44'b00011111000000000110000001100000000000000000;
			// PEs: 11, 11 -> 
			// srcs: (300, 13)(3) 1, (927) -72 --> (1127) -72:NM0, ALU, *, 
			8'd14 : rdata = 44'b00011100000000000011111111100000000000000000;
			// PEs: 11, 11 -> 11
			// srcs: (303, 17)(326) 0, (1127) -72 --> (1327) 72:NW3, ALU, -, NW3
			8'd15 : rdata = 44'b00010010000000110011111111100010110000000000;
			// PEs: 8, 11 -> 12
			// srcs: (343, 10)(805) -9, (171) 7 --> (973) -63:PEGB0, ND2, *, PENB
			8'd16 : rdata = 44'b00011111000000000110000001000000000100000000;
			// PEs: 11, 10 -> 10
			// srcs: (345, 14)(3) 1, (972) -72 --> (1172) -72:NM0, PENB, *, PEGB2
			8'd17 : rdata = 44'b00011100000000001101111111000000000010100000;
			// PEs: 11, 12 -> 11
			// srcs: (352, 18)(372) 5, (1173) -63 --> (1373) 68:NW2, PEGB4, -, NW2
			8'd18 : rdata = 44'b00010010000000101110000100000010100000000000;
			default : rdata = 44'b00000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 12) begin
	always @(*) begin
		case(address)
			// PEs: 12, 12 -> 11
			// srcs: (1, 0)(17) 8, (218) 5 --> (418) 40:ND0, NW0, *, PEGB3
			8'd0 : rdata = 44'b00011011000000000100000000000000000010110000;
			// PEs: 12, 12 -> 13
			// srcs: (2, 1)(95) 8, (296) 0 --> (496) 0:ND1, NW1, *, PENB
			8'd1 : rdata = 44'b00011011000000010100000000100000000100000000;
			// PEs: 12, 12 -> 13
			// srcs: (3, 2)(173) 3, (374) 8 --> (574) 24:ND2, NW2, *, PENB
			8'd2 : rdata = 44'b00011011000000100100000001000000000100000000;
			// PEs: 12, 12 -> 12
			// srcs: (4, 3)(128) 5, (329) 1 --> (529) 5:ND3, NW3, *, NI0
			8'd3 : rdata = 44'b00011011000000110100000001110000000000000000;
			// PEs: 15 -> 
			// srcs: (6, 4)(422) 63 --> (422) 63:PEGB7, pass, 
			8'd4 : rdata = 44'b11000111000011100000000000000000000000000000;
			// PEs: 14, 12 -> 8
			// srcs: (9, 5)(421) 28, (422) 63 --> (619) 91:PEGB6, ALU, +, PEGB0
			8'd5 : rdata = 44'b00001111000011000011111111100000000010000000;
			// PEs: 12 -> 8
			// srcs: (27, 6)(529) 5 --> (529) 5:NI0, pass, PEGB0
			8'd6 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 8, 12 -> 13
			// srcs: (189, 7)(805) -9, (17) 8 --> (819) -72:PEGB0, ND0, *, PENB
			8'd7 : rdata = 44'b00011111000000000110000000000000000100000000;
			// PEs: 12, 11 -> 11
			// srcs: (190, 11)(3) 1, (817) -36 --> (1017) -36:NM0, PENB, *, PEGB3
			8'd8 : rdata = 44'b00011100000000001101111111000000000010110000;
			// PEs: 12, 13 -> 12
			// srcs: (198, 15)(218) 5, (1019) -72 --> (1219) 77:NW0, PEGB5, -, NW0
			8'd9 : rdata = 44'b00010010000000001110000101000010000000000000;
			// PEs: 8, 12 -> 13
			// srcs: (267, 8)(805) -9, (95) 8 --> (897) -72:PEGB0, ND1, *, PENB
			8'd10 : rdata = 44'b00011111000000000110000000100000000100000000;
			// PEs: 12, 11 -> 11
			// srcs: (268, 12)(3) 1, (895) -36 --> (1095) -36:NM0, PENB, *, PEGB3
			8'd11 : rdata = 44'b00011100000000001101111111000000000010110000;
			// PEs: 12, 13 -> 12
			// srcs: (276, 16)(296) 0, (1097) -72 --> (1297) 72:NW1, PEGB5, -, NW1
			8'd12 : rdata = 44'b00010010000000011110000101000010010000000000;
			// PEs: 8, 12 -> 
			// srcs: (300, 9)(805) -9, (128) 5 --> (930) -45:PEGB0, ND3, *, 
			8'd13 : rdata = 44'b00011111000000000110000001100000000000000000;
			// PEs: 12, 12 -> 
			// srcs: (303, 13)(3) 1, (930) -45 --> (1130) -45:NM0, ALU, *, 
			8'd14 : rdata = 44'b00011100000000000011111111100000000000000000;
			// PEs: 12, 12 -> 12
			// srcs: (306, 17)(329) 1, (1130) -45 --> (1330) 46:NW3, ALU, -, NW3
			8'd15 : rdata = 44'b00010010000000110011111111100010110000000000;
			// PEs: 8, 12 -> 13
			// srcs: (345, 10)(805) -9, (173) 3 --> (975) -27:PEGB0, ND2, *, PENB
			8'd16 : rdata = 44'b00011111000000000110000001000000000100000000;
			// PEs: 12, 11 -> 11
			// srcs: (346, 14)(3) 1, (973) -63 --> (1173) -63:NM0, PENB, *, PEGB3
			8'd17 : rdata = 44'b00011100000000001101111111000000000010110000;
			// PEs: 12, 13 -> 12
			// srcs: (354, 18)(374) 8, (1175) -27 --> (1375) 35:NW2, PEGB5, -, NW2
			8'd18 : rdata = 44'b00010010000000101110000101000010100000000000;
			default : rdata = 44'b00000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 13) begin
	always @(*) begin
		case(address)
			// PEs: 13, 13 -> 11
			// srcs: (1, 0)(18) 9, (219) 8 --> (419) 72:ND0, NW0, *, PEGB3
			8'd0 : rdata = 44'b00011011000000000100000000000000000010110000;
			// PEs: 13, 13 -> 13
			// srcs: (2, 1)(96) 9, (297) 2 --> (497) 18:ND1, NW1, *, NI0
			8'd1 : rdata = 44'b00011011000000010100000000110000000000000000;
			// PEs: 13, 13 -> 13
			// srcs: (3, 2)(174) 9, (375) 6 --> (575) 54:ND2, NW2, *, NI1
			8'd2 : rdata = 44'b00011011000000100100000001010100000000000000;
			// PEs: 13, 13 -> 8
			// srcs: (4, 3)(135) 9, (336) 1 --> (536) 9:ND3, NW3, *, PEGB0
			8'd3 : rdata = 44'b00011011000000110100000001100000000010000000;
			// PEs: 12, 13 -> 9
			// srcs: (5, 4)(496) 0, (497) 18 --> (692) 18:PENB, NI0, +, PEGB1
			8'd4 : rdata = 44'b00001110111111101010000000000000000010010000;
			// PEs: 12, 13 -> 8
			// srcs: (6, 5)(574) 24, (575) 54 --> (770) 78:PENB, NI1, +, PEGB0
			8'd5 : rdata = 44'b00001110111111101010000000100000000010000000;
			// PEs: 8, 13 -> 14
			// srcs: (190, 6)(805) -9, (18) 9 --> (820) -81:PEGB0, ND0, *, PENB
			8'd6 : rdata = 44'b00011111000000000110000000000000000100000000;
			// PEs: 13, 12 -> 12
			// srcs: (192, 10)(3) 1, (819) -72 --> (1019) -72:NM0, PENB, *, PEGB4
			8'd7 : rdata = 44'b00011100000000001101111111000000000011000000;
			// PEs: 13, 14 -> 13
			// srcs: (199, 15)(219) 8, (1020) -81 --> (1220) 89:NW0, PEGB6, -, NW0
			8'd8 : rdata = 44'b00010010000000001110000110000010000000000000;
			// PEs: 8, 13 -> 13
			// srcs: (268, 7)(805) -9, (96) 9 --> (898) -81:PEGB0, ND1, *, NI0
			8'd9 : rdata = 44'b00011111000000000110000000110000000000000000;
			// PEs: 13, 12 -> 12
			// srcs: (270, 11)(3) 1, (897) -72 --> (1097) -72:NM0, PENB, *, PEGB4
			8'd10 : rdata = 44'b00011100000000001101111111000000000011000000;
			// PEs: 13, 13 -> 
			// srcs: (271, 12)(3) 1, (898) -81 --> (1098) -81:NM0, NI0, *, 
			8'd11 : rdata = 44'b00011100000000001010000000000000000000000000;
			// PEs: 13, 13 -> 13
			// srcs: (274, 16)(297) 2, (1098) -81 --> (1298) 83:NW1, ALU, -, NW1
			8'd12 : rdata = 44'b00010010000000010011111111100010010000000000;
			// PEs: 8, 13 -> 
			// srcs: (307, 8)(805) -9, (135) 9 --> (937) -81:PEGB0, ND3, *, 
			8'd13 : rdata = 44'b00011111000000000110000001100000000000000000;
			// PEs: 13, 13 -> 
			// srcs: (310, 13)(3) 1, (937) -81 --> (1137) -81:NM0, ALU, *, 
			8'd14 : rdata = 44'b00011100000000000011111111100000000000000000;
			// PEs: 13, 13 -> 13
			// srcs: (313, 17)(336) 1, (1137) -81 --> (1337) 82:NW3, ALU, -, NW3
			8'd15 : rdata = 44'b00010010000000110011111111100010110000000000;
			// PEs: 8, 13 -> 14
			// srcs: (346, 9)(805) -9, (174) 9 --> (976) -81:PEGB0, ND2, *, PENB
			8'd16 : rdata = 44'b00011111000000000110000001000000000100000000;
			// PEs: 13, 12 -> 12
			// srcs: (348, 14)(3) 1, (975) -27 --> (1175) -27:NM0, PENB, *, PEGB4
			8'd17 : rdata = 44'b00011100000000001101111111000000000011000000;
			// PEs: 13, 14 -> 13
			// srcs: (355, 18)(375) 6, (1176) -81 --> (1376) 87:NW2, PEGB6, -, NW2
			8'd18 : rdata = 44'b00010010000000101110000110000010100000000000;
			default : rdata = 44'b00000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 14) begin
	always @(*) begin
		case(address)
			// PEs: 14, 14 -> 12
			// srcs: (1, 0)(20) 7, (221) 4 --> (421) 28:ND0, NW0, *, PEGB4
			8'd0 : rdata = 44'b00011011000000000100000000000000000011000000;
			// PEs: 14, 14 -> 15
			// srcs: (2, 1)(98) 1, (299) 2 --> (499) 2:ND1, NW1, *, PENB
			8'd1 : rdata = 44'b00011011000000010100000000100000000100000000;
			// PEs: 14, 14 -> 15
			// srcs: (3, 2)(176) 6, (377) 8 --> (577) 48:ND2, NW2, *, PENB
			8'd2 : rdata = 44'b00011011000000100100000001000000000100000000;
			// PEs: 14, 14 -> 9
			// srcs: (4, 3)(138) 7, (339) 9 --> (539) 63:ND3, NW3, *, PEGB1
			8'd3 : rdata = 44'b00011011000000110100000001100000000010010000;
			// PEs: 11 -> 
			// srcs: (8, 4)(572) 35 --> (572) 35:PEGB3, pass, 
			8'd4 : rdata = 44'b11000111000001100000000000000000000000000000;
			// PEs: 10, 14 -> 8
			// srcs: (11, 5)(571) 32, (572) 35 --> (767) 67:PEGB2, ALU, +, PEGB0
			8'd5 : rdata = 44'b00001111000001000011111111100000000010000000;
			// PEs: 8, 14 -> 14
			// srcs: (192, 6)(805) -9, (20) 7 --> (822) -63:PEGB0, ND0, *, NI0
			8'd6 : rdata = 44'b00011111000000000110000000010000000000000000;
			// PEs: 14, 13 -> 13
			// srcs: (193, 10)(3) 1, (820) -81 --> (1020) -81:NM0, PENB, *, PEGB5
			8'd7 : rdata = 44'b00011100000000001101111111000000000011010000;
			// PEs: 14, 14 -> 
			// srcs: (195, 11)(3) 1, (822) -63 --> (1022) -63:NM0, NI0, *, 
			8'd8 : rdata = 44'b00011100000000001010000000000000000000000000;
			// PEs: 14, 14 -> 14
			// srcs: (198, 16)(221) 4, (1022) -63 --> (1222) 67:NW0, ALU, -, NW0
			8'd9 : rdata = 44'b00010010000000000011111111100010000000000000;
			// PEs: 8, 14 -> 
			// srcs: (270, 7)(805) -9, (98) 1 --> (900) -9:PEGB0, ND1, *, 
			8'd10 : rdata = 44'b00011111000000000110000000100000000000000000;
			// PEs: 14, 14 -> 
			// srcs: (273, 12)(3) 1, (900) -9 --> (1100) -9:NM0, ALU, *, 
			8'd11 : rdata = 44'b00011100000000000011111111100000000000000000;
			// PEs: 14, 14 -> 14
			// srcs: (276, 17)(299) 2, (1100) -9 --> (1300) 11:NW1, ALU, -, NW1
			8'd12 : rdata = 44'b00010010000000010011111111100010010000000000;
			// PEs: 8, 14 -> 
			// srcs: (310, 8)(805) -9, (138) 7 --> (940) -63:PEGB0, ND3, *, 
			8'd13 : rdata = 44'b00011111000000000110000001100000000000000000;
			// PEs: 14, 14 -> 
			// srcs: (313, 13)(3) 1, (940) -63 --> (1140) -63:NM0, ALU, *, 
			8'd14 : rdata = 44'b00011100000000000011111111100000000000000000;
			// PEs: 14, 14 -> 14
			// srcs: (316, 18)(339) 9, (1140) -63 --> (1340) 72:NW3, ALU, -, NW3
			8'd15 : rdata = 44'b00010010000000110011111111100010110000000000;
			// PEs: 8, 14 -> 14
			// srcs: (348, 9)(805) -9, (176) 6 --> (978) -54:PEGB0, ND2, *, NI0
			8'd16 : rdata = 44'b00011111000000000110000001010000000000000000;
			// PEs: 14, 13 -> 13
			// srcs: (349, 14)(3) 1, (976) -81 --> (1176) -81:NM0, PENB, *, PEGB5
			8'd17 : rdata = 44'b00011100000000001101111111000000000011010000;
			// PEs: 14, 14 -> 
			// srcs: (351, 15)(3) 1, (978) -54 --> (1178) -54:NM0, NI0, *, 
			8'd18 : rdata = 44'b00011100000000001010000000000000000000000000;
			// PEs: 14, 14 -> 14
			// srcs: (354, 19)(377) 8, (1178) -54 --> (1378) 62:NW2, ALU, -, NW2
			8'd19 : rdata = 44'b00010010000000100011111111100010100000000000;
			default : rdata = 44'b00000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 15) begin
	always @(*) begin
		case(address)
			// PEs: 15, 15 -> 12
			// srcs: (1, 0)(21) 9, (222) 7 --> (422) 63:ND0, NW0, *, PEGB4
			8'd0 : rdata = 44'b00011011000000000100000000000000000011000000;
			// PEs: 15, 15 -> 15
			// srcs: (2, 1)(99) 9, (300) 7 --> (500) 63:ND1, NW1, *, NI0
			8'd1 : rdata = 44'b00011011000000010100000000110000000000000000;
			// PEs: 15, 15 -> 15
			// srcs: (3, 2)(177) 0, (378) 1 --> (578) 0:ND2, NW2, *, NI1
			8'd2 : rdata = 44'b00011011000000100100000001010100000000000000;
			// PEs: 15, 15 -> 15
			// srcs: (4, 3)(141) 9, (342) 8 --> (542) 72:ND3, NW3, *, NI2
			8'd3 : rdata = 44'b00011011000000110100000001111000000000000000;
			// PEs: 14, 15 -> 8
			// srcs: (5, 4)(499) 2, (500) 63 --> (695) 65:PENB, NI0, +, PENB
			8'd4 : rdata = 44'b00001110111111101010000000000000000100000000;
			// PEs: 14, 15 -> 15
			// srcs: (6, 5)(577) 48, (578) 0 --> (772) 48:PENB, NI1, +, NI0
			8'd5 : rdata = 44'b00001110111111101010000000110000000000000000;
			// PEs: 15 -> 8
			// srcs: (12, 6)(542) 72 --> (542) 72:NI2, pass, PENB
			8'd6 : rdata = 44'b11000101000000100000000000000000000100000000;
			// PEs: 15 -> 8
			// srcs: (24, 7)(772) 48 --> (772) 48:NI0, pass, PENB
			8'd7 : rdata = 44'b11000101000000000000000000000000000100000000;
			// PEs: 8, 15 -> 
			// srcs: (193, 8)(805) -9, (21) 9 --> (823) -81:PEGB0, ND0, *, 
			8'd8 : rdata = 44'b00011111000000000110000000000000000000000000;
			// PEs: 15, 15 -> 
			// srcs: (196, 12)(3) 1, (823) -81 --> (1023) -81:NM0, ALU, *, 
			8'd9 : rdata = 44'b00011100000000000011111111100000000000000000;
			// PEs: 15, 15 -> 15
			// srcs: (199, 16)(222) 7, (1023) -81 --> (1223) 88:NW0, ALU, -, NW0
			8'd10 : rdata = 44'b00010010000000000011111111100010000000000000;
			// PEs: 8, 15 -> 
			// srcs: (271, 9)(805) -9, (99) 9 --> (901) -81:PEGB0, ND1, *, 
			8'd11 : rdata = 44'b00011111000000000110000000100000000000000000;
			// PEs: 15, 15 -> 
			// srcs: (274, 13)(3) 1, (901) -81 --> (1101) -81:NM0, ALU, *, 
			8'd12 : rdata = 44'b00011100000000000011111111100000000000000000;
			// PEs: 15, 15 -> 15
			// srcs: (277, 17)(300) 7, (1101) -81 --> (1301) 88:NW1, ALU, -, NW1
			8'd13 : rdata = 44'b00010010000000010011111111100010010000000000;
			// PEs: 8, 15 -> 
			// srcs: (313, 10)(805) -9, (141) 9 --> (943) -81:PEGB0, ND3, *, 
			8'd14 : rdata = 44'b00011111000000000110000001100000000000000000;
			// PEs: 15, 15 -> 
			// srcs: (316, 14)(3) 1, (943) -81 --> (1143) -81:NM0, ALU, *, 
			8'd15 : rdata = 44'b00011100000000000011111111100000000000000000;
			// PEs: 15, 15 -> 15
			// srcs: (319, 18)(342) 8, (1143) -81 --> (1343) 89:NW3, ALU, -, NW3
			8'd16 : rdata = 44'b00010010000000110011111111100010110000000000;
			// PEs: 8, 15 -> 
			// srcs: (349, 11)(805) -9, (177) 0 --> (979) 0:PEGB0, ND2, *, 
			8'd17 : rdata = 44'b00011111000000000110000001000000000000000000;
			// PEs: 15, 15 -> 
			// srcs: (352, 15)(3) 1, (979) 0 --> (1179) 0:NM0, ALU, *, 
			8'd18 : rdata = 44'b00011100000000000011111111100000000000000000;
			// PEs: 15, 15 -> 15
			// srcs: (355, 19)(378) 1, (1179) 0 --> (1379) 1:NW2, ALU, -, NW2
			8'd19 : rdata = 44'b00010010000000100011111111100010100000000000;
			default : rdata = 44'b00000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 16) begin
	always @(*) begin
		case(address)
			// PEs: 23 -> 24
			// srcs: (4, 0)(509) 12 --> (509) 12:PENB, pass, PUNB
			8'd0 : rdata = 44'b11000110111111100000000000000000001000000000;
			// PEs: 23 -> 24
			// srcs: (5, 1)(587) 28 --> (587) 28:PENB, pass, PUNB
			8'd1 : rdata = 44'b11000110111111100000000000000000001000000000;
			// PEs: 18 -> 32
			// srcs: (9, 20)(548) 0 --> (548) 0:PEGB2, pass, PUGB4
			8'd2 : rdata = 44'b11000111000001000000000000000000000000001100;
			// PEs: 23 -> 24
			// srcs: (10, 2)(432) 56 --> (432) 56:PENB, pass, PUNB
			8'd3 : rdata = 44'b11000110111111100000000000000000001000000000;
			// PEs: 32 -> 16
			// srcs: (11, 4)(417) 0 --> (417) 0:PUGB4, pass, NI0
			8'd4 : rdata = 44'b11000111000010010000000000010000000000000000;
			// PEs: 17 -> 48
			// srcs: (12, 6)(622) 46 --> (622) 46:PEGB1, pass, PUGB6
			8'd5 : rdata = 44'b11000111000000100000000000000000000000001110;
			// PEs: 18 -> 40
			// srcs: (13, 12)(697) 64 --> (697) 64:PEGB2, pass, PUGB5
			8'd6 : rdata = 44'b11000111000001000000000000000000000000001101;
			// PEs: 8 -> 17
			// srcs: (14, 3)(613) 60 --> (613) 60:PUNB, pass, PENB
			8'd7 : rdata = 44'b11000110111111110000000000000000000100000000;
			// PEs: 18 -> 56
			// srcs: (15, 7)(624) 48 --> (624) 48:PEGB2, pass, PUGB7
			8'd8 : rdata = 44'b11000111000001000000000000000000000000001111;
			// PEs: 19 -> 24
			// srcs: (16, 8)(629) 23 --> (629) 23:PEGB3, pass, PUNB
			8'd9 : rdata = 44'b11000111000001100000000000000000001000000000;
			// PEs: 20 -> 40
			// srcs: (17, 22)(554) 14 --> (554) 14:PEGB4, pass, PUGB5
			8'd10 : rdata = 44'b11000111000010000000000000000000000000001101;
			// PEs: 21 -> 0
			// srcs: (18, 23)(561) 18 --> (561) 18:PEGB5, pass, PUGB0
			8'd11 : rdata = 44'b11000111000010100000000000000000000000001000;
			// PEs: 16 -> 17
			// srcs: (21, 5)(417) 0 --> (417) 0:NI0, pass, PENB
			8'd12 : rdata = 44'b11000101000000000000000000000000000100000000;
			// PEs: 32 -> 16
			// srcs: (22, 9)(641) 51 --> (641) 51:PUGB4, pass, NI0
			8'd13 : rdata = 44'b11000111000010010000000000010000000000000000;
			// PEs: 48 -> 17
			// srcs: (23, 10)(445) 30 --> (445) 30:PUGB6, pass, PENB
			8'd14 : rdata = 44'b11000111000011010000000000000000000100000000;
			// PEs: 17 -> 56
			// srcs: (24, 19)(545) 36 --> (545) 36:PEGB1, pass, PUGB7
			8'd15 : rdata = 44'b11000111000000100000000000000000000000001111;
			// PEs: 19 -> 48
			// srcs: (25, 21)(551) 21 --> (551) 21:PEGB3, pass, PUGB6
			8'd16 : rdata = 44'b11000111000001100000000000000000000000001110;
			// PEs: 22 -> 56
			// srcs: (26, 24)(564) 0 --> (564) 0:PEGB6, pass, PUGB7
			8'd17 : rdata = 44'b11000111000011000000000000000000000000001111;
			// PEs: 23 -> 0
			// srcs: (27, 25)(567) 7 --> (567) 7:PENB, pass, PUGB0
			8'd18 : rdata = 44'b11000110111111100000000000000000000000001000;
			// PEs: 22 -> 24
			// srcs: (28, 26)(780) 56 --> (780) 56:PEGB6, pass, PUNB
			8'd19 : rdata = 44'b11000111000011000000000000000000001000000000;
			// PEs: 16 -> 17
			// srcs: (29, 11)(641) 51 --> (641) 51:NI0, pass, PENB
			8'd20 : rdata = 44'b11000101000000000000000000000000000100000000;
			// PEs: 24 -> 16
			// srcs: (30, 13)(710) 20 --> (710) 20:PUGB3, pass, NI0
			8'd21 : rdata = 44'b11000111000001110000000000010000000000000000;
			// PEs: 0 -> 17
			// srcs: (31, 14)(514) 20 --> (514) 20:PUGB0, pass, PENB
			8'd22 : rdata = 44'b11000111000000010000000000000000000100000000;
			// PEs: 17 -> 40
			// srcs: (32, 27)(614) 60 --> (614) 60:PEGB1, pass, PUGB5
			8'd23 : rdata = 44'b11000111000000100000000000000000000000001101;
			// PEs: 17 -> 0
			// srcs: (36, 28)(642) 81 --> (642) 81:PEGB1, pass, PUGB0
			8'd24 : rdata = 44'b11000111000000100000000000000000000000001000;
			// PEs: 16 -> 17
			// srcs: (37, 15)(710) 20 --> (710) 20:NI0, pass, PENB
			8'd25 : rdata = 44'b11000101000000000000000000000000000100000000;
			// PEs: 24 -> 16
			// srcs: (38, 16)(716) 46 --> (716) 46:PUGB3, pass, NI0
			8'd26 : rdata = 44'b11000111000001110000000000010000000000000000;
			// PEs: 8 -> 17
			// srcs: (39, 17)(520) 7 --> (520) 7:PUNB, pass, PENB
			8'd27 : rdata = 44'b11000110111111110000000000000000000100000000;
			// PEs: 23 -> 56
			// srcs: (40, 32)(706) 11 --> (706) 11:PENB, pass, PUGB7
			8'd28 : rdata = 44'b11000110111111100000000000000000000000001111;
			// PEs: 17 -> 24
			// srcs: (44, 33)(711) 40 --> (711) 40:PEGB1, pass, PUNB
			8'd29 : rdata = 44'b11000111000000100000000000000000001000000000;
			// PEs: 16 -> 17
			// srcs: (45, 18)(716) 46 --> (716) 46:NI0, pass, PENB
			8'd30 : rdata = 44'b11000101000000000000000000000000000100000000;
			// PEs: 0 -> 16
			// srcs: (46, 29)(696) 77 --> (696) 77:PUGB0, pass, NI0
			8'd31 : rdata = 44'b11000111000000010000000000010000000000000000;
			// PEs: 21 -> 24
			// srcs: (47, 38)(779) 42 --> (779) 42:PEGB5, pass, PUNB
			8'd32 : rdata = 44'b11000111000010100000000000000000001000000000;
			// PEs: 40 -> 17
			// srcs: (48, 30)(698) 69 --> (698) 69:PUGB5, pass, PENB
			8'd33 : rdata = 44'b11000111000010110000000000000000000100000000;
			// PEs: 17 -> 40
			// srcs: (52, 34)(717) 53 --> (717) 53:PEGB1, pass, PUGB5
			8'd34 : rdata = 44'b11000111000000100000000000000000000000001101;
			// PEs: 16 -> 17
			// srcs: (55, 31)(696) 77 --> (696) 77:NI0, pass, PENB
			8'd35 : rdata = 44'b11000101000000000000000000000000000100000000;
			// PEs: 8 -> 16
			// srcs: (56, 35)(735) 118 --> (735) 118:PUNB, pass, NI0
			8'd36 : rdata = 44'b11000110111111110000000000010000000000000000;
			// PEs: 48 -> 17
			// srcs: (57, 36)(737) 149 --> (737) 149:PUGB6, pass, PENB
			8'd37 : rdata = 44'b11000111000011010000000000000000000100000000;
			// PEs: 16 -> 17
			// srcs: (63, 37)(735) 118 --> (735) 118:NI0, pass, PENB
			8'd38 : rdata = 44'b11000101000000000000000000000000000100000000;
			// PEs: 8 -> 17
			// srcs: (64, 39)(694) 85 --> (694) 85:PUNB, pass, PENB
			8'd39 : rdata = 44'b11000110111111110000000000000000000100000000;
			// PEs: 17 -> 48
			// srcs: (70, 40)(738) 267 --> (738) 267:PEGB1, pass, PUGB6
			8'd40 : rdata = 44'b11000111000000100000000000000000000000001110;
			// PEs: 8 -> 16
			// srcs: (80, 41)(640) 249 --> (640) 249:PUNB, pass, NI0
			8'd41 : rdata = 44'b11000110111111110000000000010000000000000000;
			// PEs: 48 -> 17
			// srcs: (83, 42)(651) 315 --> (651) 315:PUGB6, pass, PENB
			8'd42 : rdata = 44'b11000111000011010000000000000000000100000000;
			// PEs: 16 -> 17
			// srcs: (90, 43)(640) 249 --> (640) 249:NI0, pass, PENB
			8'd43 : rdata = 44'b11000101000000000000000000000000000100000000;
			// PEs: 8 -> 17
			// srcs: (91, 44)(689) 409 --> (689) 409:PUNB, pass, PENB
			8'd44 : rdata = 44'b11000110111111110000000000000000000100000000;
			// PEs: 8 -> 17
			// srcs: (98, 45)(628) 523 --> (628) 523:PUNB, pass, PENB
			8'd45 : rdata = 44'b11000110111111110000000000000000000100000000;
			// PEs: 17 -> 24
			// srcs: (99, 46)(701) 640 --> (701) 640:PEGB1, pass, PUNB
			8'd46 : rdata = 44'b11000111000000100000000000000000001000000000;
			// PEs: 17 -> 24
			// srcs: (107, 47)(653) 1087 --> (653) 1087:PEGB1, pass, PUNB
			8'd47 : rdata = 44'b11000111000000100000000000000000001000000000;
			// PEs: 0 -> 17
			// srcs: (193, 48)(805) -9 --> (805) -9:PUGB0, pass, PENB
			8'd48 : rdata = 44'b11000111000000010000000000000000000100000000;
			// PEs: 0 -> 18
			// srcs: (194, 49)(805) -9 --> (805) -9:PUGB0, pass, PEGB2
			8'd49 : rdata = 44'b11000111000000010000000000000000000010100000;
			// PEs: 0 -> 19
			// srcs: (196, 50)(805) -9 --> (805) -9:PUGB0, pass, PEGB3
			8'd50 : rdata = 44'b11000111000000010000000000000000000010110000;
			// PEs: 0 -> 20
			// srcs: (197, 51)(805) -9 --> (805) -9:PUGB0, pass, PEGB4
			8'd51 : rdata = 44'b11000111000000010000000000000000000011000000;
			// PEs: 0 -> 21
			// srcs: (199, 52)(805) -9 --> (805) -9:PUGB0, pass, PEGB5
			8'd52 : rdata = 44'b11000111000000010000000000000000000011010000;
			// PEs: 0 -> 22
			// srcs: (200, 53)(805) -9 --> (805) -9:PUGB0, pass, PEGB6
			8'd53 : rdata = 44'b11000111000000010000000000000000000011100000;
			// PEs: 0 -> 23
			// srcs: (201, 54)(805) -9 --> (805) -9:PUGB0, pass, PEGB7
			8'd54 : rdata = 44'b11000111000000010000000000000000000011110000;
			// PEs: 0 -> 17
			// srcs: (271, 55)(805) -9 --> (805) -9:PUGB0, pass, PENB
			8'd55 : rdata = 44'b11000111000000010000000000000000000100000000;
			// PEs: 0 -> 18
			// srcs: (272, 56)(805) -9 --> (805) -9:PUGB0, pass, PEGB2
			8'd56 : rdata = 44'b11000111000000010000000000000000000010100000;
			// PEs: 0 -> 19
			// srcs: (274, 57)(805) -9 --> (805) -9:PUGB0, pass, PEGB3
			8'd57 : rdata = 44'b11000111000000010000000000000000000010110000;
			// PEs: 0 -> 20
			// srcs: (275, 58)(805) -9 --> (805) -9:PUGB0, pass, PEGB4
			8'd58 : rdata = 44'b11000111000000010000000000000000000011000000;
			// PEs: 0 -> 21
			// srcs: (276, 59)(805) -9 --> (805) -9:PUGB0, pass, PEGB5
			8'd59 : rdata = 44'b11000111000000010000000000000000000011010000;
			// PEs: 0 -> 22
			// srcs: (277, 60)(805) -9 --> (805) -9:PUGB0, pass, PEGB6
			8'd60 : rdata = 44'b11000111000000010000000000000000000011100000;
			// PEs: 0 -> 23
			// srcs: (278, 61)(805) -9 --> (805) -9:PUGB0, pass, PEGB7
			8'd61 : rdata = 44'b11000111000000010000000000000000000011110000;
			// PEs: 0 -> 17
			// srcs: (314, 62)(805) -9 --> (805) -9:PUGB0, pass, PENB
			8'd62 : rdata = 44'b11000111000000010000000000000000000100000000;
			// PEs: 0 -> 18
			// srcs: (317, 63)(805) -9 --> (805) -9:PUGB0, pass, PEGB2
			8'd63 : rdata = 44'b11000111000000010000000000000000000010100000;
			// PEs: 0 -> 19
			// srcs: (320, 64)(805) -9 --> (805) -9:PUGB0, pass, PEGB3
			8'd64 : rdata = 44'b11000111000000010000000000000000000010110000;
			// PEs: 0 -> 20
			// srcs: (323, 65)(805) -9 --> (805) -9:PUGB0, pass, PEGB4
			8'd65 : rdata = 44'b11000111000000010000000000000000000011000000;
			// PEs: 0 -> 21
			// srcs: (330, 66)(805) -9 --> (805) -9:PUGB0, pass, PEGB5
			8'd66 : rdata = 44'b11000111000000010000000000000000000011010000;
			// PEs: 0 -> 22
			// srcs: (333, 67)(805) -9 --> (805) -9:PUGB0, pass, PEGB6
			8'd67 : rdata = 44'b11000111000000010000000000000000000011100000;
			// PEs: 0 -> 23
			// srcs: (336, 68)(805) -9 --> (805) -9:PUGB0, pass, PEGB7
			8'd68 : rdata = 44'b11000111000000010000000000000000000011110000;
			// PEs: 0 -> 17
			// srcs: (349, 69)(805) -9 --> (805) -9:PUGB0, pass, PENB
			8'd69 : rdata = 44'b11000111000000010000000000000000000100000000;
			// PEs: 0 -> 18
			// srcs: (350, 70)(805) -9 --> (805) -9:PUGB0, pass, PEGB2
			8'd70 : rdata = 44'b11000111000000010000000000000000000010100000;
			// PEs: 0 -> 19
			// srcs: (351, 71)(805) -9 --> (805) -9:PUGB0, pass, PEGB3
			8'd71 : rdata = 44'b11000111000000010000000000000000000010110000;
			// PEs: 0 -> 20
			// srcs: (352, 72)(805) -9 --> (805) -9:PUGB0, pass, PEGB4
			8'd72 : rdata = 44'b11000111000000010000000000000000000011000000;
			// PEs: 0 -> 21
			// srcs: (353, 73)(805) -9 --> (805) -9:PUGB0, pass, PEGB5
			8'd73 : rdata = 44'b11000111000000010000000000000000000011010000;
			// PEs: 0 -> 22
			// srcs: (354, 74)(805) -9 --> (805) -9:PUGB0, pass, PEGB6
			8'd74 : rdata = 44'b11000111000000010000000000000000000011100000;
			// PEs: 0 -> 23
			// srcs: (356, 75)(805) -9 --> (805) -9:PUGB0, pass, PEGB7
			8'd75 : rdata = 44'b11000111000000010000000000000000000011110000;
			default : rdata = 44'b00000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 17) begin
	always @(*) begin
		case(address)
			// PEs: 17, 17 -> 17
			// srcs: (1, 0)(23) 5, (224) 2 --> (424) 10:ND0, NW0, *, NI0
			8'd0 : rdata = 44'b00011011000000000100000000010000000000000000;
			// PEs: 17, 17 -> 18
			// srcs: (2, 1)(101) 8, (302) 8 --> (502) 64:ND1, NW1, *, PENB
			8'd1 : rdata = 44'b00011011000000010100000000100000000100000000;
			// PEs: 17, 17 -> 21
			// srcs: (3, 2)(179) 9, (380) 2 --> (580) 18:ND2, NW2, *, PEGB5
			8'd2 : rdata = 44'b00011011000000100100000001000000000011010000;
			// PEs: 17, 17 -> 17
			// srcs: (4, 3)(144) 4, (345) 9 --> (545) 36:ND3, NW3, *, NI1
			8'd3 : rdata = 44'b00011011000000110100000001110100000000000000;
			// PEs: 17, 18 -> 16
			// srcs: (7, 4)(424) 10, (425) 36 --> (622) 46:NI0, PEGB2, +, PEGB0
			8'd4 : rdata = 44'b00001101000000001110000010000000000010000000;
			// PEs: 16 -> 17
			// srcs: (16, 5)(613) 60 --> (613) 60:PENB, pass, NI0
			8'd5 : rdata = 44'b11000110111111100000000000010000000000000000;
			// PEs: 17 -> 16
			// srcs: (19, 13)(545) 36 --> (545) 36:NI1, pass, PEGB0
			8'd6 : rdata = 44'b11000101000000010000000000000000000010000000;
			// PEs: 17, 16 -> 16
			// srcs: (23, 6)(613) 60, (417) 0 --> (614) 60:NI0, PENB, +, PEGB0
			8'd7 : rdata = 44'b00001101000000001101111111000000000010000000;
			// PEs: 16 -> 
			// srcs: (25, 7)(445) 30 --> (445) 30:PENB, pass, 
			8'd8 : rdata = 44'b11000110111111100000000000000000000000000000;
			// PEs: 16, 17 -> 16
			// srcs: (31, 8)(641) 51, (445) 30 --> (642) 81:PENB, ALU, +, PEGB0
			8'd9 : rdata = 44'b00001110111111100011111111100000000010000000;
			// PEs: 16 -> 
			// srcs: (33, 9)(514) 20 --> (514) 20:PENB, pass, 
			8'd10 : rdata = 44'b11000110111111100000000000000000000000000000;
			// PEs: 16, 17 -> 16
			// srcs: (39, 10)(710) 20, (514) 20 --> (711) 40:PENB, ALU, +, PEGB0
			8'd11 : rdata = 44'b00001110111111100011111111100000000010000000;
			// PEs: 16 -> 
			// srcs: (41, 11)(520) 7 --> (520) 7:PENB, pass, 
			8'd12 : rdata = 44'b11000110111111100000000000000000000000000000;
			// PEs: 16, 17 -> 16
			// srcs: (47, 12)(716) 46, (520) 7 --> (717) 53:PENB, ALU, +, PEGB0
			8'd13 : rdata = 44'b00001110111111100011111111100000000010000000;
			// PEs: 16 -> 
			// srcs: (50, 14)(698) 69 --> (698) 69:PENB, pass, 
			8'd14 : rdata = 44'b11000110111111100000000000000000000000000000;
			// PEs: 16, 17 -> 17
			// srcs: (57, 15)(696) 77, (698) 69 --> (699) 146:PENB, ALU, +, NI0
			8'd15 : rdata = 44'b00001110111111100011111111110000000000000000;
			// PEs: 16 -> 
			// srcs: (59, 16)(737) 149 --> (737) 149:PENB, pass, 
			8'd16 : rdata = 44'b11000110111111100000000000000000000000000000;
			// PEs: 16, 17 -> 16
			// srcs: (65, 17)(735) 118, (737) 149 --> (738) 267:PENB, ALU, +, PEGB0
			8'd17 : rdata = 44'b00001110111111100011111111100000000010000000;
			// PEs: 16, 17 -> 17
			// srcs: (67, 18)(694) 85, (699) 146 --> (700) 231:PENB, NI0, +, NI1
			8'd18 : rdata = 44'b00001110111111101010000000010100000000000000;
			// PEs: 16 -> 
			// srcs: (85, 19)(651) 315 --> (651) 315:PENB, pass, 
			8'd19 : rdata = 44'b11000110111111100000000000000000000000000000;
			// PEs: 16, 17 -> 17
			// srcs: (92, 20)(640) 249, (651) 315 --> (652) 564:PENB, ALU, +, NI0
			8'd20 : rdata = 44'b00001110111111100011111111110000000000000000;
			// PEs: 16, 17 -> 16
			// srcs: (93, 21)(689) 409, (700) 231 --> (701) 640:PENB, NI1, +, PEGB0
			8'd21 : rdata = 44'b00001110111111101010000000100000000010000000;
			// PEs: 16, 17 -> 16
			// srcs: (102, 22)(628) 523, (652) 564 --> (653) 1087:PENB, NI0, +, PEGB0
			8'd22 : rdata = 44'b00001110111111101010000000000000000010000000;
			// PEs: 16, 17 -> 18
			// srcs: (195, 23)(805) -9, (23) 5 --> (825) -45:PENB, ND0, *, PENB
			8'd23 : rdata = 44'b00011110111111100110000000000000000100000000;
			// PEs: 17, 18 -> 17
			// srcs: (204, 27)(224) 2, (1025) -45 --> (1225) 47:NW0, PEGB2, -, NW0
			8'd24 : rdata = 44'b00010010000000001110000010000010000000000000;
			// PEs: 16, 17 -> 18
			// srcs: (273, 24)(805) -9, (101) 8 --> (903) -72:PENB, ND1, *, PENB
			8'd25 : rdata = 44'b00011110111111100110000000100000000100000000;
			// PEs: 17, 18 -> 17
			// srcs: (282, 28)(302) 8, (1103) -72 --> (1303) 80:NW1, PEGB2, -, NW1
			8'd26 : rdata = 44'b00010010000000011110000010000010010000000000;
			// PEs: 16, 17 -> 18
			// srcs: (316, 25)(805) -9, (144) 4 --> (946) -36:PENB, ND3, *, PENB
			8'd27 : rdata = 44'b00011110111111100110000001100000000100000000;
			// PEs: 17, 18 -> 17
			// srcs: (325, 29)(345) 9, (1146) -36 --> (1346) 45:NW3, PEGB2, -, NW3
			8'd28 : rdata = 44'b00010010000000111110000010000010110000000000;
			// PEs: 16, 17 -> 18
			// srcs: (351, 26)(805) -9, (179) 9 --> (981) -81:PENB, ND2, *, PENB
			8'd29 : rdata = 44'b00011110111111100110000001000000000100000000;
			// PEs: 17, 18 -> 17
			// srcs: (360, 30)(380) 2, (1181) -81 --> (1381) 83:NW2, PEGB2, -, NW2
			8'd30 : rdata = 44'b00010010000000101110000010000010100000000000;
			default : rdata = 44'b00000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 18) begin
	always @(*) begin
		case(address)
			// PEs: 18, 18 -> 17
			// srcs: (1, 0)(24) 9, (225) 4 --> (425) 36:ND0, NW0, *, PEGB1
			8'd0 : rdata = 44'b00011011000000000100000000000000000010010000;
			// PEs: 18, 18 -> 18
			// srcs: (2, 1)(102) 5, (303) 0 --> (503) 0:ND1, NW1, *, NI0
			8'd1 : rdata = 44'b00011011000000010100000000110000000000000000;
			// PEs: 18, 18 -> 21
			// srcs: (3, 2)(180) 6, (381) 0 --> (581) 0:ND2, NW2, *, PEGB5
			8'd2 : rdata = 44'b00011011000000100100000001000000000011010000;
			// PEs: 18, 18 -> 16
			// srcs: (4, 3)(147) 6, (348) 0 --> (548) 0:ND3, NW3, *, PEGB0
			8'd3 : rdata = 44'b00011011000000110100000001100000000010000000;
			// PEs: 17, 18 -> 16
			// srcs: (5, 6)(502) 64, (503) 0 --> (697) 64:PENB, NI0, +, PEGB0
			8'd4 : rdata = 44'b00001110111111101010000000000000000010000000;
			// PEs: 20 -> 
			// srcs: (6, 4)(428) 48 --> (428) 48:PEGB4, pass, 
			8'd5 : rdata = 44'b11000111000010000000000000000000000000000000;
			// PEs: 19, 18 -> 16
			// srcs: (9, 5)(427) 0, (428) 48 --> (624) 48:PEGB3, ALU, +, PEGB0
			8'd6 : rdata = 44'b00001111000001100011111111100000000010000000;
			// PEs: 18, 17 -> 17
			// srcs: (198, 11)(3) 1, (825) -45 --> (1025) -45:NM0, PENB, *, PEGB1
			8'd7 : rdata = 44'b00011100000000001101111111000000000010010000;
			// PEs: 16, 18 -> 19
			// srcs: (199, 7)(805) -9, (24) 9 --> (826) -81:PEGB0, ND0, *, PENB
			8'd8 : rdata = 44'b00011111000000000110000000000000000100000000;
			// PEs: 18, 19 -> 18
			// srcs: (208, 16)(225) 4, (1026) -81 --> (1226) 85:NW0, PEGB3, -, NW0
			8'd9 : rdata = 44'b00010010000000001110000011000010000000000000;
			// PEs: 18, 17 -> 17
			// srcs: (276, 12)(3) 1, (903) -72 --> (1103) -72:NM0, PENB, *, PEGB1
			8'd10 : rdata = 44'b00011100000000001101111111000000000010010000;
			// PEs: 16, 18 -> 19
			// srcs: (277, 8)(805) -9, (102) 5 --> (904) -45:PEGB0, ND1, *, PENB
			8'd11 : rdata = 44'b00011111000000000110000000100000000100000000;
			// PEs: 18, 19 -> 18
			// srcs: (286, 17)(303) 0, (1104) -45 --> (1304) 45:NW1, PEGB3, -, NW1
			8'd12 : rdata = 44'b00010010000000011110000011000010010000000000;
			// PEs: 18, 17 -> 17
			// srcs: (319, 13)(3) 1, (946) -36 --> (1146) -36:NM0, PENB, *, PEGB1
			8'd13 : rdata = 44'b00011100000000001101111111000000000010010000;
			// PEs: 16, 18 -> 
			// srcs: (322, 9)(805) -9, (147) 6 --> (949) -54:PEGB0, ND3, *, 
			8'd14 : rdata = 44'b00011111000000000110000001100000000000000000;
			// PEs: 18, 18 -> 
			// srcs: (325, 14)(3) 1, (949) -54 --> (1149) -54:NM0, ALU, *, 
			8'd15 : rdata = 44'b00011100000000000011111111100000000000000000;
			// PEs: 18, 18 -> 18
			// srcs: (328, 18)(348) 0, (1149) -54 --> (1349) 54:NW3, ALU, -, NW3
			8'd16 : rdata = 44'b00010010000000110011111111100010110000000000;
			// PEs: 18, 17 -> 17
			// srcs: (354, 15)(3) 1, (981) -81 --> (1181) -81:NM0, PENB, *, PEGB1
			8'd17 : rdata = 44'b00011100000000001101111111000000000010010000;
			// PEs: 16, 18 -> 19
			// srcs: (355, 10)(805) -9, (180) 6 --> (982) -54:PEGB0, ND2, *, PENB
			8'd18 : rdata = 44'b00011111000000000110000001000000000100000000;
			// PEs: 18, 19 -> 18
			// srcs: (364, 19)(381) 0, (1182) -54 --> (1382) 54:NW2, PEGB3, -, NW2
			8'd19 : rdata = 44'b00010010000000101110000011000010100000000000;
			default : rdata = 44'b00000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 19) begin
	always @(*) begin
		case(address)
			// PEs: 19, 19 -> 18
			// srcs: (1, 0)(26) 7, (227) 0 --> (427) 0:ND0, NW0, *, PEGB2
			8'd0 : rdata = 44'b00011011000000000100000000000000000010100000;
			// PEs: 19, 19 -> 20
			// srcs: (2, 1)(104) 1, (305) 3 --> (505) 3:ND1, NW1, *, PENB
			8'd1 : rdata = 44'b00011011000000010100000000100000000100000000;
			// PEs: 19, 19 -> 20
			// srcs: (3, 2)(181) 4, (382) 6 --> (582) 24:ND2, NW2, *, PENB
			8'd2 : rdata = 44'b00011011000000100100000001000000000100000000;
			// PEs: 19, 19 -> 19
			// srcs: (4, 3)(150) 7, (351) 3 --> (551) 21:ND3, NW3, *, NI0
			8'd3 : rdata = 44'b00011011000000110100000001110000000000000000;
			// PEs: 22 -> 
			// srcs: (6, 4)(431) 16 --> (431) 16:PEGB6, pass, 
			8'd4 : rdata = 44'b11000111000011000000000000000000000000000000;
			// PEs: 21, 19 -> 16
			// srcs: (9, 5)(430) 7, (431) 16 --> (629) 23:PEGB5, ALU, +, PEGB0
			8'd5 : rdata = 44'b00001111000010100011111111100000000010000000;
			// PEs: 19 -> 16
			// srcs: (19, 6)(551) 21 --> (551) 21:NI0, pass, PEGB0
			8'd6 : rdata = 44'b11000101000000000000000000000000000010000000;
			// PEs: 16, 19 -> 20
			// srcs: (201, 7)(805) -9, (26) 7 --> (828) -63:PEGB0, ND0, *, PENB
			8'd7 : rdata = 44'b00011111000000000110000000000000000100000000;
			// PEs: 19, 18 -> 18
			// srcs: (202, 11)(3) 1, (826) -81 --> (1026) -81:NM0, PENB, *, PEGB2
			8'd8 : rdata = 44'b00011100000000001101111111000000000010100000;
			// PEs: 19, 20 -> 19
			// srcs: (210, 15)(227) 0, (1028) -63 --> (1228) 63:NW0, PEGB4, -, NW0
			8'd9 : rdata = 44'b00010010000000001110000100000010000000000000;
			// PEs: 16, 19 -> 20
			// srcs: (279, 8)(805) -9, (104) 1 --> (906) -9:PEGB0, ND1, *, PENB
			8'd10 : rdata = 44'b00011111000000000110000000100000000100000000;
			// PEs: 19, 18 -> 18
			// srcs: (280, 12)(3) 1, (904) -45 --> (1104) -45:NM0, PENB, *, PEGB2
			8'd11 : rdata = 44'b00011100000000001101111111000000000010100000;
			// PEs: 19, 20 -> 19
			// srcs: (288, 16)(305) 3, (1106) -9 --> (1306) 12:NW1, PEGB4, -, NW1
			8'd12 : rdata = 44'b00010010000000011110000100000010010000000000;
			// PEs: 16, 19 -> 
			// srcs: (325, 9)(805) -9, (150) 7 --> (952) -63:PEGB0, ND3, *, 
			8'd13 : rdata = 44'b00011111000000000110000001100000000000000000;
			// PEs: 19, 19 -> 
			// srcs: (328, 13)(3) 1, (952) -63 --> (1152) -63:NM0, ALU, *, 
			8'd14 : rdata = 44'b00011100000000000011111111100000000000000000;
			// PEs: 19, 19 -> 19
			// srcs: (331, 17)(351) 3, (1152) -63 --> (1352) 66:NW3, ALU, -, NW3
			8'd15 : rdata = 44'b00010010000000110011111111100010110000000000;
			// PEs: 16, 19 -> 20
			// srcs: (356, 10)(805) -9, (181) 4 --> (983) -36:PEGB0, ND2, *, PENB
			8'd16 : rdata = 44'b00011111000000000110000001000000000100000000;
			// PEs: 19, 18 -> 18
			// srcs: (358, 14)(3) 1, (982) -54 --> (1182) -54:NM0, PENB, *, PEGB2
			8'd17 : rdata = 44'b00011100000000001101111111000000000010100000;
			// PEs: 19, 20 -> 19
			// srcs: (365, 18)(382) 6, (1183) -36 --> (1383) 42:NW2, PEGB4, -, NW2
			8'd18 : rdata = 44'b00010010000000101110000100000010100000000000;
			default : rdata = 44'b00000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 20) begin
	always @(*) begin
		case(address)
			// PEs: 20, 20 -> 18
			// srcs: (1, 0)(27) 6, (228) 8 --> (428) 48:ND0, NW0, *, PEGB2
			8'd0 : rdata = 44'b00011011000000000100000000000000000010100000;
			// PEs: 20, 20 -> 20
			// srcs: (2, 1)(105) 0, (306) 4 --> (506) 0:ND1, NW1, *, NI0
			8'd1 : rdata = 44'b00011011000000010100000000110000000000000000;
			// PEs: 20, 20 -> 20
			// srcs: (3, 2)(182) 1, (383) 0 --> (583) 0:ND2, NW2, *, NI1
			8'd2 : rdata = 44'b00011011000000100100000001010100000000000000;
			// PEs: 20, 20 -> 16
			// srcs: (4, 3)(153) 7, (354) 2 --> (554) 14:ND3, NW3, *, PEGB0
			8'd3 : rdata = 44'b00011011000000110100000001100000000010000000;
			// PEs: 19, 20 -> 23
			// srcs: (5, 4)(505) 3, (506) 0 --> (704) 3:PENB, NI0, +, PEGB7
			8'd4 : rdata = 44'b00001110111111101010000000000000000011110000;
			// PEs: 19, 20 -> 21
			// srcs: (6, 5)(582) 24, (583) 0 --> (778) 24:PENB, NI1, +, PENB
			8'd5 : rdata = 44'b00001110111111101010000000100000000100000000;
			// PEs: 16, 20 -> 20
			// srcs: (202, 6)(805) -9, (27) 6 --> (829) -54:PEGB0, ND0, *, NI0
			8'd6 : rdata = 44'b00011111000000000110000000010000000000000000;
			// PEs: 20, 19 -> 19
			// srcs: (204, 10)(3) 1, (828) -63 --> (1028) -63:NM0, PENB, *, PEGB3
			8'd7 : rdata = 44'b00011100000000001101111111000000000010110000;
			// PEs: 20, 20 -> 
			// srcs: (205, 11)(3) 1, (829) -54 --> (1029) -54:NM0, NI0, *, 
			8'd8 : rdata = 44'b00011100000000001010000000000000000000000000;
			// PEs: 20, 20 -> 20
			// srcs: (208, 15)(228) 8, (1029) -54 --> (1229) 62:NW0, ALU, -, NW0
			8'd9 : rdata = 44'b00010010000000000011111111100010000000000000;
			// PEs: 16, 20 -> 21
			// srcs: (280, 7)(805) -9, (105) 0 --> (907) 0:PEGB0, ND1, *, PENB
			8'd10 : rdata = 44'b00011111000000000110000000100000000100000000;
			// PEs: 20, 19 -> 19
			// srcs: (282, 12)(3) 1, (906) -9 --> (1106) -9:NM0, PENB, *, PEGB3
			8'd11 : rdata = 44'b00011100000000001101111111000000000010110000;
			// PEs: 20, 21 -> 20
			// srcs: (289, 16)(306) 4, (1107) 0 --> (1307) 4:NW1, PEGB5, -, NW1
			8'd12 : rdata = 44'b00010010000000011110000101000010010000000000;
			// PEs: 16, 20 -> 
			// srcs: (328, 8)(805) -9, (153) 7 --> (955) -63:PEGB0, ND3, *, 
			8'd13 : rdata = 44'b00011111000000000110000001100000000000000000;
			// PEs: 20, 20 -> 
			// srcs: (331, 13)(3) 1, (955) -63 --> (1155) -63:NM0, ALU, *, 
			8'd14 : rdata = 44'b00011100000000000011111111100000000000000000;
			// PEs: 20, 20 -> 20
			// srcs: (334, 17)(354) 2, (1155) -63 --> (1355) 65:NW3, ALU, -, NW3
			8'd15 : rdata = 44'b00010010000000110011111111100010110000000000;
			// PEs: 16, 20 -> 21
			// srcs: (357, 9)(805) -9, (182) 1 --> (984) -9:PEGB0, ND2, *, PENB
			8'd16 : rdata = 44'b00011111000000000110000001000000000100000000;
			// PEs: 20, 19 -> 19
			// srcs: (359, 14)(3) 1, (983) -36 --> (1183) -36:NM0, PENB, *, PEGB3
			8'd17 : rdata = 44'b00011100000000001101111111000000000010110000;
			// PEs: 20, 21 -> 20
			// srcs: (366, 18)(383) 0, (1184) -9 --> (1384) 9:NW2, PEGB5, -, NW2
			8'd18 : rdata = 44'b00010010000000101110000101000010100000000000;
			default : rdata = 44'b00000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 21) begin
	always @(*) begin
		case(address)
			// PEs: 21, 21 -> 19
			// srcs: (1, 0)(29) 1, (230) 7 --> (430) 7:ND0, NW0, *, PEGB3
			8'd0 : rdata = 44'b00011011000000000100000000000000000010110000;
			// PEs: 21, 21 -> 22
			// srcs: (2, 1)(106) 8, (307) 1 --> (507) 8:ND1, NW1, *, PENB
			8'd1 : rdata = 44'b00011011000000010100000000100000000100000000;
			// PEs: 21, 21 -> 22
			// srcs: (3, 2)(183) 7, (384) 0 --> (584) 0:ND2, NW2, *, PENB
			8'd2 : rdata = 44'b00011011000000100100000001000000000100000000;
			// PEs: 21, 21 -> 16
			// srcs: (4, 3)(160) 3, (361) 6 --> (561) 18:ND3, NW3, *, PEGB0
			8'd3 : rdata = 44'b00011011000000110100000001100000000010000000;
			// PEs: 18 -> 
			// srcs: (8, 4)(581) 0 --> (581) 0:PEGB2, pass, 
			8'd4 : rdata = 44'b11000111000001000000000000000000000000000000;
			// PEs: 17, 21 -> 
			// srcs: (11, 5)(580) 18, (581) 0 --> (777) 18:PEGB1, ALU, +, 
			8'd5 : rdata = 44'b00001111000000100011111111100000000000000000;
			// PEs: 21, 20 -> 16
			// srcs: (14, 6)(777) 18, (778) 24 --> (779) 42:ALU, PENB, +, PEGB0
			8'd6 : rdata = 44'b00001001111111111101111111000000000010000000;
			// PEs: 16, 21 -> 22
			// srcs: (204, 7)(805) -9, (29) 1 --> (831) -9:PEGB0, ND0, *, PENB
			8'd7 : rdata = 44'b00011111000000000110000000000000000100000000;
			// PEs: 21, 22 -> 21
			// srcs: (213, 15)(230) 7, (1031) -9 --> (1231) 16:NW0, PEGB6, -, NW0
			8'd8 : rdata = 44'b00010010000000001110000110000010000000000000;
			// PEs: 16, 21 -> 21
			// srcs: (281, 8)(805) -9, (106) 8 --> (908) -72:PEGB0, ND1, *, NI0
			8'd9 : rdata = 44'b00011111000000000110000000110000000000000000;
			// PEs: 21, 20 -> 20
			// srcs: (283, 11)(3) 1, (907) 0 --> (1107) 0:NM0, PENB, *, PEGB4
			8'd10 : rdata = 44'b00011100000000001101111111000000000011000000;
			// PEs: 21, 21 -> 
			// srcs: (284, 12)(3) 1, (908) -72 --> (1108) -72:NM0, NI0, *, 
			8'd11 : rdata = 44'b00011100000000001010000000000000000000000000;
			// PEs: 21, 21 -> 21
			// srcs: (287, 16)(307) 1, (1108) -72 --> (1308) 73:NW1, ALU, -, NW1
			8'd12 : rdata = 44'b00010010000000010011111111100010010000000000;
			// PEs: 16, 21 -> 
			// srcs: (335, 9)(805) -9, (160) 3 --> (962) -27:PEGB0, ND3, *, 
			8'd13 : rdata = 44'b00011111000000000110000001100000000000000000;
			// PEs: 21, 21 -> 
			// srcs: (338, 13)(3) 1, (962) -27 --> (1162) -27:NM0, ALU, *, 
			8'd14 : rdata = 44'b00011100000000000011111111100000000000000000;
			// PEs: 21, 21 -> 21
			// srcs: (341, 17)(361) 6, (1162) -27 --> (1362) 33:NW3, ALU, -, NW3
			8'd15 : rdata = 44'b00010010000000110011111111100010110000000000;
			// PEs: 16, 21 -> 22
			// srcs: (358, 10)(805) -9, (183) 7 --> (985) -63:PEGB0, ND2, *, PENB
			8'd16 : rdata = 44'b00011111000000000110000001000000000100000000;
			// PEs: 21, 20 -> 20
			// srcs: (360, 14)(3) 1, (984) -9 --> (1184) -9:NM0, PENB, *, PEGB4
			8'd17 : rdata = 44'b00011100000000001101111111000000000011000000;
			// PEs: 21, 22 -> 21
			// srcs: (367, 18)(384) 0, (1185) -63 --> (1385) 63:NW2, PEGB6, -, NW2
			8'd18 : rdata = 44'b00010010000000101110000110000010100000000000;
			default : rdata = 44'b00000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 22) begin
	always @(*) begin
		case(address)
			// PEs: 22, 22 -> 19
			// srcs: (1, 0)(30) 8, (231) 2 --> (431) 16:ND0, NW0, *, PEGB3
			8'd0 : rdata = 44'b00011011000000000100000000000000000010110000;
			// PEs: 22, 22 -> 22
			// srcs: (2, 1)(107) 0, (308) 7 --> (508) 0:ND1, NW1, *, NI0
			8'd1 : rdata = 44'b00011011000000010100000000110000000000000000;
			// PEs: 22, 22 -> 22
			// srcs: (3, 2)(184) 8, (385) 7 --> (585) 56:ND2, NW2, *, NI1
			8'd2 : rdata = 44'b00011011000000100100000001010100000000000000;
			// PEs: 22, 22 -> 16
			// srcs: (4, 3)(163) 0, (364) 6 --> (564) 0:ND3, NW3, *, PEGB0
			8'd3 : rdata = 44'b00011011000000110100000001100000000010000000;
			// PEs: 21, 22 -> 23
			// srcs: (5, 5)(507) 8, (508) 0 --> (705) 8:PENB, NI0, +, PENB
			8'd4 : rdata = 44'b00001110111111101010000000000000000100000000;
			// PEs: 21, 22 -> 16
			// srcs: (6, 4)(584) 0, (585) 56 --> (780) 56:PENB, NI1, +, PEGB0
			8'd5 : rdata = 44'b00001110111111101010000000100000000010000000;
			// PEs: 16, 22 -> 22
			// srcs: (205, 6)(805) -9, (30) 8 --> (832) -72:PEGB0, ND0, *, NI0
			8'd6 : rdata = 44'b00011111000000000110000000010000000000000000;
			// PEs: 22, 21 -> 21
			// srcs: (207, 10)(3) 1, (831) -9 --> (1031) -9:NM0, PENB, *, PEGB5
			8'd7 : rdata = 44'b00011100000000001101111111000000000011010000;
			// PEs: 22, 22 -> 
			// srcs: (208, 11)(3) 1, (832) -72 --> (1032) -72:NM0, NI0, *, 
			8'd8 : rdata = 44'b00011100000000001010000000000000000000000000;
			// PEs: 22, 22 -> 22
			// srcs: (211, 16)(231) 2, (1032) -72 --> (1232) 74:NW0, ALU, -, NW0
			8'd9 : rdata = 44'b00010010000000000011111111100010000000000000;
			// PEs: 16, 22 -> 
			// srcs: (282, 7)(805) -9, (107) 0 --> (909) 0:PEGB0, ND1, *, 
			8'd10 : rdata = 44'b00011111000000000110000000100000000000000000;
			// PEs: 22, 22 -> 
			// srcs: (285, 12)(3) 1, (909) 0 --> (1109) 0:NM0, ALU, *, 
			8'd11 : rdata = 44'b00011100000000000011111111100000000000000000;
			// PEs: 22, 22 -> 22
			// srcs: (288, 17)(308) 7, (1109) 0 --> (1309) 7:NW1, ALU, -, NW1
			8'd12 : rdata = 44'b00010010000000010011111111100010010000000000;
			// PEs: 16, 22 -> 
			// srcs: (338, 8)(805) -9, (163) 0 --> (965) 0:PEGB0, ND3, *, 
			8'd13 : rdata = 44'b00011111000000000110000001100000000000000000;
			// PEs: 22, 22 -> 
			// srcs: (341, 13)(3) 1, (965) 0 --> (1165) 0:NM0, ALU, *, 
			8'd14 : rdata = 44'b00011100000000000011111111100000000000000000;
			// PEs: 22, 22 -> 22
			// srcs: (344, 18)(364) 6, (1165) 0 --> (1365) 6:NW3, ALU, -, NW3
			8'd15 : rdata = 44'b00010010000000110011111111100010110000000000;
			// PEs: 16, 22 -> 22
			// srcs: (359, 9)(805) -9, (184) 8 --> (986) -72:PEGB0, ND2, *, NI0
			8'd16 : rdata = 44'b00011111000000000110000001010000000000000000;
			// PEs: 22, 21 -> 21
			// srcs: (361, 14)(3) 1, (985) -63 --> (1185) -63:NM0, PENB, *, PEGB5
			8'd17 : rdata = 44'b00011100000000001101111111000000000011010000;
			// PEs: 22, 22 -> 
			// srcs: (362, 15)(3) 1, (986) -72 --> (1186) -72:NM0, NI0, *, 
			8'd18 : rdata = 44'b00011100000000001010000000000000000000000000;
			// PEs: 22, 22 -> 22
			// srcs: (365, 19)(385) 7, (1186) -72 --> (1386) 79:NW2, ALU, -, NW2
			8'd19 : rdata = 44'b00010010000000100011111111100010100000000000;
			default : rdata = 44'b00000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 23) begin
	always @(*) begin
		case(address)
			// PEs: 23, 23 -> 23
			// srcs: (1, 0)(31) 7, (232) 8 --> (432) 56:ND0, NW0, *, NI0
			8'd0 : rdata = 44'b00011011000000000100000000010000000000000000;
			// PEs: 23, 23 -> 16
			// srcs: (2, 1)(108) 2, (309) 6 --> (509) 12:ND1, NW1, *, PENB
			8'd1 : rdata = 44'b00011011000000010100000000100000000100000000;
			// PEs: 23, 23 -> 16
			// srcs: (3, 2)(186) 4, (387) 7 --> (587) 28:ND2, NW2, *, PENB
			8'd2 : rdata = 44'b00011011000000100100000001000000000100000000;
			// PEs: 23, 23 -> 23
			// srcs: (4, 3)(166) 7, (367) 1 --> (567) 7:ND3, NW3, *, NI1
			8'd3 : rdata = 44'b00011011000000110100000001110100000000000000;
			// PEs: 23 -> 16
			// srcs: (8, 4)(432) 56 --> (432) 56:NI0, pass, PENB
			8'd4 : rdata = 44'b11000101000000000000000000000000000100000000;
			// PEs: 20, 22 -> 23
			// srcs: (11, 5)(704) 3, (705) 8 --> (706) 11:PEGB4, PENB, +, NI0
			8'd5 : rdata = 44'b00001111000010001101111111010000000000000000;
			// PEs: 23 -> 16
			// srcs: (21, 6)(567) 7 --> (567) 7:NI1, pass, PENB
			8'd6 : rdata = 44'b11000101000000010000000000000000000100000000;
			// PEs: 23 -> 16
			// srcs: (35, 7)(706) 11 --> (706) 11:NI0, pass, PENB
			8'd7 : rdata = 44'b11000101000000000000000000000000000100000000;
			// PEs: 16, 23 -> 
			// srcs: (206, 8)(805) -9, (31) 7 --> (833) -63:PEGB0, ND0, *, 
			8'd8 : rdata = 44'b00011111000000000110000000000000000000000000;
			// PEs: 23, 23 -> 
			// srcs: (209, 12)(3) 1, (833) -63 --> (1033) -63:NM0, ALU, *, 
			8'd9 : rdata = 44'b00011100000000000011111111100000000000000000;
			// PEs: 23, 23 -> 23
			// srcs: (212, 16)(232) 8, (1033) -63 --> (1233) 71:NW0, ALU, -, NW0
			8'd10 : rdata = 44'b00010010000000000011111111100010000000000000;
			// PEs: 16, 23 -> 
			// srcs: (283, 9)(805) -9, (108) 2 --> (910) -18:PEGB0, ND1, *, 
			8'd11 : rdata = 44'b00011111000000000110000000100000000000000000;
			// PEs: 23, 23 -> 
			// srcs: (286, 13)(3) 1, (910) -18 --> (1110) -18:NM0, ALU, *, 
			8'd12 : rdata = 44'b00011100000000000011111111100000000000000000;
			// PEs: 23, 23 -> 23
			// srcs: (289, 17)(309) 6, (1110) -18 --> (1310) 24:NW1, ALU, -, NW1
			8'd13 : rdata = 44'b00010010000000010011111111100010010000000000;
			// PEs: 16, 23 -> 
			// srcs: (341, 10)(805) -9, (166) 7 --> (968) -63:PEGB0, ND3, *, 
			8'd14 : rdata = 44'b00011111000000000110000001100000000000000000;
			// PEs: 23, 23 -> 
			// srcs: (344, 14)(3) 1, (968) -63 --> (1168) -63:NM0, ALU, *, 
			8'd15 : rdata = 44'b00011100000000000011111111100000000000000000;
			// PEs: 23, 23 -> 23
			// srcs: (347, 18)(367) 1, (1168) -63 --> (1368) 64:NW3, ALU, -, NW3
			8'd16 : rdata = 44'b00010010000000110011111111100010110000000000;
			// PEs: 16, 23 -> 
			// srcs: (361, 11)(805) -9, (186) 4 --> (988) -36:PEGB0, ND2, *, 
			8'd17 : rdata = 44'b00011111000000000110000001000000000000000000;
			// PEs: 23, 23 -> 
			// srcs: (364, 15)(3) 1, (988) -36 --> (1188) -36:NM0, ALU, *, 
			8'd18 : rdata = 44'b00011100000000000011111111100000000000000000;
			// PEs: 23, 23 -> 23
			// srcs: (367, 19)(387) 7, (1188) -36 --> (1388) 43:NW2, ALU, -, NW2
			8'd19 : rdata = 44'b00010010000000100011111111100010100000000000;
			default : rdata = 44'b00000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 24) begin
	always @(*) begin
		case(address)
			// PEs: 16 -> 28
			// srcs: (6, 0)(509) 12 --> (509) 12:PUNB, pass, PEGB4
			8'd0 : rdata = 44'b11000110111111110000000000000000000011000000;
			// PEs: 16 -> 25
			// srcs: (7, 1)(587) 28 --> (587) 28:PUNB, pass, PENB
			8'd1 : rdata = 44'b11000110111111110000000000000000000100000000;
			// PEs: 27 -> 16
			// srcs: (10, 8)(710) 20 --> (710) 20:PEGB3, pass, PUGB2
			8'd2 : rdata = 44'b11000111000001100000000000000000000000001010;
			// PEs: 31 -> 16
			// srcs: (11, 10)(716) 46 --> (716) 46:PENB, pass, PUGB2
			8'd3 : rdata = 44'b11000110111111100000000000000000000000001010;
			// PEs: 25 -> 0
			// srcs: (14, 4)(632) 75 --> (632) 75:PEGB1, pass, PUGB0
			8'd4 : rdata = 44'b11000111000000100000000000000000000000001000;
			// PEs: 26 -> 8
			// srcs: (15, 5)(635) 18 --> (635) 18:PEGB2, pass, PUGB1
			8'd5 : rdata = 44'b11000111000001000000000000000000000000001001;
			// PEs: 27 -> 32
			// srcs: (16, 6)(637) 30 --> (637) 30:PEGB3, pass, PUNB
			8'd6 : rdata = 44'b11000111000001100000000000000000001000000000;
			// PEs: 16 -> 25
			// srcs: (17, 2)(432) 56 --> (432) 56:PUNB, pass, PENB
			8'd7 : rdata = 44'b11000110111111110000000000000000000100000000;
			// PEs: 16 -> 25
			// srcs: (18, 3)(629) 23 --> (629) 23:PUNB, pass, PENB
			8'd8 : rdata = 44'b11000110111111110000000000000000000100000000;
			// PEs: 28 -> 56
			// srcs: (19, 7)(707) 30 --> (707) 30:PEGB4, pass, PUGB7
			8'd9 : rdata = 44'b11000111000010000000000000000000000000001111;
			// PEs: 0 -> 25
			// srcs: (20, 9)(517) 0 --> (517) 0:PUGB0, pass, PENB
			8'd10 : rdata = 44'b11000111000000010000000000000000000100000000;
			// PEs: 32 -> 24
			// srcs: (21, 11)(721) 64 --> (721) 64:PUGB4, pass, NI0
			8'd11 : rdata = 44'b11000111000010010000000000010000000000000000;
			// PEs: 8 -> 25
			// srcs: (22, 12)(526) 0 --> (526) 0:PUGB1, pass, PENB
			8'd12 : rdata = 44'b11000111000000110000000000000000000100000000;
			// PEs: 27 -> 32
			// srcs: (30, 16)(576) 42 --> (576) 42:PEGB3, pass, PUNB
			8'd13 : rdata = 44'b11000111000001100000000000000000001000000000;
			// PEs: 29 -> 32
			// srcs: (31, 19)(789) 6 --> (789) 6:PEGB5, pass, PUNB
			8'd14 : rdata = 44'b11000111000010100000000000000000001000000000;
			// PEs: 31 -> 32
			// srcs: (32, 20)(791) 67 --> (791) 67:PENB, pass, PUNB
			8'd15 : rdata = 44'b11000110111111100000000000000000001000000000;
			// PEs: 24 -> 25
			// srcs: (34, 13)(721) 64 --> (721) 64:NI0, pass, PENB
			8'd16 : rdata = 44'b11000101000000000000000000000000000100000000;
			// PEs: 8 -> 25
			// srcs: (35, 14)(765) 2 --> (765) 2:PUGB1, pass, PENB
			8'd17 : rdata = 44'b11000111000000110000000000000000000100000000;
			// PEs: 8 -> 25
			// srcs: (36, 15)(767) 67 --> (767) 67:PUGB1, pass, PENB
			8'd18 : rdata = 44'b11000111000000110000000000000000000100000000;
			// PEs: 25 -> 48
			// srcs: (37, 21)(631) 99 --> (631) 99:PEGB1, pass, PUGB6
			8'd19 : rdata = 44'b11000111000000100000000000000000000000001110;
			// PEs: 25 -> 32
			// srcs: (41, 23)(722) 64 --> (722) 64:PEGB1, pass, PUNB
			8'd20 : rdata = 44'b11000111000000100000000000000000001000000000;
			// PEs: 8 -> 25
			// srcs: (47, 17)(772) 48 --> (772) 48:PUGB1, pass, PENB
			8'd21 : rdata = 44'b11000111000000110000000000000000000100000000;
			// PEs: 16 -> 25
			// srcs: (48, 18)(780) 56 --> (780) 56:PUNB, pass, PENB
			8'd22 : rdata = 44'b11000110111111110000000000000000000100000000;
			// PEs: 16 -> 28
			// srcs: (49, 22)(711) 40 --> (711) 40:PUNB, pass, PEGB4
			8'd23 : rdata = 44'b11000110111111110000000000000000000011000000;
			// PEs: 25 -> 32
			// srcs: (54, 27)(773) 48 --> (773) 48:PEGB1, pass, PUNB
			8'd24 : rdata = 44'b11000111000000100000000000000000001000000000;
			// PEs: 26 -> 32
			// srcs: (55, 31)(769) 104 --> (769) 104:PEGB2, pass, PUNB
			8'd25 : rdata = 44'b11000111000001000000000000000000001000000000;
			// PEs: 56 -> 24
			// srcs: (60, 24)(741) 60 --> (741) 60:PUGB7, pass, NI0
			8'd26 : rdata = 44'b11000111000011110000000000010000000000000000;
			// PEs: 28 -> 56
			// srcs: (61, 29)(714) 89 --> (714) 89:PEGB4, pass, PUGB7
			8'd27 : rdata = 44'b11000111000010000000000000000000000000001111;
			// PEs: 32 -> 25
			// srcs: (78, 25)(743) 32 --> (743) 32:PUGB4, pass, PENB
			8'd28 : rdata = 44'b11000111000010010000000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (85, 26)(741) 60 --> (741) 60:NI0, pass, PENB
			8'd29 : rdata = 44'b11000101000000000000000000000000000100000000;
			// PEs: 16 -> 25
			// srcs: (86, 28)(779) 42 --> (779) 42:PUNB, pass, PENB
			8'd30 : rdata = 44'b11000110111111110000000000000000000100000000;
			// PEs: 25 -> 56
			// srcs: (92, 30)(744) 92 --> (744) 92:PEGB1, pass, PUGB7
			8'd31 : rdata = 44'b11000111000000100000000000000000000000001111;
			// PEs: 29 -> 32
			// srcs: (101, 32)(788) 274 --> (788) 274:PEGB5, pass, PUNB
			8'd32 : rdata = 44'b11000111000010100000000000000000001000000000;
			// PEs: 56 -> 24
			// srcs: (117, 33)(677) 325 --> (677) 325:PUGB7, pass, NI0
			8'd33 : rdata = 44'b11000111000011110000000000010000000000000000;
			// PEs: 16 -> 25
			// srcs: (118, 34)(701) 640 --> (701) 640:PUNB, pass, PENB
			8'd34 : rdata = 44'b11000110111111110000000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (124, 35)(677) 325 --> (677) 325:NI0, pass, PENB
			8'd35 : rdata = 44'b11000101000000000000000000000000000100000000;
			// PEs: 16 -> 25
			// srcs: (125, 36)(653) 1087 --> (653) 1087:PUNB, pass, PENB
			8'd36 : rdata = 44'b11000110111111110000000000000000000100000000;
			// PEs: 25 -> 0
			// srcs: (141, 37)(703) 2052 --> (703) 2052:PEGB1, pass, PUGB0
			8'd37 : rdata = 44'b11000111000000100000000000000000000000001000;
			// PEs: 0 -> 25
			// srcs: (202, 38)(805) -9 --> (805) -9:PUGB0, pass, PENB
			8'd38 : rdata = 44'b11000111000000010000000000000000000100000000;
			// PEs: 0 -> 26
			// srcs: (203, 39)(805) -9 --> (805) -9:PUGB0, pass, PEGB2
			8'd39 : rdata = 44'b11000111000000010000000000000000000010100000;
			// PEs: 0 -> 27
			// srcs: (204, 40)(805) -9 --> (805) -9:PUGB0, pass, PEGB3
			8'd40 : rdata = 44'b11000111000000010000000000000000000010110000;
			// PEs: 0 -> 28
			// srcs: (206, 41)(805) -9 --> (805) -9:PUGB0, pass, PEGB4
			8'd41 : rdata = 44'b11000111000000010000000000000000000011000000;
			// PEs: 0 -> 29
			// srcs: (207, 42)(805) -9 --> (805) -9:PUGB0, pass, PEGB5
			8'd42 : rdata = 44'b11000111000000010000000000000000000011010000;
			// PEs: 0 -> 30
			// srcs: (209, 43)(805) -9 --> (805) -9:PUGB0, pass, PEGB6
			8'd43 : rdata = 44'b11000111000000010000000000000000000011100000;
			// PEs: 0 -> 31
			// srcs: (210, 44)(805) -9 --> (805) -9:PUGB0, pass, PEGB7
			8'd44 : rdata = 44'b11000111000000010000000000000000000011110000;
			// PEs: 0 -> 25
			// srcs: (279, 45)(805) -9 --> (805) -9:PUGB0, pass, PENB
			8'd45 : rdata = 44'b11000111000000010000000000000000000100000000;
			// PEs: 0 -> 26
			// srcs: (281, 46)(805) -9 --> (805) -9:PUGB0, pass, PEGB2
			8'd46 : rdata = 44'b11000111000000010000000000000000000010100000;
			// PEs: 0 -> 27
			// srcs: (282, 47)(805) -9 --> (805) -9:PUGB0, pass, PEGB3
			8'd47 : rdata = 44'b11000111000000010000000000000000000010110000;
			// PEs: 0 -> 28
			// srcs: (284, 48)(805) -9 --> (805) -9:PUGB0, pass, PEGB4
			8'd48 : rdata = 44'b11000111000000010000000000000000000011000000;
			// PEs: 0 -> 29
			// srcs: (285, 49)(805) -9 --> (805) -9:PUGB0, pass, PEGB5
			8'd49 : rdata = 44'b11000111000000010000000000000000000011010000;
			// PEs: 0 -> 30
			// srcs: (287, 50)(805) -9 --> (805) -9:PUGB0, pass, PEGB6
			8'd50 : rdata = 44'b11000111000000010000000000000000000011100000;
			// PEs: 0 -> 31
			// srcs: (288, 51)(805) -9 --> (805) -9:PUGB0, pass, PEGB7
			8'd51 : rdata = 44'b11000111000000010000000000000000000011110000;
			// PEs: 0 -> 25
			// srcs: (339, 52)(805) -9 --> (805) -9:PUGB0, pass, PENB
			8'd52 : rdata = 44'b11000111000000010000000000000000000100000000;
			// PEs: 0 -> 26
			// srcs: (342, 53)(805) -9 --> (805) -9:PUGB0, pass, PEGB2
			8'd53 : rdata = 44'b11000111000000010000000000000000000010100000;
			// PEs: 0 -> 27
			// srcs: (345, 54)(805) -9 --> (805) -9:PUGB0, pass, PEGB3
			8'd54 : rdata = 44'b11000111000000010000000000000000000010110000;
			// PEs: 0 -> 28
			// srcs: (348, 55)(805) -9 --> (805) -9:PUGB0, pass, PEGB4
			8'd55 : rdata = 44'b11000111000000010000000000000000000011000000;
			// PEs: 0 -> 29
			// srcs: (355, 56)(805) -9 --> (805) -9:PUGB0, pass, PEGB5
			8'd56 : rdata = 44'b11000111000000010000000000000000000011010000;
			// PEs: 0 -> 25
			// srcs: (357, 57)(805) -9 --> (805) -9:PUGB0, pass, PENB
			8'd57 : rdata = 44'b11000111000000010000000000000000000100000000;
			// PEs: 0 -> 30
			// srcs: (358, 58)(805) -9 --> (805) -9:PUGB0, pass, PEGB6
			8'd58 : rdata = 44'b11000111000000010000000000000000000011100000;
			// PEs: 0 -> 26
			// srcs: (359, 59)(805) -9 --> (805) -9:PUGB0, pass, PEGB2
			8'd59 : rdata = 44'b11000111000000010000000000000000000010100000;
			// PEs: 0 -> 27
			// srcs: (360, 60)(805) -9 --> (805) -9:PUGB0, pass, PEGB3
			8'd60 : rdata = 44'b11000111000000010000000000000000000010110000;
			// PEs: 0 -> 31
			// srcs: (361, 61)(805) -9 --> (805) -9:PUGB0, pass, PEGB7
			8'd61 : rdata = 44'b11000111000000010000000000000000000011110000;
			// PEs: 0 -> 28
			// srcs: (362, 62)(805) -9 --> (805) -9:PUGB0, pass, PEGB4
			8'd62 : rdata = 44'b11000111000000010000000000000000000011000000;
			// PEs: 0 -> 29
			// srcs: (363, 63)(805) -9 --> (805) -9:PUGB0, pass, PEGB5
			8'd63 : rdata = 44'b11000111000000010000000000000000000011010000;
			// PEs: 0 -> 30
			// srcs: (365, 64)(805) -9 --> (805) -9:PUGB0, pass, PEGB6
			8'd64 : rdata = 44'b11000111000000010000000000000000000011100000;
			// PEs: 0 -> 31
			// srcs: (366, 65)(805) -9 --> (805) -9:PUGB0, pass, PEGB7
			8'd65 : rdata = 44'b11000111000000010000000000000000000011110000;
			default : rdata = 44'b00000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 25) begin
	always @(*) begin
		case(address)
			// PEs: 25, 25 -> 25
			// srcs: (1, 0)(32) 5, (233) 4 --> (433) 20:ND0, NW0, *, NI0
			8'd0 : rdata = 44'b00011011000000000100000000010000000000000000;
			// PEs: 25, 25 -> 28
			// srcs: (2, 1)(109) 2, (310) 9 --> (510) 18:ND1, NW1, *, PEGB4
			8'd1 : rdata = 44'b00011011000000010100000000100000000011000000;
			// PEs: 25, 25 -> 25
			// srcs: (3, 2)(187) 2, (388) 9 --> (588) 18:ND2, NW2, *, NI1
			8'd2 : rdata = 44'b00011011000000100100000001010100000000000000;
			// PEs: 25, 25 -> 25
			// srcs: (4, 3)(169) 8, (370) 4 --> (570) 32:ND3, NW3, *, NI2
			8'd3 : rdata = 44'b00011011000000110100000001111000000000000000;
			// PEs: 27 -> 
			// srcs: (6, 4)(435) 45 --> (435) 45:PEGB3, pass, 
			8'd4 : rdata = 44'b11000111000001100000000000000000000000000000;
			// PEs: 26, 25 -> 24
			// srcs: (9, 5)(434) 30, (435) 45 --> (632) 75:PEGB2, ALU, +, PEGB0
			8'd5 : rdata = 44'b00001111000001000011111111100000000010000000;
			// PEs: 24, 25 -> 26
			// srcs: (10, 6)(587) 28, (588) 18 --> (783) 46:PENB, NI1, +, PENB
			8'd6 : rdata = 44'b00001110111111101010000000100000000100000000;
			// PEs: 24, 25 -> 
			// srcs: (19, 7)(432) 56, (433) 20 --> (630) 76:PENB, NI0, +, 
			8'd7 : rdata = 44'b00001110111111101010000000000000000000000000;
			// PEs: 24, 25 -> 24
			// srcs: (29, 8)(629) 23, (630) 76 --> (631) 99:PENB, ALU, +, PEGB0
			8'd8 : rdata = 44'b00001110111111100011111111100000000010000000;
			// PEs: 29, 24 -> 28
			// srcs: (30, 9)(712) 49, (517) 0 --> (713) 49:PEGB5, PENB, +, PEGB4
			8'd9 : rdata = 44'b00001111000010101101111111000000000011000000;
			// PEs: 24 -> 
			// srcs: (31, 10)(526) 0 --> (526) 0:PENB, pass, 
			8'd10 : rdata = 44'b11000110111111100000000000000000000000000000;
			// PEs: 24, 25 -> 24
			// srcs: (36, 11)(721) 64, (526) 0 --> (722) 64:PENB, ALU, +, PEGB0
			8'd11 : rdata = 44'b00001110111111100011111111100000000010000000;
			// PEs: 24, 25 -> 25
			// srcs: (37, 12)(765) 2, (570) 32 --> (766) 34:PENB, NI2, +, NI0
			8'd12 : rdata = 44'b00001110111111101010000001010000000000000000;
			// PEs: 24, 26 -> 26
			// srcs: (38, 13)(767) 67, (573) 3 --> (768) 70:PENB, PEGB2, +, PENB
			8'd13 : rdata = 44'b00001110111111101110000010000000000100000000;
			// PEs: 25 -> 26
			// srcs: (45, 18)(766) 34 --> (766) 34:NI0, pass, PENB
			8'd14 : rdata = 44'b11000101000000000000000000000000000100000000;
			// PEs: 24, 28 -> 24
			// srcs: (49, 14)(772) 48, (579) 0 --> (773) 48:PENB, PEGB4, +, PEGB0
			8'd15 : rdata = 44'b00001110111111101110000100000000000010000000;
			// PEs: 24, 29 -> 25
			// srcs: (57, 15)(780) 56, (586) 5 --> (781) 61:PENB, PEGB5, +, NI0
			8'd16 : rdata = 44'b00001110111111101110000101010000000000000000;
			// PEs: 24 -> 
			// srcs: (80, 16)(743) 32 --> (743) 32:PENB, pass, 
			8'd17 : rdata = 44'b11000110111111100000000000000000000000000000;
			// PEs: 24, 25 -> 24
			// srcs: (87, 17)(741) 60, (743) 32 --> (744) 92:PENB, ALU, +, PEGB0
			8'd18 : rdata = 44'b00001110111111100011111111100000000010000000;
			// PEs: 24, 25 -> 29
			// srcs: (88, 19)(779) 42, (781) 61 --> (782) 103:PENB, NI0, +, PEGB5
			8'd19 : rdata = 44'b00001110111111101010000000000000000011010000;
			// PEs: 24 -> 
			// srcs: (120, 20)(701) 640 --> (701) 640:PENB, pass, 
			8'd20 : rdata = 44'b11000110111111100000000000000000000000000000;
			// PEs: 24, 25 -> 
			// srcs: (126, 21)(677) 325, (701) 640 --> (702) 965:PENB, ALU, +, 
			8'd21 : rdata = 44'b00001110111111100011111111100000000000000000;
			// PEs: 24, 25 -> 24
			// srcs: (136, 22)(653) 1087, (702) 965 --> (703) 2052:PENB, ALU, +, PEGB0
			8'd22 : rdata = 44'b00001110111111100011111111100000000010000000;
			// PEs: 24, 25 -> 26
			// srcs: (204, 23)(805) -9, (32) 5 --> (834) -45:PENB, ND0, *, PENB
			8'd23 : rdata = 44'b00011110111111100110000000000000000100000000;
			// PEs: 25, 26 -> 25
			// srcs: (213, 27)(233) 4, (1034) -45 --> (1234) 49:NW0, PEGB2, -, NW0
			8'd24 : rdata = 44'b00010010000000001110000010000010000000000000;
			// PEs: 24, 25 -> 26
			// srcs: (281, 24)(805) -9, (109) 2 --> (911) -18:PENB, ND1, *, PENB
			8'd25 : rdata = 44'b00011110111111100110000000100000000100000000;
			// PEs: 25, 26 -> 25
			// srcs: (290, 28)(310) 9, (1111) -18 --> (1311) 27:NW1, PEGB2, -, NW1
			8'd26 : rdata = 44'b00010010000000011110000010000010010000000000;
			// PEs: 24, 25 -> 26
			// srcs: (341, 25)(805) -9, (169) 8 --> (971) -72:PENB, ND3, *, PENB
			8'd27 : rdata = 44'b00011110111111100110000001100000000100000000;
			// PEs: 25, 26 -> 25
			// srcs: (350, 29)(370) 4, (1171) -72 --> (1371) 76:NW3, PEGB2, -, NW3
			8'd28 : rdata = 44'b00010010000000111110000010000010110000000000;
			// PEs: 24, 25 -> 26
			// srcs: (359, 26)(805) -9, (187) 2 --> (989) -18:PENB, ND2, *, PENB
			8'd29 : rdata = 44'b00011110111111100110000001000000000100000000;
			// PEs: 25, 26 -> 25
			// srcs: (368, 30)(388) 9, (1189) -18 --> (1389) 27:NW2, PEGB2, -, NW2
			8'd30 : rdata = 44'b00010010000000101110000010000010100000000000;
			default : rdata = 44'b00000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 26) begin
	always @(*) begin
		case(address)
			// PEs: 26, 26 -> 25
			// srcs: (1, 0)(33) 5, (234) 6 --> (434) 30:ND0, NW0, *, PEGB1
			8'd0 : rdata = 44'b00011011000000000100000000000000000010010000;
			// PEs: 26, 26 -> 27
			// srcs: (2, 1)(111) 2, (312) 4 --> (512) 8:ND1, NW1, *, PENB
			8'd1 : rdata = 44'b00011011000000010100000000100000000100000000;
			// PEs: 26, 26 -> 30
			// srcs: (3, 2)(189) 7, (390) 8 --> (590) 56:ND2, NW2, *, PEGB6
			8'd2 : rdata = 44'b00011011000000100100000001000000000011100000;
			// PEs: 26, 26 -> 25
			// srcs: (4, 3)(172) 3, (373) 1 --> (573) 3:ND3, NW3, *, PEGB1
			8'd3 : rdata = 44'b00011011000000110100000001100000000010010000;
			// PEs: 29 -> 
			// srcs: (6, 4)(438) 0 --> (438) 0:PEGB5, pass, 
			8'd4 : rdata = 44'b11000111000010100000000000000000000000000000;
			// PEs: 28, 26 -> 24
			// srcs: (9, 5)(437) 18, (438) 0 --> (635) 18:PEGB4, ALU, +, PEGB0
			8'd5 : rdata = 44'b00001111000010000011111111100000000010000000;
			// PEs: 25, 30 -> 30
			// srcs: (16, 6)(783) 46, (589) 49 --> (784) 95:PENB, PEGB6, +, PEGB6
			8'd6 : rdata = 44'b00001110111111101110000110000000000011100000;
			// PEs: 25 -> 
			// srcs: (40, 7)(768) 70 --> (768) 70:PENB, pass, 
			8'd7 : rdata = 44'b11000110111111100000000000000000000000000000;
			// PEs: 25, 26 -> 24
			// srcs: (47, 8)(766) 34, (768) 70 --> (769) 104:PENB, ALU, +, PEGB0
			8'd8 : rdata = 44'b00001110111111100011111111100000000010000000;
			// PEs: 26, 25 -> 25
			// srcs: (207, 13)(3) 1, (834) -45 --> (1034) -45:NM0, PENB, *, PEGB1
			8'd9 : rdata = 44'b00011100000000001101111111000000000010010000;
			// PEs: 24, 26 -> 27
			// srcs: (208, 9)(805) -9, (33) 5 --> (835) -45:PEGB0, ND0, *, PENB
			8'd10 : rdata = 44'b00011111000000000110000000000000000100000000;
			// PEs: 26, 27 -> 26
			// srcs: (217, 18)(234) 6, (1035) -45 --> (1235) 51:NW0, PEGB3, -, NW0
			8'd11 : rdata = 44'b00010010000000001110000011000010000000000000;
			// PEs: 26, 25 -> 25
			// srcs: (284, 14)(3) 1, (911) -18 --> (1111) -18:NM0, PENB, *, PEGB1
			8'd12 : rdata = 44'b00011100000000001101111111000000000010010000;
			// PEs: 24, 26 -> 27
			// srcs: (286, 10)(805) -9, (111) 2 --> (913) -18:PEGB0, ND1, *, PENB
			8'd13 : rdata = 44'b00011111000000000110000000100000000100000000;
			// PEs: 26, 27 -> 26
			// srcs: (295, 19)(312) 4, (1113) -18 --> (1313) 22:NW1, PEGB3, -, NW1
			8'd14 : rdata = 44'b00010010000000011110000011000010010000000000;
			// PEs: 26, 25 -> 25
			// srcs: (344, 15)(3) 1, (971) -72 --> (1171) -72:NM0, PENB, *, PEGB1
			8'd15 : rdata = 44'b00011100000000001101111111000000000010010000;
			// PEs: 24, 26 -> 
			// srcs: (347, 11)(805) -9, (172) 3 --> (974) -27:PEGB0, ND3, *, 
			8'd16 : rdata = 44'b00011111000000000110000001100000000000000000;
			// PEs: 26, 26 -> 
			// srcs: (350, 16)(3) 1, (974) -27 --> (1174) -27:NM0, ALU, *, 
			8'd17 : rdata = 44'b00011100000000000011111111100000000000000000;
			// PEs: 26, 26 -> 26
			// srcs: (353, 20)(373) 1, (1174) -27 --> (1374) 28:NW3, ALU, -, NW3
			8'd18 : rdata = 44'b00010010000000110011111111100010110000000000;
			// PEs: 26, 25 -> 25
			// srcs: (362, 17)(3) 1, (989) -18 --> (1189) -18:NM0, PENB, *, PEGB1
			8'd19 : rdata = 44'b00011100000000001101111111000000000010010000;
			// PEs: 24, 26 -> 27
			// srcs: (364, 12)(805) -9, (189) 7 --> (991) -63:PEGB0, ND2, *, PENB
			8'd20 : rdata = 44'b00011111000000000110000001000000000100000000;
			// PEs: 26, 27 -> 26
			// srcs: (373, 21)(390) 8, (1191) -63 --> (1391) 71:NW2, PEGB3, -, NW2
			8'd21 : rdata = 44'b00010010000000101110000011000010100000000000;
			default : rdata = 44'b00000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 27) begin
	always @(*) begin
		case(address)
			// PEs: 27, 27 -> 25
			// srcs: (1, 0)(34) 9, (235) 5 --> (435) 45:ND0, NW0, *, PEGB1
			8'd0 : rdata = 44'b00011011000000000100000000000000000010010000;
			// PEs: 27, 27 -> 27
			// srcs: (2, 1)(112) 6, (313) 2 --> (513) 12:ND1, NW1, *, NI0
			8'd1 : rdata = 44'b00011011000000010100000000110000000000000000;
			// PEs: 27, 27 -> 30
			// srcs: (3, 2)(190) 1, (391) 8 --> (591) 8:ND2, NW2, *, PEGB6
			8'd2 : rdata = 44'b00011011000000100100000001000000000011100000;
			// PEs: 27, 27 -> 27
			// srcs: (4, 3)(175) 6, (376) 7 --> (576) 42:ND3, NW3, *, NI1
			8'd3 : rdata = 44'b00011011000000110100000001110100000000000000;
			// PEs: 26, 27 -> 24
			// srcs: (5, 6)(512) 8, (513) 12 --> (710) 20:PENB, NI0, +, PEGB0
			8'd4 : rdata = 44'b00001110111111101010000000000000000010000000;
			// PEs: 31 -> 
			// srcs: (6, 4)(441) 30 --> (441) 30:PEGB7, pass, 
			8'd5 : rdata = 44'b11000111000011100000000000000000000000000000;
			// PEs: 30, 27 -> 24
			// srcs: (9, 5)(440) 0, (441) 30 --> (637) 30:PEGB6, ALU, +, PEGB0
			8'd6 : rdata = 44'b00001111000011000011111111100000000010000000;
			// PEs: 27 -> 24
			// srcs: (25, 7)(576) 42 --> (576) 42:NI1, pass, PEGB0
			8'd7 : rdata = 44'b11000101000000010000000000000000000010000000;
			// PEs: 24, 27 -> 28
			// srcs: (209, 8)(805) -9, (34) 9 --> (836) -81:PEGB0, ND0, *, PENB
			8'd8 : rdata = 44'b00011111000000000110000000000000000100000000;
			// PEs: 27, 26 -> 26
			// srcs: (211, 12)(3) 1, (835) -45 --> (1035) -45:NM0, PENB, *, PEGB2
			8'd9 : rdata = 44'b00011100000000001101111111000000000010100000;
			// PEs: 27, 28 -> 27
			// srcs: (218, 17)(235) 5, (1036) -81 --> (1236) 86:NW0, PEGB4, -, NW0
			8'd10 : rdata = 44'b00010010000000001110000100000010000000000000;
			// PEs: 24, 27 -> 27
			// srcs: (287, 9)(805) -9, (112) 6 --> (914) -54:PEGB0, ND1, *, NI0
			8'd11 : rdata = 44'b00011111000000000110000000110000000000000000;
			// PEs: 27, 26 -> 26
			// srcs: (289, 13)(3) 1, (913) -18 --> (1113) -18:NM0, PENB, *, PEGB2
			8'd12 : rdata = 44'b00011100000000001101111111000000000010100000;
			// PEs: 27, 27 -> 
			// srcs: (290, 14)(3) 1, (914) -54 --> (1114) -54:NM0, NI0, *, 
			8'd13 : rdata = 44'b00011100000000001010000000000000000000000000;
			// PEs: 27, 27 -> 27
			// srcs: (293, 18)(313) 2, (1114) -54 --> (1314) 56:NW1, ALU, -, NW1
			8'd14 : rdata = 44'b00010010000000010011111111100010010000000000;
			// PEs: 24, 27 -> 
			// srcs: (350, 10)(805) -9, (175) 6 --> (977) -54:PEGB0, ND3, *, 
			8'd15 : rdata = 44'b00011111000000000110000001100000000000000000;
			// PEs: 27, 27 -> 
			// srcs: (353, 15)(3) 1, (977) -54 --> (1177) -54:NM0, ALU, *, 
			8'd16 : rdata = 44'b00011100000000000011111111100000000000000000;
			// PEs: 27, 27 -> 27
			// srcs: (356, 19)(376) 7, (1177) -54 --> (1377) 61:NW3, ALU, -, NW3
			8'd17 : rdata = 44'b00010010000000110011111111100010110000000000;
			// PEs: 24, 27 -> 28
			// srcs: (365, 11)(805) -9, (190) 1 --> (992) -9:PEGB0, ND2, *, PENB
			8'd18 : rdata = 44'b00011111000000000110000001000000000100000000;
			// PEs: 27, 26 -> 26
			// srcs: (367, 16)(3) 1, (991) -63 --> (1191) -63:NM0, PENB, *, PEGB2
			8'd19 : rdata = 44'b00011100000000001101111111000000000010100000;
			// PEs: 27, 28 -> 27
			// srcs: (374, 20)(391) 8, (1192) -9 --> (1392) 17:NW2, PEGB4, -, NW2
			8'd20 : rdata = 44'b00010010000000101110000100000010100000000000;
			default : rdata = 44'b00000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 28) begin
	always @(*) begin
		case(address)
			// PEs: 28, 28 -> 26
			// srcs: (1, 0)(36) 2, (237) 9 --> (437) 18:ND0, NW0, *, PEGB2
			8'd0 : rdata = 44'b00011011000000000100000000000000000010100000;
			// PEs: 28, 28 -> 29
			// srcs: (2, 1)(114) 5, (315) 9 --> (515) 45:ND1, NW1, *, PENB
			8'd1 : rdata = 44'b00011011000000010100000000100000000100000000;
			// PEs: 28, 28 -> 29
			// srcs: (3, 2)(192) 1, (393) 2 --> (593) 2:ND2, NW2, *, PENB
			8'd2 : rdata = 44'b00011011000000100100000001000000000100000000;
			// PEs: 28, 28 -> 25
			// srcs: (4, 3)(178) 0, (379) 2 --> (579) 0:ND3, NW3, *, PEGB1
			8'd3 : rdata = 44'b00011011000000110100000001100000000010010000;
			// PEs: 24 -> 
			// srcs: (11, 4)(509) 12 --> (509) 12:PEGB0, pass, 
			8'd4 : rdata = 44'b11000111000000000000000000000000000000000000;
			// PEs: 28, 25 -> 24
			// srcs: (14, 5)(509) 12, (510) 18 --> (707) 30:ALU, PEGB1, +, PEGB0
			8'd5 : rdata = 44'b00001001111111111110000001000000000010000000;
			// PEs: 24 -> 
			// srcs: (54, 6)(711) 40 --> (711) 40:PEGB0, pass, 
			8'd6 : rdata = 44'b11000111000000000000000000000000000000000000;
			// PEs: 28, 25 -> 24
			// srcs: (56, 7)(711) 40, (713) 49 --> (714) 89:ALU, PEGB1, +, PEGB0
			8'd7 : rdata = 44'b00001001111111111110000001000000000010000000;
			// PEs: 24, 28 -> 28
			// srcs: (211, 8)(805) -9, (36) 2 --> (838) -18:PEGB0, ND0, *, NI0
			8'd8 : rdata = 44'b00011111000000000110000000010000000000000000;
			// PEs: 28, 27 -> 27
			// srcs: (212, 12)(3) 1, (836) -81 --> (1036) -81:NM0, PENB, *, PEGB3
			8'd9 : rdata = 44'b00011100000000001101111111000000000010110000;
			// PEs: 28, 28 -> 
			// srcs: (214, 13)(3) 1, (838) -18 --> (1038) -18:NM0, NI0, *, 
			8'd10 : rdata = 44'b00011100000000001010000000000000000000000000;
			// PEs: 28, 28 -> 28
			// srcs: (217, 16)(237) 9, (1038) -18 --> (1238) 27:NW0, ALU, -, NW0
			8'd11 : rdata = 44'b00010010000000000011111111100010000000000000;
			// PEs: 24, 28 -> 29
			// srcs: (289, 9)(805) -9, (114) 5 --> (916) -45:PEGB0, ND1, *, PENB
			8'd12 : rdata = 44'b00011111000000000110000000100000000100000000;
			// PEs: 28, 29 -> 28
			// srcs: (298, 17)(315) 9, (1116) -45 --> (1316) 54:NW1, PEGB5, -, NW1
			8'd13 : rdata = 44'b00010010000000011110000101000010010000000000;
			// PEs: 24, 28 -> 
			// srcs: (353, 10)(805) -9, (178) 0 --> (980) 0:PEGB0, ND3, *, 
			8'd14 : rdata = 44'b00011111000000000110000001100000000000000000;
			// PEs: 28, 28 -> 
			// srcs: (356, 14)(3) 1, (980) 0 --> (1180) 0:NM0, ALU, *, 
			8'd15 : rdata = 44'b00011100000000000011111111100000000000000000;
			// PEs: 28, 28 -> 28
			// srcs: (359, 18)(379) 2, (1180) 0 --> (1380) 2:NW3, ALU, -, NW3
			8'd16 : rdata = 44'b00010010000000110011111111100010110000000000;
			// PEs: 24, 28 -> 29
			// srcs: (367, 11)(805) -9, (192) 1 --> (994) -9:PEGB0, ND2, *, PENB
			8'd17 : rdata = 44'b00011111000000000110000001000000000100000000;
			// PEs: 28, 27 -> 27
			// srcs: (368, 15)(3) 1, (992) -9 --> (1192) -9:NM0, PENB, *, PEGB3
			8'd18 : rdata = 44'b00011100000000001101111111000000000010110000;
			// PEs: 28, 29 -> 28
			// srcs: (376, 19)(393) 2, (1194) -9 --> (1394) 11:NW2, PEGB5, -, NW2
			8'd19 : rdata = 44'b00010010000000101110000101000010100000000000;
			default : rdata = 44'b00000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 29) begin
	always @(*) begin
		case(address)
			// PEs: 29, 29 -> 26
			// srcs: (1, 0)(37) 3, (238) 0 --> (438) 0:ND0, NW0, *, PEGB2
			8'd0 : rdata = 44'b00011011000000000100000000000000000010100000;
			// PEs: 29, 29 -> 29
			// srcs: (2, 1)(115) 2, (316) 2 --> (516) 4:ND1, NW1, *, NI0
			8'd1 : rdata = 44'b00011011000000010100000000110000000000000000;
			// PEs: 29, 29 -> 29
			// srcs: (3, 2)(193) 2, (394) 2 --> (594) 4:ND2, NW2, *, NI1
			8'd2 : rdata = 44'b00011011000000100100000001010100000000000000;
			// PEs: 29, 29 -> 29
			// srcs: (4, 3)(185) 5, (386) 1 --> (586) 5:ND3, NW3, *, NI2
			8'd3 : rdata = 44'b00011011000000110100000001111000000000000000;
			// PEs: 28, 29 -> 25
			// srcs: (5, 4)(515) 45, (516) 4 --> (712) 49:PENB, NI0, +, PEGB1
			8'd4 : rdata = 44'b00001110111111101010000000000000000010010000;
			// PEs: 28, 29 -> 24
			// srcs: (6, 5)(593) 2, (594) 4 --> (789) 6:PENB, NI1, +, PEGB0
			8'd5 : rdata = 44'b00001110111111101010000000100000000010000000;
			// PEs: 29 -> 25
			// srcs: (52, 6)(586) 5 --> (586) 5:NI2, pass, PEGB1
			8'd6 : rdata = 44'b11000101000000100000000000000000000010010000;
			// PEs: 25 -> 
			// srcs: (93, 7)(782) 103 --> (782) 103:PEGB1, pass, 
			8'd7 : rdata = 44'b11000111000000100000000000000000000000000000;
			// PEs: 29, 30 -> 24
			// srcs: (96, 8)(782) 103, (787) 171 --> (788) 274:ALU, PEGB6, +, PEGB0
			8'd8 : rdata = 44'b00001001111111111110000110000000000010000000;
			// PEs: 24, 29 -> 30
			// srcs: (212, 9)(805) -9, (37) 3 --> (839) -27:PEGB0, ND0, *, PENB
			8'd9 : rdata = 44'b00011111000000000110000000000000000100000000;
			// PEs: 29, 30 -> 29
			// srcs: (221, 16)(238) 0, (1039) -27 --> (1239) 27:NW0, PEGB6, -, NW0
			8'd10 : rdata = 44'b00010010000000001110000110000010000000000000;
			// PEs: 24, 29 -> 30
			// srcs: (290, 10)(805) -9, (115) 2 --> (917) -18:PEGB0, ND1, *, PENB
			8'd11 : rdata = 44'b00011111000000000110000000100000000100000000;
			// PEs: 29, 28 -> 28
			// srcs: (292, 13)(3) 1, (916) -45 --> (1116) -45:NM0, PENB, *, PEGB4
			8'd12 : rdata = 44'b00011100000000001101111111000000000011000000;
			// PEs: 29, 30 -> 29
			// srcs: (299, 17)(316) 2, (1117) -18 --> (1317) 20:NW1, PEGB6, -, NW1
			8'd13 : rdata = 44'b00010010000000011110000110000010010000000000;
			// PEs: 24, 29 -> 
			// srcs: (360, 11)(805) -9, (185) 5 --> (987) -45:PEGB0, ND3, *, 
			8'd14 : rdata = 44'b00011111000000000110000001100000000000000000;
			// PEs: 29, 29 -> 
			// srcs: (363, 14)(3) 1, (987) -45 --> (1187) -45:NM0, ALU, *, 
			8'd15 : rdata = 44'b00011100000000000011111111100000000000000000;
			// PEs: 29, 29 -> 29
			// srcs: (366, 18)(386) 1, (1187) -45 --> (1387) 46:NW3, ALU, -, NW3
			8'd16 : rdata = 44'b00010010000000110011111111100010110000000000;
			// PEs: 24, 29 -> 30
			// srcs: (368, 12)(805) -9, (193) 2 --> (995) -18:PEGB0, ND2, *, PENB
			8'd17 : rdata = 44'b00011111000000000110000001000000000100000000;
			// PEs: 29, 28 -> 28
			// srcs: (370, 15)(3) 1, (994) -9 --> (1194) -9:NM0, PENB, *, PEGB4
			8'd18 : rdata = 44'b00011100000000001101111111000000000011000000;
			// PEs: 29, 30 -> 29
			// srcs: (377, 19)(394) 2, (1195) -18 --> (1395) 20:NW2, PEGB6, -, NW2
			8'd19 : rdata = 44'b00010010000000101110000110000010100000000000;
			default : rdata = 44'b00000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 30) begin
	always @(*) begin
		case(address)
			// PEs: 30, 30 -> 27
			// srcs: (1, 0)(39) 9, (240) 0 --> (440) 0:ND0, NW0, *, PEGB3
			8'd0 : rdata = 44'b00011011000000000100000000000000000010110000;
			// PEs: 30, 30 -> 31
			// srcs: (2, 1)(117) 6, (318) 3 --> (518) 18:ND1, NW1, *, PENB
			8'd1 : rdata = 44'b00011011000000010100000000100000000100000000;
			// PEs: 30, 30 -> 31
			// srcs: (3, 2)(195) 8, (396) 4 --> (596) 32:ND2, NW2, *, PENB
			8'd2 : rdata = 44'b00011011000000100100000001000000000100000000;
			// PEs: 30, 30 -> 26
			// srcs: (4, 3)(188) 7, (389) 7 --> (589) 49:ND3, NW3, *, PEGB2
			8'd3 : rdata = 44'b00011011000000110100000001100000000010100000;
			// PEs: 27 -> 
			// srcs: (8, 4)(591) 8 --> (591) 8:PEGB3, pass, 
			8'd4 : rdata = 44'b11000111000001100000000000000000000000000000;
			// PEs: 26, 30 -> 31
			// srcs: (11, 5)(590) 56, (591) 8 --> (785) 64:PEGB2, ALU, +, PENB
			8'd5 : rdata = 44'b00001111000001000011111111100000000100000000;
			// PEs: 26 -> 
			// srcs: (21, 6)(784) 95 --> (784) 95:PEGB2, pass, 
			8'd6 : rdata = 44'b11000111000001000000000000000000000000000000;
			// PEs: 30, 31 -> 29
			// srcs: (24, 7)(784) 95, (786) 76 --> (787) 171:ALU, PEGB7, +, PEGB5
			8'd7 : rdata = 44'b00001001111111111110000111000000000011010000;
			// PEs: 24, 30 -> 31
			// srcs: (214, 8)(805) -9, (39) 9 --> (841) -81:PEGB0, ND0, *, PENB
			8'd8 : rdata = 44'b00011111000000000110000000000000000100000000;
			// PEs: 30, 29 -> 29
			// srcs: (215, 12)(3) 1, (839) -27 --> (1039) -27:NM0, PENB, *, PEGB5
			8'd9 : rdata = 44'b00011100000000001101111111000000000011010000;
			// PEs: 30, 31 -> 30
			// srcs: (223, 17)(240) 0, (1041) -81 --> (1241) 81:NW0, PEGB7, -, NW0
			8'd10 : rdata = 44'b00010010000000001110000111000010000000000000;
			// PEs: 24, 30 -> 31
			// srcs: (292, 9)(805) -9, (117) 6 --> (919) -54:PEGB0, ND1, *, PENB
			8'd11 : rdata = 44'b00011111000000000110000000100000000100000000;
			// PEs: 30, 29 -> 29
			// srcs: (293, 13)(3) 1, (917) -18 --> (1117) -18:NM0, PENB, *, PEGB5
			8'd12 : rdata = 44'b00011100000000001101111111000000000011010000;
			// PEs: 30, 31 -> 30
			// srcs: (301, 18)(318) 3, (1119) -54 --> (1319) 57:NW1, PEGB7, -, NW1
			8'd13 : rdata = 44'b00010010000000011110000111000010010000000000;
			// PEs: 24, 30 -> 
			// srcs: (363, 10)(805) -9, (188) 7 --> (990) -63:PEGB0, ND3, *, 
			8'd14 : rdata = 44'b00011111000000000110000001100000000000000000;
			// PEs: 30, 30 -> 
			// srcs: (366, 14)(3) 1, (990) -63 --> (1190) -63:NM0, ALU, *, 
			8'd15 : rdata = 44'b00011100000000000011111111100000000000000000;
			// PEs: 30, 30 -> 30
			// srcs: (369, 19)(389) 7, (1190) -63 --> (1390) 70:NW3, ALU, -, NW3
			8'd16 : rdata = 44'b00010010000000110011111111100010110000000000;
			// PEs: 24, 30 -> 30
			// srcs: (370, 11)(805) -9, (195) 8 --> (997) -72:PEGB0, ND2, *, NI0
			8'd17 : rdata = 44'b00011111000000000110000001010000000000000000;
			// PEs: 30, 29 -> 29
			// srcs: (371, 15)(3) 1, (995) -18 --> (1195) -18:NM0, PENB, *, PEGB5
			8'd18 : rdata = 44'b00011100000000001101111111000000000011010000;
			// PEs: 30, 30 -> 
			// srcs: (373, 16)(3) 1, (997) -72 --> (1197) -72:NM0, NI0, *, 
			8'd19 : rdata = 44'b00011100000000001010000000000000000000000000;
			// PEs: 30, 30 -> 30
			// srcs: (376, 20)(396) 4, (1197) -72 --> (1397) 76:NW2, ALU, -, NW2
			8'd20 : rdata = 44'b00010010000000100011111111100010100000000000;
			default : rdata = 44'b00000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 31) begin
	always @(*) begin
		case(address)
			// PEs: 31, 31 -> 27
			// srcs: (1, 0)(40) 5, (241) 6 --> (441) 30:ND0, NW0, *, PEGB3
			8'd0 : rdata = 44'b00011011000000000100000000000000000010110000;
			// PEs: 31, 31 -> 31
			// srcs: (2, 1)(118) 7, (319) 4 --> (519) 28:ND1, NW1, *, NI0
			8'd1 : rdata = 44'b00011011000000010100000000110000000000000000;
			// PEs: 31, 31 -> 31
			// srcs: (3, 2)(196) 5, (397) 7 --> (597) 35:ND2, NW2, *, NI1
			8'd2 : rdata = 44'b00011011000000100100000001010100000000000000;
			// PEs: 31, 31 -> 31
			// srcs: (4, 3)(191) 4, (392) 3 --> (592) 12:ND3, NW3, *, NI2
			8'd3 : rdata = 44'b00011011000000110100000001111000000000000000;
			// PEs: 30, 31 -> 24
			// srcs: (5, 4)(518) 18, (519) 28 --> (716) 46:PENB, NI0, +, PENB
			8'd4 : rdata = 44'b00001110111111101010000000000000000100000000;
			// PEs: 30, 31 -> 24
			// srcs: (6, 5)(596) 32, (597) 35 --> (791) 67:PENB, NI1, +, PENB
			8'd5 : rdata = 44'b00001110111111101010000000100000000100000000;
			// PEs: 30, 31 -> 30
			// srcs: (14, 6)(785) 64, (592) 12 --> (786) 76:PENB, NI2, +, PEGB6
			8'd6 : rdata = 44'b00001110111111101010000001000000000011100000;
			// PEs: 24, 31 -> 31
			// srcs: (215, 7)(805) -9, (40) 5 --> (842) -45:PEGB0, ND0, *, NI0
			8'd7 : rdata = 44'b00011111000000000110000000010000000000000000;
			// PEs: 31, 30 -> 30
			// srcs: (217, 11)(3) 1, (841) -81 --> (1041) -81:NM0, PENB, *, PEGB6
			8'd8 : rdata = 44'b00011100000000001101111111000000000011100000;
			// PEs: 31, 31 -> 
			// srcs: (218, 12)(3) 1, (842) -45 --> (1042) -45:NM0, NI0, *, 
			8'd9 : rdata = 44'b00011100000000001010000000000000000000000000;
			// PEs: 31, 31 -> 31
			// srcs: (221, 17)(241) 6, (1042) -45 --> (1242) 51:NW0, ALU, -, NW0
			8'd10 : rdata = 44'b00010010000000000011111111100010000000000000;
			// PEs: 24, 31 -> 31
			// srcs: (293, 8)(805) -9, (118) 7 --> (920) -63:PEGB0, ND1, *, NI0
			8'd11 : rdata = 44'b00011111000000000110000000110000000000000000;
			// PEs: 31, 30 -> 30
			// srcs: (295, 13)(3) 1, (919) -54 --> (1119) -54:NM0, PENB, *, PEGB6
			8'd12 : rdata = 44'b00011100000000001101111111000000000011100000;
			// PEs: 31, 31 -> 
			// srcs: (296, 14)(3) 1, (920) -63 --> (1120) -63:NM0, NI0, *, 
			8'd13 : rdata = 44'b00011100000000001010000000000000000000000000;
			// PEs: 31, 31 -> 31
			// srcs: (299, 18)(319) 4, (1120) -63 --> (1320) 67:NW1, ALU, -, NW1
			8'd14 : rdata = 44'b00010010000000010011111111100010010000000000;
			// PEs: 24, 31 -> 
			// srcs: (366, 9)(805) -9, (191) 4 --> (993) -36:PEGB0, ND3, *, 
			8'd15 : rdata = 44'b00011111000000000110000001100000000000000000;
			// PEs: 31, 31 -> 31
			// srcs: (369, 15)(3) 1, (993) -36 --> (1193) -36:NM0, ALU, *, NI0
			8'd16 : rdata = 44'b00011100000000000011111111110000000000000000;
			// PEs: 24, 31 -> 31
			// srcs: (371, 10)(805) -9, (196) 5 --> (998) -45:PEGB0, ND2, *, NI1
			8'd17 : rdata = 44'b00011111000000000110000001010100000000000000;
			// PEs: 31, 31 -> 31
			// srcs: (372, 19)(392) 3, (1193) -36 --> (1393) 39:NW3, NI0, -, NW3
			8'd18 : rdata = 44'b00010010000000111010000000000010110000000000;
			// PEs: 31, 31 -> 
			// srcs: (374, 16)(3) 1, (998) -45 --> (1198) -45:NM0, NI1, *, 
			8'd19 : rdata = 44'b00011100000000001010000000100000000000000000;
			// PEs: 31, 31 -> 31
			// srcs: (377, 20)(397) 7, (1198) -45 --> (1398) 52:NW2, ALU, -, NW2
			8'd20 : rdata = 44'b00010010000000100011111111100010100000000000;
			default : rdata = 44'b00000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 32) begin
	always @(*) begin
		case(address)
			// PEs: 39 -> 40
			// srcs: (3, 0)(452) 0 --> (452) 0:PENB, pass, PUNB
			8'd0 : rdata = 44'b11000110111111100000000000000000001000000000;
			// PEs: 39 -> 40
			// srcs: (4, 1)(530) 18 --> (530) 18:PENB, pass, PUNB
			8'd1 : rdata = 44'b11000110111111100000000000000000001000000000;
			// PEs: 39 -> 16
			// srcs: (5, 4)(417) 0 --> (417) 0:PENB, pass, PUGB2
			8'd2 : rdata = 44'b11000110111111100000000000000000000000001010;
			// PEs: 37 -> 48
			// srcs: (8, 2)(411) 9 --> (411) 9:PEGB5, pass, PUGB6
			8'd3 : rdata = 44'b11000111000010100000000000000000000000001110;
			// PEs: 38 -> 40
			// srcs: (9, 13)(646) 36 --> (646) 36:PEGB6, pass, PUNB
			8'd4 : rdata = 44'b11000111000011000000000000000000001000000000;
			// PEs: 36 -> 24
			// srcs: (10, 15)(721) 64 --> (721) 64:PEGB4, pass, PUGB3
			8'd5 : rdata = 44'b11000111000010000000000000000000000000001011;
			// PEs: 37 -> 16
			// srcs: (14, 11)(641) 51 --> (641) 51:PEGB5, pass, PUGB2
			8'd6 : rdata = 44'b11000111000010100000000000000000000000001010;
			// PEs: 38 -> 48
			// srcs: (15, 12)(643) 63 --> (643) 63:PEGB6, pass, PUGB6
			8'd7 : rdata = 44'b11000111000011000000000000000000000000001110;
			// PEs: 8 -> 33
			// srcs: (18, 3)(611) 22 --> (611) 22:PUGB1, pass, PENB
			8'd8 : rdata = 44'b11000111000000110000000000000000000100000000;
			// PEs: 8 -> 32
			// srcs: (19, 5)(617) 112 --> (617) 112:PUGB1, pass, NI0
			8'd9 : rdata = 44'b11000111000000110000000000010000000000000000;
			// PEs: 40 -> 33
			// srcs: (20, 6)(420) 0 --> (420) 0:PUGB5, pass, PENB
			8'd10 : rdata = 44'b11000111000010110000000000000000000100000000;
			// PEs: 32 -> 33
			// srcs: (26, 7)(617) 112 --> (617) 112:NI0, pass, PENB
			8'd11 : rdata = 44'b11000101000000000000000000000000000100000000;
			// PEs: 24 -> 32
			// srcs: (27, 8)(637) 30 --> (637) 30:PUNB, pass, NI0
			8'd12 : rdata = 44'b11000110111111110000000000010000000000000000;
			// PEs: 40 -> 33
			// srcs: (28, 9)(442) 0 --> (442) 0:PUGB5, pass, PENB
			8'd13 : rdata = 44'b11000111000010110000000000000000000100000000;
			// PEs: 33 -> 40
			// srcs: (29, 25)(612) 64 --> (612) 64:PEGB1, pass, PUNB
			8'd14 : rdata = 44'b11000111000000100000000000000000001000000000;
			// PEs: 33 -> 40
			// srcs: (33, 26)(618) 112 --> (618) 112:PEGB1, pass, PUNB
			8'd15 : rdata = 44'b11000111000000100000000000000000001000000000;
			// PEs: 32 -> 33
			// srcs: (34, 10)(637) 30 --> (637) 30:NI0, pass, PENB
			8'd16 : rdata = 44'b11000101000000000000000000000000000100000000;
			// PEs: 8 -> 33
			// srcs: (41, 14)(523) 18 --> (523) 18:PUGB1, pass, PENB
			8'd17 : rdata = 44'b11000111000000110000000000000000000100000000;
			// PEs: 33 -> 8
			// srcs: (42, 27)(638) 30 --> (638) 30:PEGB1, pass, PUGB1
			8'd18 : rdata = 44'b11000111000000100000000000000000000000001001;
			// PEs: 33 -> 40
			// srcs: (48, 28)(719) 30 --> (719) 30:PEGB1, pass, PUNB
			8'd19 : rdata = 44'b11000111000000100000000000000000001000000000;
			// PEs: 8 -> 33
			// srcs: (58, 16)(529) 5 --> (529) 5:PUGB1, pass, PENB
			8'd20 : rdata = 44'b11000111000000110000000000000000000100000000;
			// PEs: 48 -> 32
			// srcs: (59, 17)(742) 32 --> (742) 32:PUGB6, pass, NI0
			8'd21 : rdata = 44'b11000111000011010000000000010000000000000000;
			// PEs: 16 -> 33
			// srcs: (60, 18)(548) 0 --> (548) 0:PUGB2, pass, PENB
			8'd22 : rdata = 44'b11000111000001010000000000000000000100000000;
			// PEs: 32 -> 33
			// srcs: (66, 19)(742) 32 --> (742) 32:NI0, pass, PENB
			8'd23 : rdata = 44'b11000101000000000000000000000000000100000000;
			// PEs: 8 -> 32
			// srcs: (67, 20)(770) 78 --> (770) 78:PUGB1, pass, NI0
			8'd24 : rdata = 44'b11000111000000110000000000010000000000000000;
			// PEs: 24 -> 33
			// srcs: (68, 21)(576) 42 --> (576) 42:PUNB, pass, PENB
			8'd25 : rdata = 44'b11000110111111110000000000000000000100000000;
			// PEs: 33 -> 24
			// srcs: (73, 30)(743) 32 --> (743) 32:PEGB1, pass, PUGB3
			8'd26 : rdata = 44'b11000111000000100000000000000000000000001011;
			// PEs: 32 -> 33
			// srcs: (74, 22)(770) 78 --> (770) 78:NI0, pass, PENB
			8'd27 : rdata = 44'b11000101000000000000000000000000000100000000;
			// PEs: 24 -> 33
			// srcs: (75, 23)(789) 6 --> (789) 6:PUNB, pass, PENB
			8'd28 : rdata = 44'b11000110111111110000000000000000000100000000;
			// PEs: 24 -> 33
			// srcs: (76, 24)(791) 67 --> (791) 67:PUNB, pass, PENB
			8'd29 : rdata = 44'b11000110111111110000000000000000000100000000;
			// PEs: 24 -> 39
			// srcs: (77, 29)(722) 64 --> (722) 64:PUNB, pass, PEGB7
			8'd30 : rdata = 44'b11000110111111110000000000000000000011110000;
			// PEs: 24 -> 33
			// srcs: (78, 31)(773) 48 --> (773) 48:PUNB, pass, PENB
			8'd31 : rdata = 44'b11000110111111110000000000000000000100000000;
			// PEs: 24 -> 33
			// srcs: (79, 33)(769) 104 --> (769) 104:PUNB, pass, PENB
			8'd32 : rdata = 44'b11000110111111110000000000000000000100000000;
			// PEs: 39 -> 40
			// srcs: (86, 32)(725) 115 --> (725) 115:PENB, pass, PUNB
			8'd33 : rdata = 44'b11000110111111100000000000000000001000000000;
			// PEs: 33 -> 0
			// srcs: (101, 34)(775) 272 --> (775) 272:PEGB1, pass, PUGB0
			8'd34 : rdata = 44'b11000111000000100000000000000000000000001000;
			// PEs: 24 -> 33
			// srcs: (103, 35)(788) 274 --> (788) 274:PUNB, pass, PENB
			8'd35 : rdata = 44'b11000110111111110000000000000000000100000000;
			// PEs: 33 -> 48
			// srcs: (115, 36)(800) 542 --> (800) 542:PEGB1, pass, PUGB6
			8'd36 : rdata = 44'b11000111000000100000000000000000000000001110;
			// PEs: 0 -> 37
			// srcs: (180, 37)(805) -9 --> (805) -9:PUGB0, pass, PEGB5
			8'd37 : rdata = 44'b11000111000000010000000000000000000011010000;
			// PEs: 0 -> 38
			// srcs: (183, 38)(805) -9 --> (805) -9:PUGB0, pass, PEGB6
			8'd38 : rdata = 44'b11000111000000010000000000000000000011100000;
			// PEs: 0 -> 39
			// srcs: (186, 39)(805) -9 --> (805) -9:PUGB0, pass, PEGB7
			8'd39 : rdata = 44'b11000111000000010000000000000000000011110000;
			// PEs: 0 -> 33
			// srcs: (212, 40)(805) -9 --> (805) -9:PUGB0, pass, PENB
			8'd40 : rdata = 44'b11000111000000010000000000000000000100000000;
			// PEs: 0 -> 34
			// srcs: (213, 41)(805) -9 --> (805) -9:PUGB0, pass, PEGB2
			8'd41 : rdata = 44'b11000111000000010000000000000000000010100000;
			// PEs: 0 -> 35
			// srcs: (215, 42)(805) -9 --> (805) -9:PUGB0, pass, PEGB3
			8'd42 : rdata = 44'b11000111000000010000000000000000000010110000;
			// PEs: 0 -> 36
			// srcs: (216, 43)(805) -9 --> (805) -9:PUGB0, pass, PEGB4
			8'd43 : rdata = 44'b11000111000000010000000000000000000011000000;
			// PEs: 0 -> 37
			// srcs: (218, 44)(805) -9 --> (805) -9:PUGB0, pass, PEGB5
			8'd44 : rdata = 44'b11000111000000010000000000000000000011010000;
			// PEs: 0 -> 38
			// srcs: (219, 45)(805) -9 --> (805) -9:PUGB0, pass, PEGB6
			8'd45 : rdata = 44'b11000111000000010000000000000000000011100000;
			// PEs: 0 -> 39
			// srcs: (221, 46)(805) -9 --> (805) -9:PUGB0, pass, PEGB7
			8'd46 : rdata = 44'b11000111000000010000000000000000000011110000;
			// PEs: 0 -> 33
			// srcs: (290, 47)(805) -9 --> (805) -9:PUGB0, pass, PENB
			8'd47 : rdata = 44'b11000111000000010000000000000000000100000000;
			// PEs: 0 -> 34
			// srcs: (291, 48)(805) -9 --> (805) -9:PUGB0, pass, PEGB2
			8'd48 : rdata = 44'b11000111000000010000000000000000000010100000;
			// PEs: 0 -> 35
			// srcs: (293, 49)(805) -9 --> (805) -9:PUGB0, pass, PEGB3
			8'd49 : rdata = 44'b11000111000000010000000000000000000010110000;
			// PEs: 0 -> 36
			// srcs: (294, 50)(805) -9 --> (805) -9:PUGB0, pass, PEGB4
			8'd50 : rdata = 44'b11000111000000010000000000000000000011000000;
			// PEs: 0 -> 37
			// srcs: (296, 51)(805) -9 --> (805) -9:PUGB0, pass, PEGB5
			8'd51 : rdata = 44'b11000111000000010000000000000000000011010000;
			// PEs: 0 -> 38
			// srcs: (297, 52)(805) -9 --> (805) -9:PUGB0, pass, PEGB6
			8'd52 : rdata = 44'b11000111000000010000000000000000000011100000;
			// PEs: 0 -> 39
			// srcs: (299, 53)(805) -9 --> (805) -9:PUGB0, pass, PEGB7
			8'd53 : rdata = 44'b11000111000000010000000000000000000011110000;
			// PEs: 0 -> 33
			// srcs: (364, 54)(805) -9 --> (805) -9:PUGB0, pass, PENB
			8'd54 : rdata = 44'b11000111000000010000000000000000000100000000;
			// PEs: 0 -> 34
			// srcs: (367, 55)(805) -9 --> (805) -9:PUGB0, pass, PEGB2
			8'd55 : rdata = 44'b11000111000000010000000000000000000010100000;
			// PEs: 0 -> 33
			// srcs: (368, 56)(805) -9 --> (805) -9:PUGB0, pass, PENB
			8'd56 : rdata = 44'b11000111000000010000000000000000000100000000;
			// PEs: 0 -> 34
			// srcs: (369, 57)(805) -9 --> (805) -9:PUGB0, pass, PEGB2
			8'd57 : rdata = 44'b11000111000000010000000000000000000010100000;
			// PEs: 0 -> 35
			// srcs: (370, 58)(805) -9 --> (805) -9:PUGB0, pass, PEGB3
			8'd58 : rdata = 44'b11000111000000010000000000000000000010110000;
			// PEs: 0 -> 35
			// srcs: (371, 59)(805) -9 --> (805) -9:PUGB0, pass, PEGB3
			8'd59 : rdata = 44'b11000111000000010000000000000000000010110000;
			// PEs: 0 -> 36
			// srcs: (372, 60)(805) -9 --> (805) -9:PUGB0, pass, PEGB4
			8'd60 : rdata = 44'b11000111000000010000000000000000000011000000;
			// PEs: 0 -> 36
			// srcs: (373, 61)(805) -9 --> (805) -9:PUGB0, pass, PEGB4
			8'd61 : rdata = 44'b11000111000000010000000000000000000011000000;
			default : rdata = 44'b00000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 33) begin
	always @(*) begin
		case(address)
			// PEs: 33, 33 -> 37
			// srcs: (1, 0)(42) 6, (243) 5 --> (443) 30:ND0, NW0, *, PEGB5
			8'd0 : rdata = 44'b00011011000000000100000000000000000011010000;
			// PEs: 33, 33 -> 34
			// srcs: (2, 1)(120) 0, (321) 7 --> (521) 0:ND1, NW1, *, PENB
			8'd1 : rdata = 44'b00011011000000010100000000100000000100000000;
			// PEs: 33, 33 -> 34
			// srcs: (3, 2)(198) 0, (399) 2 --> (599) 0:ND2, NW2, *, PENB
			8'd2 : rdata = 44'b00011011000000100100000001000000000100000000;
			// PEs: 33, 33 -> 33
			// srcs: (4, 3)(194) 6, (395) 1 --> (595) 6:ND3, NW3, *, NI0
			8'd3 : rdata = 44'b00011011000000110100000001110000000000000000;
			// PEs: 32, 38 -> 32
			// srcs: (21, 4)(611) 22, (414) 42 --> (612) 64:PENB, PEGB6, +, PEGB0
			8'd4 : rdata = 44'b00001110111111101110000110000000000010000000;
			// PEs: 32 -> 
			// srcs: (22, 5)(420) 0 --> (420) 0:PENB, pass, 
			8'd5 : rdata = 44'b11000110111111100000000000000000000000000000;
			// PEs: 32, 33 -> 32
			// srcs: (28, 6)(617) 112, (420) 0 --> (618) 112:PENB, ALU, +, PEGB0
			8'd6 : rdata = 44'b00001110111111100011111111100000000010000000;
			// PEs: 32 -> 
			// srcs: (30, 7)(442) 0 --> (442) 0:PENB, pass, 
			8'd7 : rdata = 44'b11000110111111100000000000000000000000000000;
			// PEs: 32, 33 -> 32
			// srcs: (36, 8)(637) 30, (442) 0 --> (638) 30:PENB, ALU, +, PEGB0
			8'd8 : rdata = 44'b00001110111111100011111111100000000010000000;
			// PEs: 34, 32 -> 32
			// srcs: (43, 9)(718) 12, (523) 18 --> (719) 30:PEGB2, PENB, +, PEGB0
			8'd9 : rdata = 44'b00001111000001001101111111000000000010000000;
			// PEs: 38, 32 -> 39
			// srcs: (60, 10)(723) 46, (529) 5 --> (724) 51:PEGB6, PENB, +, PEGB7
			8'd10 : rdata = 44'b00001111000011001101111111000000000011110000;
			// PEs: 32 -> 
			// srcs: (62, 11)(548) 0 --> (548) 0:PENB, pass, 
			8'd11 : rdata = 44'b11000110111111100000000000000000000000000000;
			// PEs: 32, 33 -> 32
			// srcs: (68, 12)(742) 32, (548) 0 --> (743) 32:PENB, ALU, +, PEGB0
			8'd12 : rdata = 44'b00001110111111100011111111100000000010000000;
			// PEs: 32 -> 
			// srcs: (70, 13)(576) 42 --> (576) 42:PENB, pass, 
			8'd13 : rdata = 44'b11000110111111100000000000000000000000000000;
			// PEs: 32, 33 -> 33
			// srcs: (76, 14)(770) 78, (576) 42 --> (771) 120:PENB, ALU, +, NI1
			8'd14 : rdata = 44'b00001110111111100011111111110100000000000000;
			// PEs: 32, 33 -> 33
			// srcs: (77, 15)(789) 6, (595) 6 --> (790) 12:PENB, NI0, +, NI2
			8'd15 : rdata = 44'b00001110111111101010000000011000000000000000;
			// PEs: 32, 34 -> 34
			// srcs: (85, 16)(791) 67, (598) 40 --> (792) 107:PENB, PEGB2, +, PENB
			8'd16 : rdata = 44'b00001110111111101110000010000000000100000000;
			// PEs: 33, 32 -> 33
			// srcs: (86, 17)(771) 120, (773) 48 --> (774) 168:NI1, PENB, +, NI0
			8'd17 : rdata = 44'b00001101000000011101111111010000000000000000;
			// PEs: 33 -> 34
			// srcs: (92, 18)(790) 12 --> (790) 12:NI2, pass, PENB
			8'd18 : rdata = 44'b11000101000000100000000000000000000100000000;
			// PEs: 32, 33 -> 32
			// srcs: (96, 19)(769) 104, (774) 168 --> (775) 272:PENB, NI0, +, PEGB0
			8'd19 : rdata = 44'b00001110111111101010000000000000000010000000;
			// PEs: 32, 35 -> 32
			// srcs: (110, 20)(788) 274, (799) 268 --> (800) 542:PENB, PEGB3, +, PEGB0
			8'd20 : rdata = 44'b00001110111111101110000011000000000010000000;
			// PEs: 32, 33 -> 34
			// srcs: (214, 21)(805) -9, (42) 6 --> (844) -54:PENB, ND0, *, PENB
			8'd21 : rdata = 44'b00011110111111100110000000000000000100000000;
			// PEs: 33, 34 -> 33
			// srcs: (223, 25)(243) 5, (1044) -54 --> (1244) 59:NW0, PEGB2, -, NW0
			8'd22 : rdata = 44'b00010010000000001110000010000010000000000000;
			// PEs: 32, 33 -> 34
			// srcs: (292, 22)(805) -9, (120) 0 --> (922) 0:PENB, ND1, *, PENB
			8'd23 : rdata = 44'b00011110111111100110000000100000000100000000;
			// PEs: 33, 34 -> 33
			// srcs: (301, 26)(321) 7, (1122) 0 --> (1322) 7:NW1, PEGB2, -, NW1
			8'd24 : rdata = 44'b00010010000000011110000010000010010000000000;
			// PEs: 32, 33 -> 34
			// srcs: (366, 23)(805) -9, (194) 6 --> (996) -54:PENB, ND3, *, PENB
			8'd25 : rdata = 44'b00011110111111100110000001100000000100000000;
			// PEs: 32, 33 -> 34
			// srcs: (370, 24)(805) -9, (198) 0 --> (1000) 0:PENB, ND2, *, PENB
			8'd26 : rdata = 44'b00011110111111100110000001000000000100000000;
			// PEs: 33, 34 -> 33
			// srcs: (375, 27)(395) 1, (1196) -54 --> (1396) 55:NW3, PEGB2, -, NW3
			8'd27 : rdata = 44'b00010010000000111110000010000010110000000000;
			// PEs: 33, 34 -> 33
			// srcs: (379, 28)(399) 2, (1200) 0 --> (1400) 2:NW2, PEGB2, -, NW2
			8'd28 : rdata = 44'b00010010000000101110000010000010100000000000;
			default : rdata = 44'b00000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 34) begin
	always @(*) begin
		case(address)
			// PEs: 34, 34 -> 37
			// srcs: (1, 0)(43) 3, (244) 7 --> (444) 21:ND0, NW0, *, PEGB5
			8'd0 : rdata = 44'b00011011000000000100000000000000000011010000;
			// PEs: 34, 34 -> 34
			// srcs: (2, 1)(121) 3, (322) 4 --> (522) 12:ND1, NW1, *, NI0
			8'd1 : rdata = 44'b00011011000000010100000000110000000000000000;
			// PEs: 34, 34 -> 34
			// srcs: (3, 2)(199) 6, (400) 6 --> (600) 36:ND2, NW2, *, NI1
			8'd2 : rdata = 44'b00011011000000100100000001010100000000000000;
			// PEs: 34, 34 -> 34
			// srcs: (4, 3)(197) 8, (398) 5 --> (598) 40:ND3, NW3, *, NI2
			8'd3 : rdata = 44'b00011011000000110100000001111000000000000000;
			// PEs: 33, 34 -> 33
			// srcs: (5, 4)(521) 0, (522) 12 --> (718) 12:PENB, NI0, +, PEGB1
			8'd4 : rdata = 44'b00001110111111101010000000000000000010010000;
			// PEs: 33, 34 -> 35
			// srcs: (6, 5)(599) 0, (600) 36 --> (794) 36:PENB, NI1, +, PENB
			8'd5 : rdata = 44'b00001110111111101010000000100000000100000000;
			// PEs: 34 -> 33
			// srcs: (80, 6)(598) 40 --> (598) 40:NI2, pass, PEGB1
			8'd6 : rdata = 44'b11000101000000100000000000000000000010010000;
			// PEs: 33 -> 
			// srcs: (87, 7)(792) 107 --> (792) 107:PENB, pass, 
			8'd7 : rdata = 44'b11000110111111100000000000000000000000000000;
			// PEs: 33, 34 -> 35
			// srcs: (94, 8)(790) 12, (792) 107 --> (793) 119:PENB, ALU, +, PENB
			8'd8 : rdata = 44'b00001110111111100011111111100000000100000000;
			// PEs: 34, 33 -> 33
			// srcs: (217, 13)(3) 1, (844) -54 --> (1044) -54:NM0, PENB, *, PEGB1
			8'd9 : rdata = 44'b00011100000000001101111111000000000010010000;
			// PEs: 32, 34 -> 35
			// srcs: (218, 9)(805) -9, (43) 3 --> (845) -27:PEGB0, ND0, *, PENB
			8'd10 : rdata = 44'b00011111000000000110000000000000000100000000;
			// PEs: 34, 35 -> 34
			// srcs: (227, 18)(244) 7, (1045) -27 --> (1245) 34:NW0, PEGB3, -, NW0
			8'd11 : rdata = 44'b00010010000000001110000011000010000000000000;
			// PEs: 34, 33 -> 33
			// srcs: (295, 14)(3) 1, (922) 0 --> (1122) 0:NM0, PENB, *, PEGB1
			8'd12 : rdata = 44'b00011100000000001101111111000000000010010000;
			// PEs: 32, 34 -> 35
			// srcs: (296, 10)(805) -9, (121) 3 --> (923) -27:PEGB0, ND1, *, PENB
			8'd13 : rdata = 44'b00011111000000000110000000100000000100000000;
			// PEs: 34, 35 -> 34
			// srcs: (305, 19)(322) 4, (1123) -27 --> (1323) 31:NW1, PEGB3, -, NW1
			8'd14 : rdata = 44'b00010010000000011110000011000010010000000000;
			// PEs: 34, 33 -> 33
			// srcs: (369, 15)(3) 1, (996) -54 --> (1196) -54:NM0, PENB, *, PEGB1
			8'd15 : rdata = 44'b00011100000000001101111111000000000010010000;
			// PEs: 32, 34 -> 34
			// srcs: (372, 11)(805) -9, (197) 8 --> (999) -72:PEGB0, ND3, *, NI0
			8'd16 : rdata = 44'b00011111000000000110000001110000000000000000;
			// PEs: 34, 33 -> 33
			// srcs: (373, 17)(3) 1, (1000) 0 --> (1200) 0:NM0, PENB, *, PEGB1
			8'd17 : rdata = 44'b00011100000000001101111111000000000010010000;
			// PEs: 32, 34 -> 35
			// srcs: (374, 12)(805) -9, (199) 6 --> (1001) -54:PEGB0, ND2, *, PENB
			8'd18 : rdata = 44'b00011111000000000110000001000000000100000000;
			// PEs: 34, 34 -> 
			// srcs: (375, 16)(3) 1, (999) -72 --> (1199) -72:NM0, NI0, *, 
			8'd19 : rdata = 44'b00011100000000001010000000000000000000000000;
			// PEs: 34, 34 -> 34
			// srcs: (378, 20)(398) 5, (1199) -72 --> (1399) 77:NW3, ALU, -, NW3
			8'd20 : rdata = 44'b00010010000000110011111111100010110000000000;
			// PEs: 34, 35 -> 34
			// srcs: (383, 21)(400) 6, (1201) -54 --> (1401) 60:NW2, PEGB3, -, NW2
			8'd21 : rdata = 44'b00010010000000101110000011000010100000000000;
			default : rdata = 44'b00000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 35) begin
	always @(*) begin
		case(address)
			// PEs: 35, 35 -> 38
			// srcs: (1, 0)(45) 9, (246) 7 --> (446) 63:ND0, NW0, *, PEGB6
			8'd0 : rdata = 44'b00011011000000000100000000000000000011100000;
			// PEs: 35, 35 -> 36
			// srcs: (2, 1)(123) 8, (324) 8 --> (524) 64:ND1, NW1, *, PENB
			8'd1 : rdata = 44'b00011011000000010100000000100000000100000000;
			// PEs: 35, 35 -> 36
			// srcs: (3, 2)(201) 3, (402) 2 --> (602) 6:ND2, NW2, *, PENB
			8'd2 : rdata = 44'b00011011000000100100000001000000000100000000;
			// PEs: 35, 35 -> 
			// srcs: (4, 3)(200) 1, (401) 3 --> (601) 3:ND3, NW3, *, 
			8'd3 : rdata = 44'b00011011000000110100000001100000000000000000;
			// PEs: 34, 35 -> 36
			// srcs: (9, 4)(794) 36, (601) 3 --> (795) 39:PENB, ALU, +, PENB
			8'd4 : rdata = 44'b00001110111111100011111111100000000100000000;
			// PEs: 34, 36 -> 33
			// srcs: (100, 5)(793) 119, (798) 149 --> (799) 268:PENB, PEGB4, +, PEGB1
			8'd5 : rdata = 44'b00001110111111101110000100000000000010010000;
			// PEs: 32, 35 -> 35
			// srcs: (220, 6)(805) -9, (45) 9 --> (847) -81:PEGB0, ND0, *, NI0
			8'd6 : rdata = 44'b00011111000000000110000000010000000000000000;
			// PEs: 35, 34 -> 34
			// srcs: (221, 10)(3) 1, (845) -27 --> (1045) -27:NM0, PENB, *, PEGB2
			8'd7 : rdata = 44'b00011100000000001101111111000000000010100000;
			// PEs: 35, 35 -> 
			// srcs: (223, 11)(3) 1, (847) -81 --> (1047) -81:NM0, NI0, *, 
			8'd8 : rdata = 44'b00011100000000001010000000000000000000000000;
			// PEs: 35, 35 -> 35
			// srcs: (226, 15)(246) 7, (1047) -81 --> (1247) 88:NW0, ALU, -, NW0
			8'd9 : rdata = 44'b00010010000000000011111111100010000000000000;
			// PEs: 32, 35 -> 36
			// srcs: (298, 7)(805) -9, (123) 8 --> (925) -72:PEGB0, ND1, *, PENB
			8'd10 : rdata = 44'b00011111000000000110000000100000000100000000;
			// PEs: 35, 34 -> 34
			// srcs: (299, 12)(3) 1, (923) -27 --> (1123) -27:NM0, PENB, *, PEGB2
			8'd11 : rdata = 44'b00011100000000001101111111000000000010100000;
			// PEs: 35, 36 -> 35
			// srcs: (307, 16)(324) 8, (1125) -72 --> (1325) 80:NW1, PEGB4, -, NW1
			8'd12 : rdata = 44'b00010010000000011110000100000010010000000000;
			// PEs: 32, 35 -> 35
			// srcs: (375, 8)(805) -9, (200) 1 --> (1002) -9:PEGB0, ND3, *, NI0
			8'd13 : rdata = 44'b00011111000000000110000001110000000000000000;
			// PEs: 32, 35 -> 36
			// srcs: (376, 9)(805) -9, (201) 3 --> (1003) -27:PEGB0, ND2, *, PENB
			8'd14 : rdata = 44'b00011111000000000110000001000000000100000000;
			// PEs: 35, 34 -> 34
			// srcs: (377, 13)(3) 1, (1001) -54 --> (1201) -54:NM0, PENB, *, PEGB2
			8'd15 : rdata = 44'b00011100000000001101111111000000000010100000;
			// PEs: 35, 35 -> 
			// srcs: (378, 14)(3) 1, (1002) -9 --> (1202) -9:NM0, NI0, *, 
			8'd16 : rdata = 44'b00011100000000001010000000000000000000000000;
			// PEs: 35, 35 -> 35
			// srcs: (381, 17)(401) 3, (1202) -9 --> (1402) 12:NW3, ALU, -, NW3
			8'd17 : rdata = 44'b00010010000000110011111111100010110000000000;
			// PEs: 35, 36 -> 35
			// srcs: (385, 18)(402) 2, (1203) -27 --> (1403) 29:NW2, PEGB4, -, NW2
			8'd18 : rdata = 44'b00010010000000101110000100000010100000000000;
			default : rdata = 44'b00000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 36) begin
	always @(*) begin
		case(address)
			// PEs: 36, 36 -> 38
			// srcs: (1, 0)(46) 1, (247) 0 --> (447) 0:ND0, NW0, *, PEGB6
			8'd0 : rdata = 44'b00011011000000000100000000000000000011100000;
			// PEs: 36, 36 -> 36
			// srcs: (2, 1)(124) 0, (325) 5 --> (525) 0:ND1, NW1, *, NI0
			8'd1 : rdata = 44'b00011011000000010100000000110000000000000000;
			// PEs: 36, 36 -> 36
			// srcs: (3, 2)(202) 8, (403) 9 --> (603) 72:ND2, NW2, *, NI1
			8'd2 : rdata = 44'b00011011000000100100000001010100000000000000;
			// PEs: 36, 36 -> 36
			// srcs: (4, 3)(203) 4, (404) 8 --> (604) 32:ND3, NW3, *, NI2
			8'd3 : rdata = 44'b00011011000000110100000001111000000000000000;
			// PEs: 35, 36 -> 32
			// srcs: (5, 4)(524) 64, (525) 0 --> (721) 64:PENB, NI0, +, PEGB0
			8'd4 : rdata = 44'b00001110111111101010000000000000000010000000;
			// PEs: 35, 36 -> 
			// srcs: (6, 5)(602) 6, (603) 72 --> (796) 78:PENB, NI1, +, 
			8'd5 : rdata = 44'b00001110111111101010000000100000000000000000;
			// PEs: 36, 36 -> 
			// srcs: (9, 6)(796) 78, (604) 32 --> (797) 110:ALU, NI2, +, 
			8'd6 : rdata = 44'b00001001111111111010000001000000000000000000;
			// PEs: 35, 36 -> 35
			// srcs: (12, 7)(795) 39, (797) 110 --> (798) 149:PENB, ALU, +, PEGB3
			8'd7 : rdata = 44'b00001110111111100011111111100000000010110000;
			// PEs: 32, 36 -> 37
			// srcs: (221, 8)(805) -9, (46) 1 --> (848) -9:PEGB0, ND0, *, PENB
			8'd8 : rdata = 44'b00011111000000000110000000000000000100000000;
			// PEs: 36, 37 -> 36
			// srcs: (230, 14)(247) 0, (1048) -9 --> (1248) 9:NW0, PEGB5, -, NW0
			8'd9 : rdata = 44'b00010010000000001110000101000010000000000000;
			// PEs: 32, 36 -> 37
			// srcs: (299, 9)(805) -9, (124) 0 --> (926) 0:PEGB0, ND1, *, PENB
			8'd10 : rdata = 44'b00011111000000000110000000100000000100000000;
			// PEs: 36, 35 -> 35
			// srcs: (301, 12)(3) 1, (925) -72 --> (1125) -72:NM0, PENB, *, PEGB3
			8'd11 : rdata = 44'b00011100000000001101111111000000000010110000;
			// PEs: 36, 37 -> 36
			// srcs: (308, 15)(325) 5, (1126) 0 --> (1326) 5:NW1, PEGB5, -, NW1
			8'd12 : rdata = 44'b00010010000000011110000101000010010000000000;
			// PEs: 32, 36 -> 37
			// srcs: (377, 10)(805) -9, (202) 8 --> (1004) -72:PEGB0, ND2, *, PENB
			8'd13 : rdata = 44'b00011111000000000110000001000000000100000000;
			// PEs: 32, 36 -> 37
			// srcs: (378, 11)(805) -9, (203) 4 --> (1005) -36:PEGB0, ND3, *, PENB
			8'd14 : rdata = 44'b00011111000000000110000001100000000100000000;
			// PEs: 36, 35 -> 35
			// srcs: (379, 13)(3) 1, (1003) -27 --> (1203) -27:NM0, PENB, *, PEGB3
			8'd15 : rdata = 44'b00011100000000001101111111000000000010110000;
			// PEs: 36, 37 -> 36
			// srcs: (386, 16)(403) 9, (1204) -72 --> (1404) 81:NW2, PEGB5, -, NW2
			8'd16 : rdata = 44'b00010010000000101110000101000010100000000000;
			// PEs: 36, 37 -> 36
			// srcs: (387, 17)(404) 8, (1205) -36 --> (1405) 44:NW3, PEGB5, -, NW3
			8'd17 : rdata = 44'b00010010000000111110000101000010110000000000;
			default : rdata = 44'b00000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 37) begin
	always @(*) begin
		case(address)
			// PEs: 37, 37 -> 38
			// srcs: (1, 0)(48) 4, (249) 8 --> (449) 32:ND0, NW0, *, PENB
			8'd0 : rdata = 44'b00011011000000000100000000000000000100000000;
			// PEs: 37, 37 -> 38
			// srcs: (2, 1)(126) 1, (327) 6 --> (527) 6:ND1, NW1, *, PENB
			8'd1 : rdata = 44'b00011011000000010100000000100000000100000000;
			// PEs: 37, 37 -> 32
			// srcs: (3, 2)(10) 9, (211) 1 --> (411) 9:ND2, NW2, *, PEGB0
			8'd2 : rdata = 44'b00011011000000100100000001000000000010000000;
			// PEs: 34 -> 
			// srcs: (6, 3)(444) 21 --> (444) 21:PEGB2, pass, 
			8'd3 : rdata = 44'b11000111000001000000000000000000000000000000;
			// PEs: 33, 37 -> 32
			// srcs: (9, 4)(443) 30, (444) 21 --> (641) 51:PEGB1, ALU, +, PEGB0
			8'd4 : rdata = 44'b00001111000000100011111111100000000010000000;
			// PEs: 32, 37 -> 
			// srcs: (185, 5)(805) -9, (10) 9 --> (812) -81:PEGB0, ND2, *, 
			8'd5 : rdata = 44'b00011111000000000110000001000000000000000000;
			// PEs: 37, 37 -> 
			// srcs: (188, 8)(3) 1, (812) -81 --> (1012) -81:NM0, ALU, *, 
			8'd6 : rdata = 44'b00011100000000000011111111100000000000000000;
			// PEs: 37, 37 -> 37
			// srcs: (191, 14)(211) 1, (1012) -81 --> (1212) 82:NW2, ALU, -, NW2
			8'd7 : rdata = 44'b00010010000000100011111111100010100000000000;
			// PEs: 32, 37 -> 37
			// srcs: (223, 6)(805) -9, (48) 4 --> (850) -36:PEGB0, ND0, *, NI0
			8'd8 : rdata = 44'b00011111000000000110000000010000000000000000;
			// PEs: 37, 36 -> 36
			// srcs: (224, 9)(3) 1, (848) -9 --> (1048) -9:NM0, PENB, *, PEGB4
			8'd9 : rdata = 44'b00011100000000001101111111000000000011000000;
			// PEs: 37, 37 -> 
			// srcs: (226, 10)(3) 1, (850) -36 --> (1050) -36:NM0, NI0, *, 
			8'd10 : rdata = 44'b00011100000000001010000000000000000000000000;
			// PEs: 37, 37 -> 37
			// srcs: (229, 15)(249) 8, (1050) -36 --> (1250) 44:NW0, ALU, -, NW0
			8'd11 : rdata = 44'b00010010000000000011111111100010000000000000;
			// PEs: 32, 37 -> 38
			// srcs: (301, 7)(805) -9, (126) 1 --> (928) -9:PEGB0, ND1, *, PENB
			8'd12 : rdata = 44'b00011111000000000110000000100000000100000000;
			// PEs: 37, 36 -> 36
			// srcs: (302, 11)(3) 1, (926) 0 --> (1126) 0:NM0, PENB, *, PEGB4
			8'd13 : rdata = 44'b00011100000000001101111111000000000011000000;
			// PEs: 37, 38 -> 37
			// srcs: (310, 16)(327) 6, (1128) -9 --> (1328) 15:NW1, PEGB6, -, NW1
			8'd14 : rdata = 44'b00010010000000011110000110000010010000000000;
			// PEs: 37, 36 -> 36
			// srcs: (380, 12)(3) 1, (1004) -72 --> (1204) -72:NM0, PENB, *, PEGB4
			8'd15 : rdata = 44'b00011100000000001101111111000000000011000000;
			// PEs: 37, 36 -> 36
			// srcs: (381, 13)(3) 1, (1005) -36 --> (1205) -36:NM0, PENB, *, PEGB4
			8'd16 : rdata = 44'b00011100000000001101111111000000000011000000;
			default : rdata = 44'b00000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 38) begin
	always @(*) begin
		case(address)
			// PEs: 38, 38 -> 38
			// srcs: (1, 0)(49) 4, (250) 1 --> (450) 4:ND0, NW0, *, NI0
			8'd0 : rdata = 44'b00011011000000000100000000010000000000000000;
			// PEs: 38, 38 -> 38
			// srcs: (2, 1)(127) 8, (328) 5 --> (528) 40:ND1, NW1, *, NI1
			8'd1 : rdata = 44'b00011011000000010100000000110100000000000000;
			// PEs: 38, 38 -> 33
			// srcs: (3, 2)(13) 6, (214) 7 --> (414) 42:ND2, NW2, *, PEGB1
			8'd2 : rdata = 44'b00011011000000100100000001000000000010010000;
			// PEs: 37, 38 -> 32
			// srcs: (4, 5)(449) 32, (450) 4 --> (646) 36:PENB, NI0, +, PEGB0
			8'd3 : rdata = 44'b00001110111111101010000000000000000010000000;
			// PEs: 37, 38 -> 33
			// srcs: (5, 6)(527) 6, (528) 40 --> (723) 46:PENB, NI1, +, PEGB1
			8'd4 : rdata = 44'b00001110111111101010000000100000000010010000;
			// PEs: 36 -> 
			// srcs: (6, 3)(447) 0 --> (447) 0:PEGB4, pass, 
			8'd5 : rdata = 44'b11000111000010000000000000000000000000000000;
			// PEs: 35, 38 -> 32
			// srcs: (9, 4)(446) 63, (447) 0 --> (643) 63:PEGB3, ALU, +, PEGB0
			8'd6 : rdata = 44'b00001111000001100011111111100000000010000000;
			// PEs: 32, 38 -> 
			// srcs: (188, 7)(805) -9, (13) 6 --> (815) -54:PEGB0, ND2, *, 
			8'd7 : rdata = 44'b00011111000000000110000001000000000000000000;
			// PEs: 38, 38 -> 
			// srcs: (191, 10)(3) 1, (815) -54 --> (1015) -54:NM0, ALU, *, 
			8'd8 : rdata = 44'b00011100000000000011111111100000000000000000;
			// PEs: 38, 38 -> 38
			// srcs: (194, 12)(214) 7, (1015) -54 --> (1215) 61:NW2, ALU, -, NW2
			8'd9 : rdata = 44'b00010010000000100011111111100010100000000000;
			// PEs: 32, 38 -> 39
			// srcs: (224, 8)(805) -9, (49) 4 --> (851) -36:PEGB0, ND0, *, PENB
			8'd10 : rdata = 44'b00011111000000000110000000000000000100000000;
			// PEs: 38, 39 -> 38
			// srcs: (233, 13)(250) 1, (1051) -36 --> (1251) 37:NW0, PEGB7, -, NW0
			8'd11 : rdata = 44'b00010010000000001110000111000010000000000000;
			// PEs: 32, 38 -> 39
			// srcs: (302, 9)(805) -9, (127) 8 --> (929) -72:PEGB0, ND1, *, PENB
			8'd12 : rdata = 44'b00011111000000000110000000100000000100000000;
			// PEs: 38, 37 -> 37
			// srcs: (304, 11)(3) 1, (928) -9 --> (1128) -9:NM0, PENB, *, PEGB5
			8'd13 : rdata = 44'b00011100000000001101111111000000000011010000;
			// PEs: 38, 39 -> 38
			// srcs: (311, 14)(328) 5, (1129) -72 --> (1329) 77:NW1, PEGB7, -, NW1
			8'd14 : rdata = 44'b00010010000000011110000111000010010000000000;
			default : rdata = 44'b00000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 39) begin
	always @(*) begin
		case(address)
			// PEs: 39, 39 -> 32
			// srcs: (1, 0)(51) 0, (252) 3 --> (452) 0:ND0, NW0, *, PENB
			8'd0 : rdata = 44'b00011011000000000100000000000000000100000000;
			// PEs: 39, 39 -> 32
			// srcs: (2, 1)(129) 9, (330) 2 --> (530) 18:ND1, NW1, *, PENB
			8'd1 : rdata = 44'b00011011000000010100000000100000000100000000;
			// PEs: 39, 39 -> 32
			// srcs: (3, 2)(16) 0, (217) 7 --> (417) 0:ND2, NW2, *, PENB
			8'd2 : rdata = 44'b00011011000000100100000001000000000100000000;
			// PEs: 32 -> 
			// srcs: (82, 3)(722) 64 --> (722) 64:PEGB0, pass, 
			8'd3 : rdata = 44'b11000111000000000000000000000000000000000000;
			// PEs: 39, 33 -> 32
			// srcs: (84, 4)(722) 64, (724) 51 --> (725) 115:ALU, PEGB1, +, PENB
			8'd4 : rdata = 44'b00001001111111111110000001000000000100000000;
			// PEs: 32, 39 -> 
			// srcs: (191, 5)(805) -9, (16) 0 --> (818) 0:PEGB0, ND2, *, 
			8'd5 : rdata = 44'b00011111000000000110000001000000000000000000;
			// PEs: 39, 39 -> 
			// srcs: (194, 8)(3) 1, (818) 0 --> (1018) 0:NM0, ALU, *, 
			8'd6 : rdata = 44'b00011100000000000011111111100000000000000000;
			// PEs: 39, 39 -> 39
			// srcs: (197, 13)(217) 7, (1018) 0 --> (1218) 7:NW2, ALU, -, NW2
			8'd7 : rdata = 44'b00010010000000100011111111100010100000000000;
			// PEs: 32, 39 -> 39
			// srcs: (226, 6)(805) -9, (51) 0 --> (853) 0:PEGB0, ND0, *, NI0
			8'd8 : rdata = 44'b00011111000000000110000000010000000000000000;
			// PEs: 39, 38 -> 38
			// srcs: (227, 9)(3) 1, (851) -36 --> (1051) -36:NM0, PENB, *, PEGB6
			8'd9 : rdata = 44'b00011100000000001101111111000000000011100000;
			// PEs: 39, 39 -> 
			// srcs: (229, 10)(3) 1, (853) 0 --> (1053) 0:NM0, NI0, *, 
			8'd10 : rdata = 44'b00011100000000001010000000000000000000000000;
			// PEs: 39, 39 -> 39
			// srcs: (232, 14)(252) 3, (1053) 0 --> (1253) 3:NW0, ALU, -, NW0
			8'd11 : rdata = 44'b00010010000000000011111111100010000000000000;
			// PEs: 32, 39 -> 39
			// srcs: (304, 7)(805) -9, (129) 9 --> (931) -81:PEGB0, ND1, *, NI0
			8'd12 : rdata = 44'b00011111000000000110000000110000000000000000;
			// PEs: 39, 38 -> 38
			// srcs: (305, 11)(3) 1, (929) -72 --> (1129) -72:NM0, PENB, *, PEGB6
			8'd13 : rdata = 44'b00011100000000001101111111000000000011100000;
			// PEs: 39, 39 -> 
			// srcs: (307, 12)(3) 1, (931) -81 --> (1131) -81:NM0, NI0, *, 
			8'd14 : rdata = 44'b00011100000000001010000000000000000000000000;
			// PEs: 39, 39 -> 39
			// srcs: (310, 15)(330) 2, (1131) -81 --> (1331) 83:NW1, ALU, -, NW1
			8'd15 : rdata = 44'b00010010000000010011111111100010010000000000;
			default : rdata = 44'b00000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 40) begin
	always @(*) begin
		case(address)
			// PEs: 32 -> 41
			// srcs: (5, 0)(452) 0 --> (452) 0:PUNB, pass, PENB
			8'd0 : rdata = 44'b11000110111111110000000000000000000100000000;
			// PEs: 32 -> 41
			// srcs: (6, 1)(530) 18 --> (530) 18:PUNB, pass, PENB
			8'd1 : rdata = 44'b11000110111111110000000000000000000100000000;
			// PEs: 41 -> 32
			// srcs: (8, 2)(420) 0 --> (420) 0:PEGB1, pass, PUGB4
			8'd2 : rdata = 44'b11000111000000100000000000000000000000001100;
			// PEs: 43 -> 48
			// srcs: (9, 4)(426) 0 --> (426) 0:PEGB3, pass, PUNB
			8'd3 : rdata = 44'b11000111000001100000000000000000001000000000;
			// PEs: 44 -> 56
			// srcs: (10, 5)(429) 4 --> (429) 4:PEGB4, pass, PUGB7
			8'd4 : rdata = 44'b11000111000010000000000000000000000000001111;
			// PEs: 45 -> 0
			// srcs: (11, 6)(436) 9 --> (436) 9:PEGB5, pass, PUGB0
			8'd5 : rdata = 44'b11000111000010100000000000000000000000001000;
			// PEs: 46 -> 8
			// srcs: (12, 7)(439) 18 --> (439) 18:PEGB6, pass, PUGB1
			8'd6 : rdata = 44'b11000111000011000000000000000000000000001001;
			// PEs: 47 -> 32
			// srcs: (13, 8)(442) 0 --> (442) 0:PENB, pass, PUGB4
			8'd7 : rdata = 44'b11000110111111100000000000000000000000001100;
			// PEs: 41 -> 48
			// srcs: (14, 12)(648) 36 --> (648) 36:PEGB1, pass, PUNB
			8'd8 : rdata = 44'b11000111000000100000000000000000001000000000;
			// PEs: 47 -> 48
			// srcs: (15, 13)(657) 46 --> (657) 46:PENB, pass, PUNB
			8'd9 : rdata = 44'b11000110111111100000000000000000001000000000;
			// PEs: 47 -> 8
			// srcs: (16, 18)(734) 55 --> (734) 55:PENB, pass, PUGB1
			8'd10 : rdata = 44'b11000110111111100000000000000000000000001001;
			// PEs: 8 -> 41
			// srcs: (20, 3)(619) 91 --> (619) 91:PUGB1, pass, PENB
			8'd11 : rdata = 44'b11000111000000110000000000000000000100000000;
			// PEs: 32 -> 40
			// srcs: (21, 9)(646) 36 --> (646) 36:PUNB, pass, NI0
			8'd12 : rdata = 44'b11000110111111110000000000010000000000000000;
			// PEs: 48 -> 41
			// srcs: (22, 10)(451) 9 --> (451) 9:PUGB6, pass, PENB
			8'd13 : rdata = 44'b11000111000011010000000000000000000100000000;
			// PEs: 40 -> 41
			// srcs: (28, 11)(646) 36 --> (646) 36:NI0, pass, PENB
			8'd14 : rdata = 44'b11000101000000000000000000000000000100000000;
			// PEs: 16 -> 40
			// srcs: (29, 14)(697) 64 --> (697) 64:PUGB2, pass, NI0
			8'd15 : rdata = 44'b11000111000001010000000000010000000000000000;
			// PEs: 0 -> 41
			// srcs: (30, 15)(504) 5 --> (504) 5:PUGB0, pass, PENB
			8'd16 : rdata = 44'b11000111000000010000000000000000000100000000;
			// PEs: 41 -> 48
			// srcs: (35, 26)(647) 45 --> (647) 45:PEGB1, pass, PUNB
			8'd17 : rdata = 44'b11000111000000100000000000000000001000000000;
			// PEs: 40 -> 41
			// srcs: (36, 16)(697) 64 --> (697) 64:NI0, pass, PENB
			8'd18 : rdata = 44'b11000101000000000000000000000000000100000000;
			// PEs: 8 -> 41
			// srcs: (37, 17)(536) 9 --> (536) 9:PUGB1, pass, PENB
			8'd19 : rdata = 44'b11000111000000110000000000000000000100000000;
			// PEs: 56 -> 40
			// srcs: (38, 19)(747) 67 --> (747) 67:PUGB7, pass, NI0
			8'd20 : rdata = 44'b11000111000011110000000000010000000000000000;
			// PEs: 16 -> 41
			// srcs: (39, 20)(554) 14 --> (554) 14:PUGB2, pass, PENB
			8'd21 : rdata = 44'b11000111000001010000000000000000000100000000;
			// PEs: 42 -> 48
			// srcs: (40, 27)(656) 12 --> (656) 12:PEGB2, pass, PUNB
			8'd22 : rdata = 44'b11000111000001000000000000000000001000000000;
			// PEs: 41 -> 16
			// srcs: (43, 28)(698) 69 --> (698) 69:PEGB1, pass, PUGB2
			8'd23 : rdata = 44'b11000111000000100000000000000000000000001010;
			// PEs: 40 -> 41
			// srcs: (45, 21)(747) 67 --> (747) 67:NI0, pass, PENB
			8'd24 : rdata = 44'b11000101000000000000000000000000000100000000;
			// PEs: 32 -> 40
			// srcs: (46, 22)(612) 64 --> (612) 64:PUNB, pass, NI0
			8'd25 : rdata = 44'b11000110111111110000000000010000000000000000;
			// PEs: 16 -> 41
			// srcs: (47, 23)(614) 60 --> (614) 60:PUGB2, pass, PENB
			8'd26 : rdata = 44'b11000111000001010000000000000000000100000000;
			// PEs: 32 -> 46
			// srcs: (48, 25)(618) 112 --> (618) 112:PUNB, pass, PEGB6
			8'd27 : rdata = 44'b11000110111111110000000000000000000011100000;
			// PEs: 41 -> 48
			// srcs: (52, 32)(748) 81 --> (748) 81:PEGB1, pass, PUNB
			8'd28 : rdata = 44'b11000111000000100000000000000000001000000000;
			// PEs: 40 -> 41
			// srcs: (53, 24)(612) 64 --> (612) 64:NI0, pass, PENB
			8'd29 : rdata = 44'b11000101000000000000000000000000000100000000;
			// PEs: 44 -> 48
			// srcs: (54, 36)(733) 170 --> (733) 170:PEGB4, pass, PUNB
			8'd30 : rdata = 44'b11000111000010000000000000000000001000000000;
			// PEs: 16 -> 40
			// srcs: (57, 29)(717) 53 --> (717) 53:PUGB2, pass, NI0
			8'd31 : rdata = 44'b11000111000001010000000000010000000000000000;
			// PEs: 32 -> 41
			// srcs: (58, 30)(719) 30 --> (719) 30:PUNB, pass, PENB
			8'd32 : rdata = 44'b11000110111111110000000000000000000100000000;
			// PEs: 46 -> 56
			// srcs: (60, 34)(621) 218 --> (621) 218:PEGB6, pass, PUGB7
			8'd33 : rdata = 44'b11000111000011000000000000000000000000001111;
			// PEs: 40 -> 41
			// srcs: (64, 31)(717) 53 --> (717) 53:NI0, pass, PENB
			8'd34 : rdata = 44'b11000101000000000000000000000000000100000000;
			// PEs: 48 -> 41
			// srcs: (65, 33)(610) 83 --> (610) 83:PUGB6, pass, PENB
			8'd35 : rdata = 44'b11000111000011010000000000000000000100000000;
			// PEs: 41 -> 8
			// srcs: (72, 37)(616) 207 --> (616) 207:PEGB1, pass, PUGB1
			8'd36 : rdata = 44'b11000111000000100000000000000000000000001001;
			// PEs: 32 -> 41
			// srcs: (88, 35)(725) 115 --> (725) 115:PUNB, pass, PENB
			8'd37 : rdata = 44'b11000110111111110000000000000000000100000000;
			// PEs: 56 -> 41
			// srcs: (92, 38)(715) 144 --> (715) 144:PUGB7, pass, PENB
			8'd38 : rdata = 44'b11000111000011110000000000000000000100000000;
			// PEs: 56 -> 41
			// srcs: (126, 39)(751) 724 --> (751) 724:PUGB7, pass, PENB
			8'd39 : rdata = 44'b11000111000011110000000000000000000100000000;
			// PEs: 41 -> 48
			// srcs: (134, 40)(752) 1066 --> (752) 1066:PEGB1, pass, PUNB
			8'd40 : rdata = 44'b11000111000000100000000000000000001000000000;
			// PEs: 0 -> 41
			// srcs: (189, 41)(805) -9 --> (805) -9:PUGB0, pass, PENB
			8'd41 : rdata = 44'b11000111000000010000000000000000000100000000;
			// PEs: 0 -> 42
			// srcs: (192, 42)(805) -9 --> (805) -9:PUGB0, pass, PEGB2
			8'd42 : rdata = 44'b11000111000000010000000000000000000010100000;
			// PEs: 0 -> 43
			// srcs: (195, 43)(805) -9 --> (805) -9:PUGB0, pass, PEGB3
			8'd43 : rdata = 44'b11000111000000010000000000000000000010110000;
			// PEs: 0 -> 44
			// srcs: (198, 44)(805) -9 --> (805) -9:PUGB0, pass, PEGB4
			8'd44 : rdata = 44'b11000111000000010000000000000000000011000000;
			// PEs: 0 -> 45
			// srcs: (205, 45)(805) -9 --> (805) -9:PUGB0, pass, PEGB5
			8'd45 : rdata = 44'b11000111000000010000000000000000000011010000;
			// PEs: 0 -> 46
			// srcs: (208, 46)(805) -9 --> (805) -9:PUGB0, pass, PEGB6
			8'd46 : rdata = 44'b11000111000000010000000000000000000011100000;
			// PEs: 0 -> 47
			// srcs: (211, 47)(805) -9 --> (805) -9:PUGB0, pass, PEGB7
			8'd47 : rdata = 44'b11000111000000010000000000000000000011110000;
			// PEs: 0 -> 41
			// srcs: (222, 48)(805) -9 --> (805) -9:PUGB0, pass, PENB
			8'd48 : rdata = 44'b11000111000000010000000000000000000100000000;
			// PEs: 0 -> 42
			// srcs: (224, 49)(805) -9 --> (805) -9:PUGB0, pass, PEGB2
			8'd49 : rdata = 44'b11000111000000010000000000000000000010100000;
			// PEs: 0 -> 43
			// srcs: (225, 50)(805) -9 --> (805) -9:PUGB0, pass, PEGB3
			8'd50 : rdata = 44'b11000111000000010000000000000000000010110000;
			// PEs: 0 -> 44
			// srcs: (226, 51)(805) -9 --> (805) -9:PUGB0, pass, PEGB4
			8'd51 : rdata = 44'b11000111000000010000000000000000000011000000;
			// PEs: 0 -> 45
			// srcs: (227, 52)(805) -9 --> (805) -9:PUGB0, pass, PEGB5
			8'd52 : rdata = 44'b11000111000000010000000000000000000011010000;
			// PEs: 0 -> 46
			// srcs: (228, 53)(805) -9 --> (805) -9:PUGB0, pass, PEGB6
			8'd53 : rdata = 44'b11000111000000010000000000000000000011100000;
			// PEs: 0 -> 47
			// srcs: (229, 54)(805) -9 --> (805) -9:PUGB0, pass, PEGB7
			8'd54 : rdata = 44'b11000111000000010000000000000000000011110000;
			// PEs: 0 -> 41
			// srcs: (300, 55)(805) -9 --> (805) -9:PUGB0, pass, PENB
			8'd55 : rdata = 44'b11000111000000010000000000000000000100000000;
			// PEs: 0 -> 42
			// srcs: (301, 56)(805) -9 --> (805) -9:PUGB0, pass, PEGB2
			8'd56 : rdata = 44'b11000111000000010000000000000000000010100000;
			// PEs: 0 -> 43
			// srcs: (302, 57)(805) -9 --> (805) -9:PUGB0, pass, PEGB3
			8'd57 : rdata = 44'b11000111000000010000000000000000000010110000;
			// PEs: 0 -> 44
			// srcs: (303, 58)(805) -9 --> (805) -9:PUGB0, pass, PEGB4
			8'd58 : rdata = 44'b11000111000000010000000000000000000011000000;
			// PEs: 0 -> 45
			// srcs: (304, 59)(805) -9 --> (805) -9:PUGB0, pass, PEGB5
			8'd59 : rdata = 44'b11000111000000010000000000000000000011010000;
			// PEs: 0 -> 46
			// srcs: (306, 60)(805) -9 --> (805) -9:PUGB0, pass, PEGB6
			8'd60 : rdata = 44'b11000111000000010000000000000000000011100000;
			// PEs: 0 -> 47
			// srcs: (307, 61)(805) -9 --> (805) -9:PUGB0, pass, PEGB7
			8'd61 : rdata = 44'b11000111000000010000000000000000000011110000;
			default : rdata = 44'b00000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 41) begin
	always @(*) begin
		case(address)
			// PEs: 41, 41 -> 41
			// srcs: (1, 0)(52) 6, (253) 6 --> (453) 36:ND0, NW0, *, NI0
			8'd0 : rdata = 44'b00011011000000000100000000010000000000000000;
			// PEs: 41, 41 -> 41
			// srcs: (2, 1)(130) 6, (331) 6 --> (531) 36:ND1, NW1, *, NI1
			8'd1 : rdata = 44'b00011011000000010100000000110100000000000000;
			// PEs: 41, 41 -> 40
			// srcs: (3, 2)(19) 0, (220) 9 --> (420) 0:ND2, NW2, *, PEGB0
			8'd2 : rdata = 44'b00011011000000100100000001000000000010000000;
			// PEs: 40, 41 -> 40
			// srcs: (8, 3)(452) 0, (453) 36 --> (648) 36:PENB, NI0, +, PEGB0
			8'd3 : rdata = 44'b00001110111111101010000000000000000010000000;
			// PEs: 40, 41 -> 44
			// srcs: (9, 4)(530) 18, (531) 36 --> (728) 54:PENB, NI1, +, PEGB4
			8'd4 : rdata = 44'b00001110111111101010000000100000000011000000;
			// PEs: 40, 42 -> 46
			// srcs: (22, 5)(619) 91, (423) 15 --> (620) 106:PENB, PEGB2, +, PEGB6
			8'd5 : rdata = 44'b00001110111111101110000010000000000011100000;
			// PEs: 40 -> 
			// srcs: (24, 6)(451) 9 --> (451) 9:PENB, pass, 
			8'd6 : rdata = 44'b11000110111111100000000000000000000000000000;
			// PEs: 40, 41 -> 40
			// srcs: (30, 7)(646) 36, (451) 9 --> (647) 45:PENB, ALU, +, PEGB0
			8'd7 : rdata = 44'b00001110111111100011111111100000000010000000;
			// PEs: 40 -> 
			// srcs: (32, 8)(504) 5 --> (504) 5:PENB, pass, 
			8'd8 : rdata = 44'b11000110111111100000000000000000000000000000;
			// PEs: 40, 41 -> 40
			// srcs: (38, 9)(697) 64, (504) 5 --> (698) 69:PENB, ALU, +, PEGB0
			8'd9 : rdata = 44'b00001110111111100011111111100000000010000000;
			// PEs: 45, 40 -> 44
			// srcs: (39, 10)(731) 7, (536) 9 --> (732) 16:PEGB5, PENB, +, PEGB4
			8'd10 : rdata = 44'b00001111000010101101111111000000000011000000;
			// PEs: 40 -> 
			// srcs: (41, 11)(554) 14 --> (554) 14:PENB, pass, 
			8'd11 : rdata = 44'b11000110111111100000000000000000000000000000;
			// PEs: 40, 41 -> 40
			// srcs: (47, 12)(747) 67, (554) 14 --> (748) 81:PENB, ALU, +, PEGB0
			8'd12 : rdata = 44'b00001110111111100011111111100000000010000000;
			// PEs: 40 -> 
			// srcs: (49, 13)(614) 60 --> (614) 60:PENB, pass, 
			8'd13 : rdata = 44'b11000110111111100000000000000000000000000000;
			// PEs: 40, 41 -> 41
			// srcs: (55, 14)(612) 64, (614) 60 --> (615) 124:PENB, ALU, +, NI0
			8'd14 : rdata = 44'b00001110111111100011111111110000000000000000;
			// PEs: 40 -> 
			// srcs: (60, 15)(719) 30 --> (719) 30:PENB, pass, 
			8'd15 : rdata = 44'b11000110111111100000000000000000000000000000;
			// PEs: 40, 41 -> 41
			// srcs: (66, 16)(717) 53, (719) 30 --> (720) 83:PENB, ALU, +, NI1
			8'd16 : rdata = 44'b00001110111111100011111111110100000000000000;
			// PEs: 40, 41 -> 40
			// srcs: (67, 17)(610) 83, (615) 124 --> (616) 207:PENB, NI0, +, PEGB0
			8'd17 : rdata = 44'b00001110111111101010000000000000000010000000;
			// PEs: 41, 40 -> 
			// srcs: (91, 18)(720) 83, (725) 115 --> (726) 198:NI1, PENB, +, 
			8'd18 : rdata = 44'b00001101000000011101111111000000000000000000;
			// PEs: 40, 41 -> 
			// srcs: (104, 19)(715) 144, (726) 198 --> (727) 342:PENB, ALU, +, 
			8'd19 : rdata = 44'b00001110111111100011111111100000000000000000;
			// PEs: 41, 40 -> 40
			// srcs: (129, 20)(727) 342, (751) 724 --> (752) 1066:ALU, PENB, +, PEGB0
			8'd20 : rdata = 44'b00001001111111111101111111000000000010000000;
			// PEs: 40, 41 -> 42
			// srcs: (191, 21)(805) -9, (19) 0 --> (821) 0:PENB, ND2, *, PENB
			8'd21 : rdata = 44'b00011110111111100110000001000000000100000000;
			// PEs: 41, 42 -> 41
			// srcs: (200, 24)(220) 9, (1021) 0 --> (1221) 9:NW2, PEGB2, -, NW2
			8'd22 : rdata = 44'b00010010000000101110000010000010100000000000;
			// PEs: 40, 41 -> 42
			// srcs: (224, 22)(805) -9, (52) 6 --> (854) -54:PENB, ND0, *, PENB
			8'd23 : rdata = 44'b00011110111111100110000000000000000100000000;
			// PEs: 41, 42 -> 41
			// srcs: (233, 25)(253) 6, (1054) -54 --> (1254) 60:NW0, PEGB2, -, NW0
			8'd24 : rdata = 44'b00010010000000001110000010000010000000000000;
			// PEs: 40, 41 -> 42
			// srcs: (302, 23)(805) -9, (130) 6 --> (932) -54:PENB, ND1, *, PENB
			8'd25 : rdata = 44'b00011110111111100110000000100000000100000000;
			// PEs: 41, 42 -> 41
			// srcs: (311, 26)(331) 6, (1132) -54 --> (1332) 60:NW1, PEGB2, -, NW1
			8'd26 : rdata = 44'b00010010000000011110000010000010010000000000;
			default : rdata = 44'b00000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 42) begin
	always @(*) begin
		case(address)
			// PEs: 42, 42 -> 43
			// srcs: (1, 0)(54) 5, (255) 0 --> (455) 0:ND0, NW0, *, PENB
			8'd0 : rdata = 44'b00011011000000000100000000000000000100000000;
			// PEs: 42, 42 -> 43
			// srcs: (2, 1)(131) 9, (332) 4 --> (532) 36:ND1, NW1, *, PENB
			8'd1 : rdata = 44'b00011011000000010100000000100000000100000000;
			// PEs: 42, 42 -> 41
			// srcs: (3, 2)(22) 3, (223) 5 --> (423) 15:ND2, NW2, *, PEGB1
			8'd2 : rdata = 44'b00011011000000100100000001000000000010010000;
			// PEs: 45 -> 
			// srcs: (9, 3)(655) 0 --> (655) 0:PEGB5, pass, 
			8'd3 : rdata = 44'b11000111000010100000000000000000000000000000;
			// PEs: 43, 42 -> 40
			// srcs: (12, 4)(654) 12, (655) 0 --> (656) 12:PEGB3, ALU, +, PEGB0
			8'd4 : rdata = 44'b00001111000001100011111111100000000010000000;
			// PEs: 42, 41 -> 41
			// srcs: (194, 8)(3) 1, (821) 0 --> (1021) 0:NM0, PENB, *, PEGB1
			8'd5 : rdata = 44'b00011100000000001101111111000000000010010000;
			// PEs: 40, 42 -> 
			// srcs: (197, 5)(805) -9, (22) 3 --> (824) -27:PEGB0, ND2, *, 
			8'd6 : rdata = 44'b00011111000000000110000001000000000000000000;
			// PEs: 42, 42 -> 
			// srcs: (200, 9)(3) 1, (824) -27 --> (1024) -27:NM0, ALU, *, 
			8'd7 : rdata = 44'b00011100000000000011111111100000000000000000;
			// PEs: 42, 42 -> 42
			// srcs: (203, 12)(223) 5, (1024) -27 --> (1224) 32:NW2, ALU, -, NW2
			8'd8 : rdata = 44'b00010010000000100011111111100010100000000000;
			// PEs: 42, 41 -> 41
			// srcs: (227, 10)(3) 1, (854) -54 --> (1054) -54:NM0, PENB, *, PEGB1
			8'd9 : rdata = 44'b00011100000000001101111111000000000010010000;
			// PEs: 40, 42 -> 43
			// srcs: (229, 6)(805) -9, (54) 5 --> (856) -45:PEGB0, ND0, *, PENB
			8'd10 : rdata = 44'b00011111000000000110000000000000000100000000;
			// PEs: 42, 43 -> 42
			// srcs: (238, 13)(255) 0, (1056) -45 --> (1256) 45:NW0, PEGB3, -, NW0
			8'd11 : rdata = 44'b00010010000000001110000011000010000000000000;
			// PEs: 42, 41 -> 41
			// srcs: (305, 11)(3) 1, (932) -54 --> (1132) -54:NM0, PENB, *, PEGB1
			8'd12 : rdata = 44'b00011100000000001101111111000000000010010000;
			// PEs: 40, 42 -> 43
			// srcs: (306, 7)(805) -9, (131) 9 --> (933) -81:PEGB0, ND1, *, PENB
			8'd13 : rdata = 44'b00011111000000000110000000100000000100000000;
			// PEs: 42, 43 -> 42
			// srcs: (315, 14)(332) 4, (1133) -81 --> (1333) 85:NW1, PEGB3, -, NW1
			8'd14 : rdata = 44'b00010010000000011110000011000010010000000000;
			default : rdata = 44'b00000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 43) begin
	always @(*) begin
		case(address)
			// PEs: 43, 43 -> 43
			// srcs: (1, 0)(55) 6, (256) 2 --> (456) 12:ND0, NW0, *, NI0
			8'd0 : rdata = 44'b00011011000000000100000000010000000000000000;
			// PEs: 43, 43 -> 43
			// srcs: (2, 1)(132) 8, (333) 8 --> (533) 64:ND1, NW1, *, NI1
			8'd1 : rdata = 44'b00011011000000010100000000110100000000000000;
			// PEs: 43, 43 -> 40
			// srcs: (3, 2)(25) 4, (226) 0 --> (426) 0:ND2, NW2, *, PEGB0
			8'd2 : rdata = 44'b00011011000000100100000001000000000010000000;
			// PEs: 42, 43 -> 42
			// srcs: (4, 3)(455) 0, (456) 12 --> (654) 12:PENB, NI0, +, PEGB2
			8'd3 : rdata = 44'b00001110111111101010000000000000000010100000;
			// PEs: 42, 43 -> 44
			// srcs: (5, 4)(532) 36, (533) 64 --> (729) 100:PENB, NI1, +, PENB
			8'd4 : rdata = 44'b00001110111111101010000000100000000100000000;
			// PEs: 40, 43 -> 
			// srcs: (200, 5)(805) -9, (25) 4 --> (827) -36:PEGB0, ND2, *, 
			8'd5 : rdata = 44'b00011111000000000110000001000000000000000000;
			// PEs: 43, 43 -> 
			// srcs: (203, 8)(3) 1, (827) -36 --> (1027) -36:NM0, ALU, *, 
			8'd6 : rdata = 44'b00011100000000000011111111100000000000000000;
			// PEs: 43, 43 -> 43
			// srcs: (206, 11)(226) 0, (1027) -36 --> (1227) 36:NW2, ALU, -, NW2
			8'd7 : rdata = 44'b00010010000000100011111111100010100000000000;
			// PEs: 40, 43 -> 44
			// srcs: (230, 6)(805) -9, (55) 6 --> (857) -54:PEGB0, ND0, *, PENB
			8'd8 : rdata = 44'b00011111000000000110000000000000000100000000;
			// PEs: 43, 42 -> 42
			// srcs: (232, 9)(3) 1, (856) -45 --> (1056) -45:NM0, PENB, *, PEGB2
			8'd9 : rdata = 44'b00011100000000001101111111000000000010100000;
			// PEs: 43, 44 -> 43
			// srcs: (239, 12)(256) 2, (1057) -54 --> (1257) 56:NW0, PEGB4, -, NW0
			8'd10 : rdata = 44'b00010010000000001110000100000010000000000000;
			// PEs: 40, 43 -> 44
			// srcs: (307, 7)(805) -9, (132) 8 --> (934) -72:PEGB0, ND1, *, PENB
			8'd11 : rdata = 44'b00011111000000000110000000100000000100000000;
			// PEs: 43, 42 -> 42
			// srcs: (309, 10)(3) 1, (933) -81 --> (1133) -81:NM0, PENB, *, PEGB2
			8'd12 : rdata = 44'b00011100000000001101111111000000000010100000;
			// PEs: 43, 44 -> 43
			// srcs: (316, 13)(333) 8, (1134) -72 --> (1334) 80:NW1, PEGB4, -, NW1
			8'd13 : rdata = 44'b00010010000000011110000100000010010000000000;
			default : rdata = 44'b00000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 44) begin
	always @(*) begin
		case(address)
			// PEs: 44, 44 -> 45
			// srcs: (1, 0)(56) 0, (257) 6 --> (457) 0:ND0, NW0, *, PENB
			8'd0 : rdata = 44'b00011011000000000100000000000000000100000000;
			// PEs: 44, 44 -> 45
			// srcs: (2, 1)(133) 7, (334) 1 --> (534) 7:ND1, NW1, *, PENB
			8'd1 : rdata = 44'b00011011000000010100000000100000000100000000;
			// PEs: 44, 44 -> 40
			// srcs: (3, 2)(28) 1, (229) 4 --> (429) 4:ND2, NW2, *, PEGB0
			8'd2 : rdata = 44'b00011011000000100100000001000000000010000000;
			// PEs: 41, 43 -> 
			// srcs: (15, 3)(728) 54, (729) 100 --> (730) 154:PEGB1, PENB, +, 
			8'd3 : rdata = 44'b00001111000000101101111111000000000000000000;
			// PEs: 44, 41 -> 40
			// srcs: (45, 4)(730) 154, (732) 16 --> (733) 170:ALU, PEGB1, +, PEGB0
			8'd4 : rdata = 44'b00001001111111111110000001000000000010000000;
			// PEs: 40, 44 -> 
			// srcs: (203, 5)(805) -9, (28) 1 --> (830) -9:PEGB0, ND2, *, 
			8'd5 : rdata = 44'b00011111000000000110000001000000000000000000;
			// PEs: 44, 44 -> 
			// srcs: (206, 8)(3) 1, (830) -9 --> (1030) -9:NM0, ALU, *, 
			8'd6 : rdata = 44'b00011100000000000011111111100000000000000000;
			// PEs: 44, 44 -> 44
			// srcs: (209, 11)(229) 4, (1030) -9 --> (1230) 13:NW2, ALU, -, NW2
			8'd7 : rdata = 44'b00010010000000100011111111100010100000000000;
			// PEs: 40, 44 -> 45
			// srcs: (231, 6)(805) -9, (56) 0 --> (858) 0:PEGB0, ND0, *, PENB
			8'd8 : rdata = 44'b00011111000000000110000000000000000100000000;
			// PEs: 44, 43 -> 43
			// srcs: (233, 9)(3) 1, (857) -54 --> (1057) -54:NM0, PENB, *, PEGB3
			8'd9 : rdata = 44'b00011100000000001101111111000000000010110000;
			// PEs: 44, 45 -> 44
			// srcs: (240, 12)(257) 6, (1058) 0 --> (1258) 6:NW0, PEGB5, -, NW0
			8'd10 : rdata = 44'b00010010000000001110000101000010000000000000;
			// PEs: 40, 44 -> 45
			// srcs: (308, 7)(805) -9, (133) 7 --> (935) -63:PEGB0, ND1, *, PENB
			8'd11 : rdata = 44'b00011111000000000110000000100000000100000000;
			// PEs: 44, 43 -> 43
			// srcs: (310, 10)(3) 1, (934) -72 --> (1134) -72:NM0, PENB, *, PEGB3
			8'd12 : rdata = 44'b00011100000000001101111111000000000010110000;
			// PEs: 44, 45 -> 44
			// srcs: (317, 13)(334) 1, (1135) -63 --> (1335) 64:NW1, PEGB5, -, NW1
			8'd13 : rdata = 44'b00010010000000011110000101000010010000000000;
			default : rdata = 44'b00000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 45) begin
	always @(*) begin
		case(address)
			// PEs: 45, 45 -> 45
			// srcs: (1, 0)(57) 6, (258) 0 --> (458) 0:ND0, NW0, *, NI0
			8'd0 : rdata = 44'b00011011000000000100000000010000000000000000;
			// PEs: 45, 45 -> 45
			// srcs: (2, 1)(134) 3, (335) 0 --> (535) 0:ND1, NW1, *, NI1
			8'd1 : rdata = 44'b00011011000000010100000000110100000000000000;
			// PEs: 45, 45 -> 40
			// srcs: (3, 2)(35) 9, (236) 1 --> (436) 9:ND2, NW2, *, PEGB0
			8'd2 : rdata = 44'b00011011000000100100000001000000000010000000;
			// PEs: 44, 45 -> 42
			// srcs: (4, 4)(457) 0, (458) 0 --> (655) 0:PENB, NI0, +, PEGB2
			8'd3 : rdata = 44'b00001110111111101010000000000000000010100000;
			// PEs: 44, 45 -> 41
			// srcs: (5, 3)(534) 7, (535) 0 --> (731) 7:PENB, NI1, +, PEGB1
			8'd4 : rdata = 44'b00001110111111101010000000100000000010010000;
			// PEs: 40, 45 -> 
			// srcs: (210, 5)(805) -9, (35) 9 --> (837) -81:PEGB0, ND2, *, 
			8'd5 : rdata = 44'b00011111000000000110000001000000000000000000;
			// PEs: 45, 45 -> 
			// srcs: (213, 8)(3) 1, (837) -81 --> (1037) -81:NM0, ALU, *, 
			8'd6 : rdata = 44'b00011100000000000011111111100000000000000000;
			// PEs: 45, 45 -> 45
			// srcs: (216, 11)(236) 1, (1037) -81 --> (1237) 82:NW2, ALU, -, NW2
			8'd7 : rdata = 44'b00010010000000100011111111100010100000000000;
			// PEs: 40, 45 -> 46
			// srcs: (232, 6)(805) -9, (57) 6 --> (859) -54:PEGB0, ND0, *, PENB
			8'd8 : rdata = 44'b00011111000000000110000000000000000100000000;
			// PEs: 45, 44 -> 44
			// srcs: (234, 9)(3) 1, (858) 0 --> (1058) 0:NM0, PENB, *, PEGB4
			8'd9 : rdata = 44'b00011100000000001101111111000000000011000000;
			// PEs: 45, 46 -> 45
			// srcs: (241, 12)(258) 0, (1059) -54 --> (1259) 54:NW0, PEGB6, -, NW0
			8'd10 : rdata = 44'b00010010000000001110000110000010000000000000;
			// PEs: 40, 45 -> 46
			// srcs: (309, 7)(805) -9, (134) 3 --> (936) -27:PEGB0, ND1, *, PENB
			8'd11 : rdata = 44'b00011111000000000110000000100000000100000000;
			// PEs: 45, 44 -> 44
			// srcs: (311, 10)(3) 1, (935) -63 --> (1135) -63:NM0, PENB, *, PEGB4
			8'd12 : rdata = 44'b00011100000000001101111111000000000011000000;
			// PEs: 45, 46 -> 45
			// srcs: (318, 13)(335) 0, (1136) -27 --> (1336) 27:NW1, PEGB6, -, NW1
			8'd13 : rdata = 44'b00010010000000011110000110000010010000000000;
			default : rdata = 44'b00000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 46) begin
	always @(*) begin
		case(address)
			// PEs: 46, 46 -> 47
			// srcs: (1, 0)(58) 2, (259) 5 --> (459) 10:ND0, NW0, *, PENB
			8'd0 : rdata = 44'b00011011000000000100000000000000000100000000;
			// PEs: 46, 46 -> 47
			// srcs: (2, 1)(136) 2, (337) 5 --> (537) 10:ND1, NW1, *, PENB
			8'd1 : rdata = 44'b00011011000000010100000000100000000100000000;
			// PEs: 46, 46 -> 40
			// srcs: (3, 2)(38) 9, (239) 2 --> (439) 18:ND2, NW2, *, PEGB0
			8'd2 : rdata = 44'b00011011000000100100000001000000000010000000;
			// PEs: 40 -> 
			// srcs: (53, 3)(618) 112 --> (618) 112:PEGB0, pass, 
			8'd3 : rdata = 44'b11000111000000000000000000000000000000000000;
			// PEs: 46, 41 -> 40
			// srcs: (55, 4)(618) 112, (620) 106 --> (621) 218:ALU, PEGB1, +, PEGB0
			8'd4 : rdata = 44'b00001001111111111110000001000000000010000000;
			// PEs: 40, 46 -> 
			// srcs: (213, 5)(805) -9, (38) 9 --> (840) -81:PEGB0, ND2, *, 
			8'd5 : rdata = 44'b00011111000000000110000001000000000000000000;
			// PEs: 46, 46 -> 
			// srcs: (216, 8)(3) 1, (840) -81 --> (1040) -81:NM0, ALU, *, 
			8'd6 : rdata = 44'b00011100000000000011111111100000000000000000;
			// PEs: 46, 46 -> 46
			// srcs: (219, 12)(239) 2, (1040) -81 --> (1240) 83:NW2, ALU, -, NW2
			8'd7 : rdata = 44'b00010010000000100011111111100010100000000000;
			// PEs: 40, 46 -> 47
			// srcs: (233, 6)(805) -9, (58) 2 --> (860) -18:PEGB0, ND0, *, PENB
			8'd8 : rdata = 44'b00011111000000000110000000000000000100000000;
			// PEs: 46, 45 -> 45
			// srcs: (235, 9)(3) 1, (859) -54 --> (1059) -54:NM0, PENB, *, PEGB5
			8'd9 : rdata = 44'b00011100000000001101111111000000000011010000;
			// PEs: 46, 47 -> 46
			// srcs: (242, 13)(259) 5, (1060) -18 --> (1260) 23:NW0, PEGB7, -, NW0
			8'd10 : rdata = 44'b00010010000000001110000111000010000000000000;
			// PEs: 40, 46 -> 46
			// srcs: (311, 7)(805) -9, (136) 2 --> (938) -18:PEGB0, ND1, *, NI0
			8'd11 : rdata = 44'b00011111000000000110000000110000000000000000;
			// PEs: 46, 45 -> 45
			// srcs: (312, 10)(3) 1, (936) -27 --> (1136) -27:NM0, PENB, *, PEGB5
			8'd12 : rdata = 44'b00011100000000001101111111000000000011010000;
			// PEs: 46, 46 -> 
			// srcs: (314, 11)(3) 1, (938) -18 --> (1138) -18:NM0, NI0, *, 
			8'd13 : rdata = 44'b00011100000000001010000000000000000000000000;
			// PEs: 46, 46 -> 46
			// srcs: (317, 14)(337) 5, (1138) -18 --> (1338) 23:NW1, ALU, -, NW1
			8'd14 : rdata = 44'b00010010000000010011111111100010010000000000;
			default : rdata = 44'b00000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 47) begin
	always @(*) begin
		case(address)
			// PEs: 47, 47 -> 47
			// srcs: (1, 0)(59) 9, (260) 4 --> (460) 36:ND0, NW0, *, NI0
			8'd0 : rdata = 44'b00011011000000000100000000010000000000000000;
			// PEs: 47, 47 -> 47
			// srcs: (2, 1)(137) 9, (338) 5 --> (538) 45:ND1, NW1, *, NI1
			8'd1 : rdata = 44'b00011011000000010100000000110100000000000000;
			// PEs: 47, 47 -> 40
			// srcs: (3, 2)(41) 0, (242) 4 --> (442) 0:ND2, NW2, *, PENB
			8'd2 : rdata = 44'b00011011000000100100000001000000000100000000;
			// PEs: 46, 47 -> 40
			// srcs: (4, 3)(459) 10, (460) 36 --> (657) 46:PENB, NI0, +, PENB
			8'd3 : rdata = 44'b00001110111111101010000000000000000100000000;
			// PEs: 46, 47 -> 40
			// srcs: (5, 4)(537) 10, (538) 45 --> (734) 55:PENB, NI1, +, PENB
			8'd4 : rdata = 44'b00001110111111101010000000100000000100000000;
			// PEs: 40, 47 -> 
			// srcs: (216, 5)(805) -9, (41) 0 --> (843) 0:PEGB0, ND2, *, 
			8'd5 : rdata = 44'b00011111000000000110000001000000000000000000;
			// PEs: 47, 47 -> 
			// srcs: (219, 8)(3) 1, (843) 0 --> (1043) 0:NM0, ALU, *, 
			8'd6 : rdata = 44'b00011100000000000011111111100000000000000000;
			// PEs: 47, 47 -> 47
			// srcs: (222, 12)(242) 4, (1043) 0 --> (1243) 4:NW2, ALU, -, NW2
			8'd7 : rdata = 44'b00010010000000100011111111100010100000000000;
			// PEs: 40, 47 -> 47
			// srcs: (234, 6)(805) -9, (59) 9 --> (861) -81:PEGB0, ND0, *, NI0
			8'd8 : rdata = 44'b00011111000000000110000000010000000000000000;
			// PEs: 47, 46 -> 46
			// srcs: (236, 9)(3) 1, (860) -18 --> (1060) -18:NM0, PENB, *, PEGB6
			8'd9 : rdata = 44'b00011100000000001101111111000000000011100000;
			// PEs: 47, 47 -> 
			// srcs: (237, 10)(3) 1, (861) -81 --> (1061) -81:NM0, NI0, *, 
			8'd10 : rdata = 44'b00011100000000001010000000000000000000000000;
			// PEs: 47, 47 -> 47
			// srcs: (240, 13)(260) 4, (1061) -81 --> (1261) 85:NW0, ALU, -, NW0
			8'd11 : rdata = 44'b00010010000000000011111111100010000000000000;
			// PEs: 40, 47 -> 
			// srcs: (312, 7)(805) -9, (137) 9 --> (939) -81:PEGB0, ND1, *, 
			8'd12 : rdata = 44'b00011111000000000110000000100000000000000000;
			// PEs: 47, 47 -> 
			// srcs: (315, 11)(3) 1, (939) -81 --> (1139) -81:NM0, ALU, *, 
			8'd13 : rdata = 44'b00011100000000000011111111100000000000000000;
			// PEs: 47, 47 -> 47
			// srcs: (318, 14)(338) 5, (1139) -81 --> (1339) 86:NW1, ALU, -, NW1
			8'd14 : rdata = 44'b00010010000000010011111111100010010000000000;
			default : rdata = 44'b00000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 48) begin
	always @(*) begin
		case(address)
			// PEs: 55 -> 56
			// srcs: (3, 0)(471) 8 --> (471) 8:PENB, pass, PUNB
			8'd0 : rdata = 44'b11000110111111100000000000000000001000000000;
			// PEs: 55 -> 56
			// srcs: (4, 1)(549) 48 --> (549) 48:PENB, pass, PUNB
			8'd1 : rdata = 44'b11000110111111100000000000000000001000000000;
			// PEs: 49 -> 16
			// srcs: (8, 8)(445) 30 --> (445) 30:PEGB1, pass, PUGB2
			8'd2 : rdata = 44'b11000111000000100000000000000000000000001010;
			// PEs: 51 -> 40
			// srcs: (9, 10)(451) 9 --> (451) 9:PEGB3, pass, PUGB5
			8'd3 : rdata = 44'b11000111000001100000000000000000000000001101;
			// PEs: 54 -> 56
			// srcs: (10, 13)(666) 48 --> (666) 48:PEGB6, pass, PUNB
			8'd4 : rdata = 44'b11000111000011000000000000000000001000000000;
			// PEs: 52 -> 56
			// srcs: (11, 15)(740) 24 --> (740) 24:PEGB4, pass, PUNB
			8'd5 : rdata = 44'b11000111000010000000000000000000001000000000;
			// PEs: 54 -> 32
			// srcs: (12, 16)(742) 32 --> (742) 32:PEGB6, pass, PUGB4
			8'd6 : rdata = 44'b11000111000011000000000000000000000000001100;
			// PEs: 32 -> 48
			// srcs: (13, 3)(411) 9 --> (411) 9:PUGB4, pass, NI0
			8'd7 : rdata = 44'b11000111000010010000000000010000000000000000;
			// PEs: 0 -> 49
			// srcs: (19, 2)(608) 0 --> (608) 0:PUGB0, pass, PENB
			8'd8 : rdata = 44'b11000111000000010000000000000000000100000000;
			// PEs: 0 -> 55
			// srcs: (22, 20)(607) 74 --> (607) 74:PUGB0, pass, PEGB7
			8'd9 : rdata = 44'b11000111000000010000000000000000000011110000;
			// PEs: 48 -> 49
			// srcs: (26, 4)(411) 9 --> (411) 9:NI0, pass, PENB
			8'd10 : rdata = 44'b11000101000000000000000000000000000100000000;
			// PEs: 16 -> 48
			// srcs: (27, 5)(622) 46 --> (622) 46:PUGB2, pass, NI0
			8'd11 : rdata = 44'b11000111000001010000000000010000000000000000;
			// PEs: 40 -> 49
			// srcs: (28, 6)(426) 0 --> (426) 0:PUNB, pass, PENB
			8'd12 : rdata = 44'b11000110111111110000000000000000000100000000;
			// PEs: 48 -> 49
			// srcs: (34, 7)(622) 46 --> (622) 46:NI0, pass, PENB
			8'd13 : rdata = 44'b11000101000000000000000000000000000100000000;
			// PEs: 32 -> 49
			// srcs: (35, 9)(643) 63 --> (643) 63:PUGB4, pass, PENB
			8'd14 : rdata = 44'b11000111000010010000000000000000000100000000;
			// PEs: 40 -> 49
			// srcs: (36, 11)(648) 36 --> (648) 36:PUNB, pass, PENB
			8'd15 : rdata = 44'b11000110111111110000000000000000000100000000;
			// PEs: 40 -> 49
			// srcs: (37, 12)(657) 46 --> (657) 46:PUNB, pass, PENB
			8'd16 : rdata = 44'b11000110111111110000000000000000000100000000;
			// PEs: 8 -> 49
			// srcs: (38, 14)(542) 72 --> (542) 72:PUGB1, pass, PENB
			8'd17 : rdata = 44'b11000111000000110000000000000000000100000000;
			// PEs: 56 -> 48
			// srcs: (39, 17)(745) 93 --> (745) 93:PUGB7, pass, NI0
			8'd18 : rdata = 44'b11000111000011110000000000010000000000000000;
			// PEs: 49 -> 56
			// srcs: (41, 21)(623) 46 --> (623) 46:PEGB1, pass, PUNB
			8'd19 : rdata = 44'b11000111000000100000000000000000001000000000;
			// PEs: 49 -> 0
			// srcs: (42, 25)(644) 99 --> (644) 99:PEGB1, pass, PUGB0
			8'd20 : rdata = 44'b11000111000000100000000000000000000000001000;
			// PEs: 16 -> 49
			// srcs: (43, 18)(551) 21 --> (551) 21:PUGB2, pass, PENB
			8'd21 : rdata = 44'b11000111000001010000000000000000000100000000;
			// PEs: 49 -> 16
			// srcs: (45, 28)(737) 149 --> (737) 149:PEGB1, pass, PUGB2
			8'd22 : rdata = 44'b11000111000000100000000000000000000000001010;
			// PEs: 55 -> 40
			// srcs: (46, 30)(610) 83 --> (610) 83:PENB, pass, PUGB5
			8'd23 : rdata = 44'b11000110111111100000000000000000000000001101;
			// PEs: 48 -> 49
			// srcs: (49, 19)(745) 93 --> (745) 93:NI0, pass, PENB
			8'd24 : rdata = 44'b11000101000000000000000000000000000100000000;
			// PEs: 24 -> 48
			// srcs: (50, 22)(631) 99 --> (631) 99:PUGB3, pass, NI0
			8'd25 : rdata = 44'b11000111000001110000000000010000000000000000;
			// PEs: 0 -> 49
			// srcs: (51, 23)(633) 84 --> (633) 84:PUGB0, pass, PENB
			8'd26 : rdata = 44'b11000111000000010000000000000000000100000000;
			// PEs: 48 -> 49
			// srcs: (57, 24)(631) 99 --> (631) 99:NI0, pass, PENB
			8'd27 : rdata = 44'b11000101000000000000000000000000000100000000;
			// PEs: 40 -> 49
			// srcs: (58, 26)(647) 45 --> (647) 45:PUNB, pass, PENB
			8'd28 : rdata = 44'b11000110111111110000000000000000000100000000;
			// PEs: 40 -> 49
			// srcs: (59, 27)(656) 12 --> (656) 12:PUNB, pass, PENB
			8'd29 : rdata = 44'b11000110111111110000000000000000000100000000;
			// PEs: 40 -> 53
			// srcs: (60, 29)(748) 81 --> (748) 81:PUNB, pass, PEGB5
			8'd30 : rdata = 44'b11000110111111110000000000000000000011010000;
			// PEs: 49 -> 8
			// srcs: (64, 31)(634) 183 --> (634) 183:PEGB1, pass, PUGB1
			8'd31 : rdata = 44'b11000111000000100000000000000000000000001001;
			// PEs: 0 -> 49
			// srcs: (67, 32)(645) 180 --> (645) 180:PUGB0, pass, PENB
			8'd32 : rdata = 44'b11000111000000010000000000000000000100000000;
			// PEs: 40 -> 48
			// srcs: (68, 33)(733) 170 --> (733) 170:PUNB, pass, NI0
			8'd33 : rdata = 44'b11000110111111110000000000010000000000000000;
			// PEs: 53 -> 56
			// srcs: (72, 36)(749) 195 --> (749) 195:PEGB5, pass, PUNB
			8'd34 : rdata = 44'b11000111000010100000000000000000001000000000;
			// PEs: 50 -> 56
			// srcs: (73, 38)(665) 184 --> (665) 184:PEGB2, pass, PUNB
			8'd35 : rdata = 44'b11000111000001000000000000000000001000000000;
			// PEs: 16 -> 49
			// srcs: (75, 34)(738) 267 --> (738) 267:PUGB2, pass, PENB
			8'd36 : rdata = 44'b11000111000001010000000000000000000100000000;
			// PEs: 49 -> 16
			// srcs: (78, 37)(651) 315 --> (651) 315:PEGB1, pass, PUGB2
			8'd37 : rdata = 44'b11000111000000100000000000000000000000001010;
			// PEs: 48 -> 49
			// srcs: (82, 35)(733) 170 --> (733) 170:NI0, pass, PENB
			8'd38 : rdata = 44'b11000101000000000000000000000000000100000000;
			// PEs: 49 -> 56
			// srcs: (89, 39)(739) 437 --> (739) 437:PEGB1, pass, PUNB
			8'd39 : rdata = 44'b11000111000000100000000000000000001000000000;
			// PEs: 0 -> 48
			// srcs: (119, 40)(776) 448 --> (776) 448:PUGB0, pass, NI0
			8'd40 : rdata = 44'b11000111000000010000000000010000000000000000;
			// PEs: 32 -> 49
			// srcs: (120, 41)(800) 542 --> (800) 542:PUGB4, pass, PENB
			8'd41 : rdata = 44'b11000111000010010000000000000000000100000000;
			// PEs: 48 -> 49
			// srcs: (127, 42)(776) 448 --> (776) 448:NI0, pass, PENB
			8'd42 : rdata = 44'b11000101000000000000000000000000000100000000;
			// PEs: 40 -> 49
			// srcs: (136, 43)(752) 1066 --> (752) 1066:PUNB, pass, PENB
			8'd43 : rdata = 44'b11000110111111110000000000000000000100000000;
			// PEs: 49 -> 0
			// srcs: (144, 44)(802) 2056 --> (802) 2056:PEGB1, pass, PUGB0
			8'd44 : rdata = 44'b11000111000000100000000000000000000000001000;
			// PEs: 0 -> 49
			// srcs: (214, 45)(805) -9 --> (805) -9:PUGB0, pass, PENB
			8'd45 : rdata = 44'b11000111000000010000000000000000000100000000;
			// PEs: 0 -> 50
			// srcs: (217, 46)(805) -9 --> (805) -9:PUGB0, pass, PEGB2
			8'd46 : rdata = 44'b11000111000000010000000000000000000010100000;
			// PEs: 0 -> 51
			// srcs: (220, 47)(805) -9 --> (805) -9:PUGB0, pass, PEGB3
			8'd47 : rdata = 44'b11000111000000010000000000000000000010110000;
			// PEs: 0 -> 52
			// srcs: (223, 48)(805) -9 --> (805) -9:PUGB0, pass, PEGB4
			8'd48 : rdata = 44'b11000111000000010000000000000000000011000000;
			// PEs: 0 -> 53
			// srcs: (230, 49)(805) -9 --> (805) -9:PUGB0, pass, PEGB5
			8'd49 : rdata = 44'b11000111000000010000000000000000000011010000;
			// PEs: 0 -> 49
			// srcs: (231, 50)(805) -9 --> (805) -9:PUGB0, pass, PENB
			8'd50 : rdata = 44'b11000111000000010000000000000000000100000000;
			// PEs: 0 -> 50
			// srcs: (232, 51)(805) -9 --> (805) -9:PUGB0, pass, PEGB2
			8'd51 : rdata = 44'b11000111000000010000000000000000000010100000;
			// PEs: 0 -> 54
			// srcs: (233, 52)(805) -9 --> (805) -9:PUGB0, pass, PEGB6
			8'd52 : rdata = 44'b11000111000000010000000000000000000011100000;
			// PEs: 0 -> 51
			// srcs: (234, 53)(805) -9 --> (805) -9:PUGB0, pass, PEGB3
			8'd53 : rdata = 44'b11000111000000010000000000000000000010110000;
			// PEs: 0 -> 52
			// srcs: (235, 54)(805) -9 --> (805) -9:PUGB0, pass, PEGB4
			8'd54 : rdata = 44'b11000111000000010000000000000000000011000000;
			// PEs: 0 -> 55
			// srcs: (236, 55)(805) -9 --> (805) -9:PUGB0, pass, PEGB7
			8'd55 : rdata = 44'b11000111000000010000000000000000000011110000;
			// PEs: 0 -> 53
			// srcs: (237, 56)(805) -9 --> (805) -9:PUGB0, pass, PEGB5
			8'd56 : rdata = 44'b11000111000000010000000000000000000011010000;
			// PEs: 0 -> 54
			// srcs: (238, 57)(805) -9 --> (805) -9:PUGB0, pass, PEGB6
			8'd57 : rdata = 44'b11000111000000010000000000000000000011100000;
			// PEs: 0 -> 55
			// srcs: (240, 58)(805) -9 --> (805) -9:PUGB0, pass, PEGB7
			8'd58 : rdata = 44'b11000111000000010000000000000000000011110000;
			// PEs: 0 -> 49
			// srcs: (309, 59)(805) -9 --> (805) -9:PUGB0, pass, PENB
			8'd59 : rdata = 44'b11000111000000010000000000000000000100000000;
			// PEs: 0 -> 50
			// srcs: (310, 60)(805) -9 --> (805) -9:PUGB0, pass, PEGB2
			8'd60 : rdata = 44'b11000111000000010000000000000000000010100000;
			// PEs: 0 -> 51
			// srcs: (312, 61)(805) -9 --> (805) -9:PUGB0, pass, PEGB3
			8'd61 : rdata = 44'b11000111000000010000000000000000000010110000;
			// PEs: 0 -> 52
			// srcs: (313, 62)(805) -9 --> (805) -9:PUGB0, pass, PEGB4
			8'd62 : rdata = 44'b11000111000000010000000000000000000011000000;
			// PEs: 0 -> 53
			// srcs: (315, 63)(805) -9 --> (805) -9:PUGB0, pass, PEGB5
			8'd63 : rdata = 44'b11000111000000010000000000000000000011010000;
			// PEs: 0 -> 54
			// srcs: (316, 64)(805) -9 --> (805) -9:PUGB0, pass, PEGB6
			8'd64 : rdata = 44'b11000111000000010000000000000000000011100000;
			// PEs: 0 -> 55
			// srcs: (318, 65)(805) -9 --> (805) -9:PUGB0, pass, PEGB7
			8'd65 : rdata = 44'b11000111000000010000000000000000000011110000;
			default : rdata = 44'b00000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 49) begin
	always @(*) begin
		case(address)
			// PEs: 49, 49 -> 50
			// srcs: (1, 0)(61) 9, (262) 0 --> (462) 0:ND0, NW0, *, PENB
			8'd0 : rdata = 44'b00011011000000000100000000000000000100000000;
			// PEs: 49, 49 -> 50
			// srcs: (2, 1)(139) 5, (340) 7 --> (540) 35:ND1, NW1, *, PENB
			8'd1 : rdata = 44'b00011011000000010100000000100000000100000000;
			// PEs: 49, 49 -> 48
			// srcs: (3, 2)(44) 6, (245) 5 --> (445) 30:ND2, NW2, *, PEGB0
			8'd2 : rdata = 44'b00011011000000100100000001000000000010000000;
			// PEs: 48 -> 
			// srcs: (21, 3)(608) 0 --> (608) 0:PENB, pass, 
			8'd3 : rdata = 44'b11000110111111100000000000000000000000000000;
			// PEs: 49, 48 -> 55
			// srcs: (28, 4)(608) 0, (411) 9 --> (609) 9:ALU, PENB, +, PEGB7
			8'd4 : rdata = 44'b00001001111111111101111111000000000011110000;
			// PEs: 48 -> 
			// srcs: (30, 5)(426) 0 --> (426) 0:PENB, pass, 
			8'd5 : rdata = 44'b11000110111111100000000000000000000000000000;
			// PEs: 48, 49 -> 48
			// srcs: (36, 6)(622) 46, (426) 0 --> (623) 46:PENB, ALU, +, PEGB0
			8'd6 : rdata = 44'b00001110111111100011111111100000000010000000;
			// PEs: 48, 50 -> 48
			// srcs: (37, 7)(643) 63, (448) 36 --> (644) 99:PENB, PEGB2, +, PEGB0
			8'd7 : rdata = 44'b00001110111111101110000010000000000010000000;
			// PEs: 48, 52 -> 49
			// srcs: (38, 8)(648) 36, (454) 54 --> (649) 90:PENB, PEGB4, +, NI0
			8'd8 : rdata = 44'b00001110111111101110000100010000000000000000;
			// PEs: 48, 53 -> 49
			// srcs: (39, 9)(657) 46, (461) 6 --> (658) 52:PENB, PEGB5, +, NI1
			8'd9 : rdata = 44'b00001110111111101110000101010100000000000000;
			// PEs: 50, 48 -> 48
			// srcs: (40, 10)(736) 77, (542) 72 --> (737) 149:PEGB2, PENB, +, PEGB0
			8'd10 : rdata = 44'b00001111000001001101111111000000000010000000;
			// PEs: 48 -> 
			// srcs: (45, 11)(551) 21 --> (551) 21:PENB, pass, 
			8'd11 : rdata = 44'b11000110111111100000000000000000000000000000;
			// PEs: 48, 49 -> 53
			// srcs: (51, 12)(745) 93, (551) 21 --> (746) 114:PENB, ALU, +, PEGB5
			8'd12 : rdata = 44'b00001110111111100011111111100000000011010000;
			// PEs: 48 -> 
			// srcs: (53, 13)(633) 84 --> (633) 84:PENB, pass, 
			8'd13 : rdata = 44'b11000110111111100000000000000000000000000000;
			// PEs: 48, 49 -> 48
			// srcs: (59, 14)(631) 99, (633) 84 --> (634) 183:PENB, ALU, +, PEGB0
			8'd14 : rdata = 44'b00001110111111100011111111100000000010000000;
			// PEs: 48, 49 -> 49
			// srcs: (60, 15)(647) 45, (649) 90 --> (650) 135:PENB, NI0, +, NI2
			8'd15 : rdata = 44'b00001110111111101010000000011000000000000000;
			// PEs: 48, 49 -> 50
			// srcs: (61, 16)(656) 12, (658) 52 --> (659) 64:PENB, NI1, +, PENB
			8'd16 : rdata = 44'b00001110111111101010000000100000000100000000;
			// PEs: 48, 49 -> 48
			// srcs: (73, 17)(645) 180, (650) 135 --> (651) 315:PENB, NI2, +, PEGB0
			8'd17 : rdata = 44'b00001110111111101010000001000000000010000000;
			// PEs: 48 -> 
			// srcs: (77, 18)(738) 267 --> (738) 267:PENB, pass, 
			8'd18 : rdata = 44'b11000110111111100000000000000000000000000000;
			// PEs: 48, 49 -> 48
			// srcs: (84, 19)(733) 170, (738) 267 --> (739) 437:PENB, ALU, +, PEGB0
			8'd19 : rdata = 44'b00001110111111100011111111100000000010000000;
			// PEs: 48 -> 
			// srcs: (122, 20)(800) 542 --> (800) 542:PENB, pass, 
			8'd20 : rdata = 44'b11000110111111100000000000000000000000000000;
			// PEs: 48, 49 -> 
			// srcs: (129, 21)(776) 448, (800) 542 --> (801) 990:PENB, ALU, +, 
			8'd21 : rdata = 44'b00001110111111100011111111100000000000000000;
			// PEs: 48, 49 -> 48
			// srcs: (139, 22)(752) 1066, (801) 990 --> (802) 2056:PENB, ALU, +, PEGB0
			8'd22 : rdata = 44'b00001110111111100011111111100000000010000000;
			// PEs: 48, 49 -> 50
			// srcs: (216, 23)(805) -9, (44) 6 --> (846) -54:PENB, ND2, *, PENB
			8'd23 : rdata = 44'b00011110111111100110000001000000000100000000;
			// PEs: 49, 50 -> 49
			// srcs: (225, 26)(245) 5, (1046) -54 --> (1246) 59:NW2, PEGB2, -, NW2
			8'd24 : rdata = 44'b00010010000000101110000010000010100000000000;
			// PEs: 48, 49 -> 50
			// srcs: (233, 24)(805) -9, (61) 9 --> (863) -81:PENB, ND0, *, PENB
			8'd25 : rdata = 44'b00011110111111100110000000000000000100000000;
			// PEs: 49, 50 -> 49
			// srcs: (242, 27)(262) 0, (1063) -81 --> (1263) 81:NW0, PEGB2, -, NW0
			8'd26 : rdata = 44'b00010010000000001110000010000010000000000000;
			// PEs: 48, 49 -> 50
			// srcs: (311, 25)(805) -9, (139) 5 --> (941) -45:PENB, ND1, *, PENB
			8'd27 : rdata = 44'b00011110111111100110000000100000000100000000;
			// PEs: 49, 50 -> 49
			// srcs: (320, 28)(340) 7, (1141) -45 --> (1341) 52:NW1, PEGB2, -, NW1
			8'd28 : rdata = 44'b00010010000000011110000010000010010000000000;
			default : rdata = 44'b00000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 50) begin
	always @(*) begin
		case(address)
			// PEs: 50, 50 -> 50
			// srcs: (1, 0)(62) 8, (263) 5 --> (463) 40:ND0, NW0, *, NI0
			8'd0 : rdata = 44'b00011011000000000100000000010000000000000000;
			// PEs: 50, 50 -> 50
			// srcs: (2, 1)(140) 6, (341) 7 --> (541) 42:ND1, NW1, *, NI1
			8'd1 : rdata = 44'b00011011000000010100000000110100000000000000;
			// PEs: 50, 50 -> 49
			// srcs: (3, 2)(47) 4, (248) 9 --> (448) 36:ND2, NW2, *, PEGB1
			8'd2 : rdata = 44'b00011011000000100100000001000000000010010000;
			// PEs: 49, 50 -> 51
			// srcs: (4, 3)(462) 0, (463) 40 --> (660) 40:PENB, NI0, +, PENB
			8'd3 : rdata = 44'b00001110111111101010000000000000000100000000;
			// PEs: 49, 50 -> 49
			// srcs: (5, 4)(540) 35, (541) 42 --> (736) 77:PENB, NI1, +, PEGB1
			8'd4 : rdata = 44'b00001110111111101010000000100000000010010000;
			// PEs: 49, 51 -> 48
			// srcs: (67, 5)(659) 64, (664) 120 --> (665) 184:PENB, PEGB3, +, PEGB0
			8'd5 : rdata = 44'b00001110111111101110000011000000000010000000;
			// PEs: 50, 49 -> 49
			// srcs: (219, 9)(3) 1, (846) -54 --> (1046) -54:NM0, PENB, *, PEGB1
			8'd6 : rdata = 44'b00011100000000001101111111000000000010010000;
			// PEs: 48, 50 -> 
			// srcs: (222, 6)(805) -9, (47) 4 --> (849) -36:PEGB0, ND2, *, 
			8'd7 : rdata = 44'b00011111000000000110000001000000000000000000;
			// PEs: 50, 50 -> 
			// srcs: (225, 10)(3) 1, (849) -36 --> (1049) -36:NM0, ALU, *, 
			8'd8 : rdata = 44'b00011100000000000011111111100000000000000000;
			// PEs: 50, 50 -> 50
			// srcs: (228, 13)(248) 9, (1049) -36 --> (1249) 45:NW2, ALU, -, NW2
			8'd9 : rdata = 44'b00010010000000100011111111100010100000000000;
			// PEs: 50, 49 -> 49
			// srcs: (236, 11)(3) 1, (863) -81 --> (1063) -81:NM0, PENB, *, PEGB1
			8'd10 : rdata = 44'b00011100000000001101111111000000000010010000;
			// PEs: 48, 50 -> 51
			// srcs: (237, 7)(805) -9, (62) 8 --> (864) -72:PEGB0, ND0, *, PENB
			8'd11 : rdata = 44'b00011111000000000110000000000000000100000000;
			// PEs: 50, 51 -> 50
			// srcs: (246, 14)(263) 5, (1064) -72 --> (1264) 77:NW0, PEGB3, -, NW0
			8'd12 : rdata = 44'b00010010000000001110000011000010000000000000;
			// PEs: 50, 49 -> 49
			// srcs: (314, 12)(3) 1, (941) -45 --> (1141) -45:NM0, PENB, *, PEGB1
			8'd13 : rdata = 44'b00011100000000001101111111000000000010010000;
			// PEs: 48, 50 -> 51
			// srcs: (315, 8)(805) -9, (140) 6 --> (942) -54:PEGB0, ND1, *, PENB
			8'd14 : rdata = 44'b00011111000000000110000000100000000100000000;
			// PEs: 50, 51 -> 50
			// srcs: (324, 15)(341) 7, (1142) -54 --> (1342) 61:NW1, PEGB3, -, NW1
			8'd15 : rdata = 44'b00010010000000011110000011000010010000000000;
			default : rdata = 44'b00000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 51) begin
	always @(*) begin
		case(address)
			// PEs: 51, 51 -> 52
			// srcs: (1, 0)(64) 5, (265) 6 --> (465) 30:ND0, NW0, *, PENB
			8'd0 : rdata = 44'b00011011000000000100000000000000000100000000;
			// PEs: 51, 51 -> 52
			// srcs: (2, 1)(142) 4, (343) 3 --> (543) 12:ND1, NW1, *, PENB
			8'd1 : rdata = 44'b00011011000000010100000000100000000100000000;
			// PEs: 51, 51 -> 48
			// srcs: (3, 2)(50) 9, (251) 1 --> (451) 9:ND2, NW2, *, PEGB0
			8'd2 : rdata = 44'b00011011000000100100000001000000000010000000;
			// PEs: 50, 54 -> 
			// srcs: (10, 3)(660) 40, (464) 14 --> (661) 54:PENB, PEGB6, +, 
			8'd3 : rdata = 44'b00001110111111101110000110000000000000000000;
			// PEs: 51, 53 -> 50
			// srcs: (16, 4)(661) 54, (663) 66 --> (664) 120:ALU, PEGB5, +, PEGB2
			8'd4 : rdata = 44'b00001001111111111110000101000000000010100000;
			// PEs: 48, 51 -> 
			// srcs: (225, 5)(805) -9, (50) 9 --> (852) -81:PEGB0, ND2, *, 
			8'd5 : rdata = 44'b00011111000000000110000001000000000000000000;
			// PEs: 51, 51 -> 
			// srcs: (228, 8)(3) 1, (852) -81 --> (1052) -81:NM0, ALU, *, 
			8'd6 : rdata = 44'b00011100000000000011111111100000000000000000;
			// PEs: 51, 51 -> 51
			// srcs: (231, 12)(251) 1, (1052) -81 --> (1252) 82:NW2, ALU, -, NW2
			8'd7 : rdata = 44'b00010010000000100011111111100010100000000000;
			// PEs: 48, 51 -> 52
			// srcs: (239, 6)(805) -9, (64) 5 --> (866) -45:PEGB0, ND0, *, PENB
			8'd8 : rdata = 44'b00011111000000000110000000000000000100000000;
			// PEs: 51, 50 -> 50
			// srcs: (240, 9)(3) 1, (864) -72 --> (1064) -72:NM0, PENB, *, PEGB2
			8'd9 : rdata = 44'b00011100000000001101111111000000000010100000;
			// PEs: 51, 52 -> 51
			// srcs: (248, 13)(265) 6, (1066) -45 --> (1266) 51:NW0, PEGB4, -, NW0
			8'd10 : rdata = 44'b00010010000000001110000100000010000000000000;
			// PEs: 48, 51 -> 51
			// srcs: (317, 7)(805) -9, (142) 4 --> (944) -36:PEGB0, ND1, *, NI0
			8'd11 : rdata = 44'b00011111000000000110000000110000000000000000;
			// PEs: 51, 50 -> 50
			// srcs: (318, 10)(3) 1, (942) -54 --> (1142) -54:NM0, PENB, *, PEGB2
			8'd12 : rdata = 44'b00011100000000001101111111000000000010100000;
			// PEs: 51, 51 -> 
			// srcs: (320, 11)(3) 1, (944) -36 --> (1144) -36:NM0, NI0, *, 
			8'd13 : rdata = 44'b00011100000000001010000000000000000000000000;
			// PEs: 51, 51 -> 51
			// srcs: (323, 14)(343) 3, (1144) -36 --> (1344) 39:NW1, ALU, -, NW1
			8'd14 : rdata = 44'b00010010000000010011111111100010010000000000;
			default : rdata = 44'b00000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 52) begin
	always @(*) begin
		case(address)
			// PEs: 52, 52 -> 52
			// srcs: (1, 0)(65) 9, (266) 1 --> (466) 9:ND0, NW0, *, NI0
			8'd0 : rdata = 44'b00011011000000000100000000010000000000000000;
			// PEs: 52, 52 -> 52
			// srcs: (2, 1)(143) 4, (344) 3 --> (544) 12:ND1, NW1, *, NI1
			8'd1 : rdata = 44'b00011011000000010100000000110100000000000000;
			// PEs: 52, 52 -> 49
			// srcs: (3, 2)(53) 9, (254) 6 --> (454) 54:ND2, NW2, *, PEGB1
			8'd2 : rdata = 44'b00011011000000100100000001000000000010010000;
			// PEs: 51, 52 -> 53
			// srcs: (4, 3)(465) 30, (466) 9 --> (662) 39:PENB, NI0, +, PENB
			8'd3 : rdata = 44'b00001110111111101010000000000000000100000000;
			// PEs: 51, 52 -> 48
			// srcs: (5, 4)(543) 12, (544) 12 --> (740) 24:PENB, NI1, +, PEGB0
			8'd4 : rdata = 44'b00001110111111101010000000100000000010000000;
			// PEs: 48, 52 -> 
			// srcs: (228, 5)(805) -9, (53) 9 --> (855) -81:PEGB0, ND2, *, 
			8'd5 : rdata = 44'b00011111000000000110000001000000000000000000;
			// PEs: 52, 52 -> 
			// srcs: (231, 8)(3) 1, (855) -81 --> (1055) -81:NM0, ALU, *, 
			8'd6 : rdata = 44'b00011100000000000011111111100000000000000000;
			// PEs: 52, 52 -> 52
			// srcs: (234, 11)(254) 6, (1055) -81 --> (1255) 87:NW2, ALU, -, NW2
			8'd7 : rdata = 44'b00010010000000100011111111100010100000000000;
			// PEs: 48, 52 -> 52
			// srcs: (240, 6)(805) -9, (65) 9 --> (867) -81:PEGB0, ND0, *, NI0
			8'd8 : rdata = 44'b00011111000000000110000000010000000000000000;
			// PEs: 52, 51 -> 51
			// srcs: (242, 9)(3) 1, (866) -45 --> (1066) -45:NM0, PENB, *, PEGB3
			8'd9 : rdata = 44'b00011100000000001101111111000000000010110000;
			// PEs: 52, 52 -> 
			// srcs: (243, 10)(3) 1, (867) -81 --> (1067) -81:NM0, NI0, *, 
			8'd10 : rdata = 44'b00011100000000001010000000000000000000000000;
			// PEs: 52, 52 -> 52
			// srcs: (246, 12)(266) 1, (1067) -81 --> (1267) 82:NW0, ALU, -, NW0
			8'd11 : rdata = 44'b00010010000000000011111111100010000000000000;
			// PEs: 48, 52 -> 53
			// srcs: (318, 7)(805) -9, (143) 4 --> (945) -36:PEGB0, ND1, *, PENB
			8'd12 : rdata = 44'b00011111000000000110000000100000000100000000;
			// PEs: 52, 53 -> 52
			// srcs: (327, 13)(344) 3, (1145) -36 --> (1345) 39:NW1, PEGB5, -, NW1
			8'd13 : rdata = 44'b00010010000000011110000101000010010000000000;
			default : rdata = 44'b00000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 53) begin
	always @(*) begin
		case(address)
			// PEs: 53, 53 -> 54
			// srcs: (1, 0)(67) 5, (268) 9 --> (468) 45:ND0, NW0, *, PENB
			8'd0 : rdata = 44'b00011011000000000100000000000000000100000000;
			// PEs: 53, 53 -> 54
			// srcs: (2, 1)(145) 8, (346) 4 --> (546) 32:ND1, NW1, *, PENB
			8'd1 : rdata = 44'b00011011000000010100000000100000000100000000;
			// PEs: 53, 53 -> 49
			// srcs: (3, 2)(60) 3, (261) 2 --> (461) 6:ND2, NW2, *, PEGB1
			8'd2 : rdata = 44'b00011011000000100100000001000000000010010000;
			// PEs: 52, 55 -> 51
			// srcs: (10, 3)(662) 39, (467) 27 --> (663) 66:PENB, PEGB7, +, PEGB3
			8'd3 : rdata = 44'b00001110111111101110000111000000000010110000;
			// PEs: 48 -> 
			// srcs: (65, 4)(748) 81 --> (748) 81:PEGB0, pass, 
			8'd4 : rdata = 44'b11000111000000000000000000000000000000000000;
			// PEs: 49, 53 -> 48
			// srcs: (67, 5)(746) 114, (748) 81 --> (749) 195:PEGB1, ALU, +, PEGB0
			8'd5 : rdata = 44'b00001111000000100011111111100000000010000000;
			// PEs: 48, 53 -> 
			// srcs: (235, 6)(805) -9, (60) 3 --> (862) -27:PEGB0, ND2, *, 
			8'd6 : rdata = 44'b00011111000000000110000001000000000000000000;
			// PEs: 53, 53 -> 
			// srcs: (238, 9)(3) 1, (862) -27 --> (1062) -27:NM0, ALU, *, 
			8'd7 : rdata = 44'b00011100000000000011111111100000000000000000;
			// PEs: 53, 53 -> 53
			// srcs: (241, 11)(261) 2, (1062) -27 --> (1262) 29:NW2, ALU, -, NW2
			8'd8 : rdata = 44'b00010010000000100011111111100010100000000000;
			// PEs: 48, 53 -> 54
			// srcs: (242, 7)(805) -9, (67) 5 --> (869) -45:PEGB0, ND0, *, PENB
			8'd9 : rdata = 44'b00011111000000000110000000000000000100000000;
			// PEs: 53, 54 -> 53
			// srcs: (251, 12)(268) 9, (1069) -45 --> (1269) 54:NW0, PEGB6, -, NW0
			8'd10 : rdata = 44'b00010010000000001110000110000010000000000000;
			// PEs: 48, 53 -> 54
			// srcs: (320, 8)(805) -9, (145) 8 --> (947) -72:PEGB0, ND1, *, PENB
			8'd11 : rdata = 44'b00011111000000000110000000100000000100000000;
			// PEs: 53, 52 -> 52
			// srcs: (321, 10)(3) 1, (945) -36 --> (1145) -36:NM0, PENB, *, PEGB4
			8'd12 : rdata = 44'b00011100000000001101111111000000000011000000;
			// PEs: 53, 54 -> 53
			// srcs: (329, 13)(346) 4, (1147) -72 --> (1347) 76:NW1, PEGB6, -, NW1
			8'd13 : rdata = 44'b00010010000000011110000110000010010000000000;
			default : rdata = 44'b00000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 54) begin
	always @(*) begin
		case(address)
			// PEs: 54, 54 -> 54
			// srcs: (1, 0)(68) 1, (269) 3 --> (469) 3:ND0, NW0, *, NI0
			8'd0 : rdata = 44'b00011011000000000100000000010000000000000000;
			// PEs: 54, 54 -> 54
			// srcs: (2, 1)(146) 1, (347) 0 --> (547) 0:ND1, NW1, *, NI1
			8'd1 : rdata = 44'b00011011000000010100000000110100000000000000;
			// PEs: 54, 54 -> 51
			// srcs: (3, 2)(63) 2, (264) 7 --> (464) 14:ND2, NW2, *, PEGB3
			8'd2 : rdata = 44'b00011011000000100100000001000000000010110000;
			// PEs: 53, 54 -> 48
			// srcs: (4, 3)(468) 45, (469) 3 --> (666) 48:PENB, NI0, +, PEGB0
			8'd3 : rdata = 44'b00001110111111101010000000000000000010000000;
			// PEs: 53, 54 -> 48
			// srcs: (5, 4)(546) 32, (547) 0 --> (742) 32:PENB, NI1, +, PEGB0
			8'd4 : rdata = 44'b00001110111111101010000000100000000010000000;
			// PEs: 48, 54 -> 
			// srcs: (238, 5)(805) -9, (63) 2 --> (865) -18:PEGB0, ND2, *, 
			8'd5 : rdata = 44'b00011111000000000110000001000000000000000000;
			// PEs: 54, 54 -> 54
			// srcs: (241, 8)(3) 1, (865) -18 --> (1065) -18:NM0, ALU, *, NI0
			8'd6 : rdata = 44'b00011100000000000011111111110000000000000000;
			// PEs: 48, 54 -> 55
			// srcs: (243, 6)(805) -9, (68) 1 --> (870) -9:PEGB0, ND0, *, PENB
			8'd7 : rdata = 44'b00011111000000000110000000000000000100000000;
			// PEs: 54, 54 -> 54
			// srcs: (244, 12)(264) 7, (1065) -18 --> (1265) 25:NW2, NI0, -, NW2
			8'd8 : rdata = 44'b00010010000000101010000000000010100000000000;
			// PEs: 54, 53 -> 53
			// srcs: (245, 9)(3) 1, (869) -45 --> (1069) -45:NM0, PENB, *, PEGB5
			8'd9 : rdata = 44'b00011100000000001101111111000000000011010000;
			// PEs: 54, 55 -> 54
			// srcs: (252, 13)(269) 3, (1070) -9 --> (1270) 12:NW0, PEGB7, -, NW0
			8'd10 : rdata = 44'b00010010000000001110000111000010000000000000;
			// PEs: 48, 54 -> 54
			// srcs: (321, 7)(805) -9, (146) 1 --> (948) -9:PEGB0, ND1, *, NI0
			8'd11 : rdata = 44'b00011111000000000110000000110000000000000000;
			// PEs: 54, 53 -> 53
			// srcs: (323, 10)(3) 1, (947) -72 --> (1147) -72:NM0, PENB, *, PEGB5
			8'd12 : rdata = 44'b00011100000000001101111111000000000011010000;
			// PEs: 54, 54 -> 
			// srcs: (324, 11)(3) 1, (948) -9 --> (1148) -9:NM0, NI0, *, 
			8'd13 : rdata = 44'b00011100000000001010000000000000000000000000;
			// PEs: 54, 54 -> 54
			// srcs: (327, 14)(347) 0, (1148) -9 --> (1348) 9:NW1, ALU, -, NW1
			8'd14 : rdata = 44'b00010010000000010011111111100010010000000000;
			default : rdata = 44'b00000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 55) begin
	always @(*) begin
		case(address)
			// PEs: 55, 55 -> 48
			// srcs: (1, 0)(70) 2, (271) 4 --> (471) 8:ND0, NW0, *, PENB
			8'd0 : rdata = 44'b00011011000000000100000000000000000100000000;
			// PEs: 55, 55 -> 48
			// srcs: (2, 1)(148) 6, (349) 8 --> (549) 48:ND1, NW1, *, PENB
			8'd1 : rdata = 44'b00011011000000010100000000100000000100000000;
			// PEs: 55, 55 -> 53
			// srcs: (3, 2)(66) 3, (267) 9 --> (467) 27:ND2, NW2, *, PEGB5
			8'd2 : rdata = 44'b00011011000000100100000001000000000011010000;
			// PEs: 49 -> 
			// srcs: (33, 3)(609) 9 --> (609) 9:PEGB1, pass, 
			8'd3 : rdata = 44'b11000111000000100000000000000000000000000000;
			// PEs: 48, 55 -> 48
			// srcs: (43, 4)(607) 74, (609) 9 --> (610) 83:PEGB0, ALU, +, PENB
			8'd4 : rdata = 44'b00001111000000000011111111100000000100000000;
			// PEs: 48, 55 -> 
			// srcs: (241, 5)(805) -9, (66) 3 --> (868) -27:PEGB0, ND2, *, 
			8'd5 : rdata = 44'b00011111000000000110000001000000000000000000;
			// PEs: 55, 55 -> 55
			// srcs: (244, 8)(3) 1, (868) -27 --> (1068) -27:NM0, ALU, *, NI0
			8'd6 : rdata = 44'b00011100000000000011111111110000000000000000;
			// PEs: 48, 55 -> 55
			// srcs: (245, 6)(805) -9, (70) 2 --> (872) -18:PEGB0, ND0, *, NI1
			8'd7 : rdata = 44'b00011111000000000110000000010100000000000000;
			// PEs: 55, 54 -> 54
			// srcs: (246, 9)(3) 1, (870) -9 --> (1070) -9:NM0, PENB, *, PEGB6
			8'd8 : rdata = 44'b00011100000000001101111111000000000011100000;
			// PEs: 55, 55 -> 55
			// srcs: (247, 12)(267) 9, (1068) -27 --> (1268) 36:NW2, NI0, -, NW2
			8'd9 : rdata = 44'b00010010000000101010000000000010100000000000;
			// PEs: 55, 55 -> 
			// srcs: (248, 10)(3) 1, (872) -18 --> (1072) -18:NM0, NI1, *, 
			8'd10 : rdata = 44'b00011100000000001010000000100000000000000000;
			// PEs: 55, 55 -> 55
			// srcs: (251, 13)(271) 4, (1072) -18 --> (1272) 22:NW0, ALU, -, NW0
			8'd11 : rdata = 44'b00010010000000000011111111100010000000000000;
			// PEs: 48, 55 -> 
			// srcs: (323, 7)(805) -9, (148) 6 --> (950) -54:PEGB0, ND1, *, 
			8'd12 : rdata = 44'b00011111000000000110000000100000000000000000;
			// PEs: 55, 55 -> 
			// srcs: (326, 11)(3) 1, (950) -54 --> (1150) -54:NM0, ALU, *, 
			8'd13 : rdata = 44'b00011100000000000011111111100000000000000000;
			// PEs: 55, 55 -> 55
			// srcs: (329, 14)(349) 8, (1150) -54 --> (1350) 62:NW1, ALU, -, NW1
			8'd14 : rdata = 44'b00010010000000010011111111100010010000000000;
			default : rdata = 44'b00000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 56) begin
	always @(*) begin
		case(address)
			// PEs: 48 -> 57
			// srcs: (5, 0)(471) 8 --> (471) 8:PUNB, pass, PENB
			8'd0 : rdata = 44'b11000110111111110000000000000000000100000000;
			// PEs: 48 -> 57
			// srcs: (6, 1)(549) 48 --> (549) 48:PUNB, pass, PENB
			8'd1 : rdata = 44'b11000110111111110000000000000000000100000000;
			// PEs: 63 -> 0
			// srcs: (7, 6)(678) 62 --> (678) 62:PENB, pass, PUNB
			8'd2 : rdata = 44'b11000110111111100000000000000000001000000000;
			// PEs: 61 -> 0
			// srcs: (8, 7)(486) 72 --> (486) 72:PEGB5, pass, PUNB
			8'd3 : rdata = 44'b11000111000010100000000000000000001000000000;
			// PEs: 62 -> 0
			// srcs: (9, 8)(489) 32 --> (489) 32:PEGB6, pass, PUNB
			8'd4 : rdata = 44'b11000111000011000000000000000000001000000000;
			// PEs: 59 -> 40
			// srcs: (10, 17)(747) 67 --> (747) 67:PEGB3, pass, PUGB5
			8'd5 : rdata = 44'b11000111000001100000000000000000000000001101;
			// PEs: 63 -> 8
			// srcs: (14, 9)(492) 0 --> (492) 0:PENB, pass, PUGB1
			8'd6 : rdata = 44'b11000110111111100000000000000000000000001001;
			// PEs: 57 -> 48
			// srcs: (15, 16)(745) 93 --> (745) 93:PEGB1, pass, PUGB6
			8'd7 : rdata = 44'b11000111000000100000000000000000000000001110;
			// PEs: 62 -> 0
			// srcs: (16, 24)(755) 48 --> (755) 48:PEGB6, pass, PUNB
			8'd8 : rdata = 44'b11000111000011000000000000000000001000000000;
			// PEs: 16 -> 56
			// srcs: (20, 2)(624) 48 --> (624) 48:PUGB2, pass, NI0
			8'd9 : rdata = 44'b11000111000001010000000000010000000000000000;
			// PEs: 40 -> 57
			// srcs: (21, 3)(429) 4 --> (429) 4:PUGB5, pass, PENB
			8'd10 : rdata = 44'b11000111000010110000000000000000000100000000;
			// PEs: 56 -> 57
			// srcs: (27, 4)(624) 48 --> (624) 48:NI0, pass, PENB
			8'd11 : rdata = 44'b11000101000000000000000000000000000100000000;
			// PEs: 48 -> 57
			// srcs: (28, 5)(666) 48 --> (666) 48:PUNB, pass, PENB
			8'd12 : rdata = 44'b11000110111111110000000000000000000100000000;
			// PEs: 24 -> 56
			// srcs: (29, 10)(707) 30 --> (707) 30:PUGB3, pass, NI0
			8'd13 : rdata = 44'b11000111000001110000000000010000000000000000;
			// PEs: 0 -> 57
			// srcs: (30, 11)(511) 14 --> (511) 14:PUGB0, pass, PENB
			8'd14 : rdata = 44'b11000111000000010000000000000000000100000000;
			// PEs: 56 -> 57
			// srcs: (36, 12)(707) 30 --> (707) 30:NI0, pass, PENB
			8'd15 : rdata = 44'b11000101000000000000000000000000000100000000;
			// PEs: 48 -> 56
			// srcs: (37, 13)(740) 24 --> (740) 24:PUNB, pass, NI0
			8'd16 : rdata = 44'b11000110111111110000000000010000000000000000;
			// PEs: 16 -> 57
			// srcs: (42, 14)(545) 36 --> (545) 36:PUGB2, pass, PENB
			8'd17 : rdata = 44'b11000111000001010000000000000000000100000000;
			// PEs: 56 -> 57
			// srcs: (48, 15)(740) 24 --> (740) 24:NI0, pass, PENB
			8'd18 : rdata = 44'b11000101000000000000000000000000000100000000;
			// PEs: 0 -> 56
			// srcs: (49, 18)(759) 57 --> (759) 57:PUGB0, pass, NI0
			8'd19 : rdata = 44'b11000111000000010000000000010000000000000000;
			// PEs: 16 -> 57
			// srcs: (50, 19)(564) 0 --> (564) 0:PUGB2, pass, PENB
			8'd20 : rdata = 44'b11000111000001010000000000000000000100000000;
			// PEs: 57 -> 24
			// srcs: (55, 23)(741) 60 --> (741) 60:PEGB1, pass, PUGB3
			8'd21 : rdata = 44'b11000111000000100000000000000000000000001011;
			// PEs: 56 -> 57
			// srcs: (56, 20)(759) 57 --> (759) 57:NI0, pass, PENB
			8'd22 : rdata = 44'b11000101000000000000000000000000000100000000;
			// PEs: 48 -> 57
			// srcs: (57, 21)(623) 46 --> (623) 46:PUNB, pass, PENB
			8'd23 : rdata = 44'b11000110111111110000000000000000000100000000;
			// PEs: 57 -> 0
			// srcs: (63, 25)(760) 57 --> (760) 57:PEGB1, pass, PUNB
			8'd24 : rdata = 44'b11000111000000100000000000000000001000000000;
			// PEs: 16 -> 57
			// srcs: (67, 22)(706) 11 --> (706) 11:PUGB2, pass, PENB
			8'd25 : rdata = 44'b11000111000001010000000000000000000100000000;
			// PEs: 40 -> 57
			// srcs: (68, 26)(621) 218 --> (621) 218:PUGB5, pass, PENB
			8'd26 : rdata = 44'b11000111000010110000000000000000000100000000;
			// PEs: 24 -> 57
			// srcs: (69, 27)(714) 89 --> (714) 89:PUGB3, pass, PENB
			8'd27 : rdata = 44'b11000111000001110000000000000000000100000000;
			// PEs: 57 -> 8
			// srcs: (77, 31)(627) 316 --> (627) 316:PEGB1, pass, PUGB1
			8'd28 : rdata = 44'b11000111000000100000000000000000000000001001;
			// PEs: 57 -> 40
			// srcs: (87, 33)(715) 144 --> (715) 144:PEGB1, pass, PUGB5
			8'd29 : rdata = 44'b11000111000000100000000000000000000000001101;
			// PEs: 24 -> 56
			// srcs: (97, 28)(744) 92 --> (744) 92:PUGB3, pass, NI0
			8'd30 : rdata = 44'b11000111000001110000000000010000000000000000;
			// PEs: 48 -> 57
			// srcs: (98, 29)(749) 195 --> (749) 195:PUNB, pass, PENB
			8'd31 : rdata = 44'b11000110111111110000000000000000000100000000;
			// PEs: 56 -> 57
			// srcs: (104, 30)(744) 92 --> (744) 92:NI0, pass, PENB
			8'd32 : rdata = 44'b11000101000000000000000000000000000100000000;
			// PEs: 48 -> 57
			// srcs: (105, 32)(665) 184 --> (665) 184:PUNB, pass, PENB
			8'd33 : rdata = 44'b11000110111111110000000000000000000100000000;
			// PEs: 48 -> 57
			// srcs: (106, 34)(739) 437 --> (739) 437:PUNB, pass, PENB
			8'd34 : rdata = 44'b11000110111111110000000000000000000100000000;
			// PEs: 57 -> 24
			// srcs: (112, 35)(677) 325 --> (677) 325:PEGB1, pass, PUGB3
			8'd35 : rdata = 44'b11000111000000100000000000000000000000001011;
			// PEs: 57 -> 40
			// srcs: (121, 36)(751) 724 --> (751) 724:PEGB1, pass, PUGB5
			8'd36 : rdata = 44'b11000111000000100000000000000000000000001101;
			// PEs: 0 -> 57
			// srcs: (239, 37)(805) -9 --> (805) -9:PUGB0, pass, PENB
			8'd37 : rdata = 44'b11000111000000010000000000000000000100000000;
			// PEs: 0 -> 57
			// srcs: (241, 38)(805) -9 --> (805) -9:PUGB0, pass, PENB
			8'd38 : rdata = 44'b11000111000000010000000000000000000100000000;
			// PEs: 0 -> 58
			// srcs: (242, 39)(805) -9 --> (805) -9:PUGB0, pass, PEGB2
			8'd39 : rdata = 44'b11000111000000010000000000000000000010100000;
			// PEs: 0 -> 58
			// srcs: (243, 40)(805) -9 --> (805) -9:PUGB0, pass, PEGB2
			8'd40 : rdata = 44'b11000111000000010000000000000000000010100000;
			// PEs: 0 -> 59
			// srcs: (244, 41)(805) -9 --> (805) -9:PUGB0, pass, PEGB3
			8'd41 : rdata = 44'b11000111000000010000000000000000000010110000;
			// PEs: 0 -> 59
			// srcs: (245, 42)(805) -9 --> (805) -9:PUGB0, pass, PEGB3
			8'd42 : rdata = 44'b11000111000000010000000000000000000010110000;
			// PEs: 0 -> 60
			// srcs: (246, 43)(805) -9 --> (805) -9:PUGB0, pass, PEGB4
			8'd43 : rdata = 44'b11000111000000010000000000000000000011000000;
			// PEs: 0 -> 61
			// srcs: (247, 44)(805) -9 --> (805) -9:PUGB0, pass, PEGB5
			8'd44 : rdata = 44'b11000111000000010000000000000000000011010000;
			// PEs: 0 -> 60
			// srcs: (248, 45)(805) -9 --> (805) -9:PUGB0, pass, PEGB4
			8'd45 : rdata = 44'b11000111000000010000000000000000000011000000;
			// PEs: 0 -> 62
			// srcs: (249, 46)(805) -9 --> (805) -9:PUGB0, pass, PEGB6
			8'd46 : rdata = 44'b11000111000000010000000000000000000011100000;
			// PEs: 0 -> 63
			// srcs: (250, 47)(805) -9 --> (805) -9:PUGB0, pass, PEGB7
			8'd47 : rdata = 44'b11000111000000010000000000000000000011110000;
			// PEs: 0 -> 61
			// srcs: (255, 48)(805) -9 --> (805) -9:PUGB0, pass, PEGB5
			8'd48 : rdata = 44'b11000111000000010000000000000000000011010000;
			// PEs: 0 -> 62
			// srcs: (258, 49)(805) -9 --> (805) -9:PUGB0, pass, PEGB6
			8'd49 : rdata = 44'b11000111000000010000000000000000000011100000;
			// PEs: 0 -> 63
			// srcs: (261, 50)(805) -9 --> (805) -9:PUGB0, pass, PEGB7
			8'd50 : rdata = 44'b11000111000000010000000000000000000011110000;
			// PEs: 0 -> 57
			// srcs: (319, 51)(805) -9 --> (805) -9:PUGB0, pass, PENB
			8'd51 : rdata = 44'b11000111000000010000000000000000000100000000;
			// PEs: 0 -> 58
			// srcs: (321, 52)(805) -9 --> (805) -9:PUGB0, pass, PEGB2
			8'd52 : rdata = 44'b11000111000000010000000000000000000010100000;
			// PEs: 0 -> 59
			// srcs: (322, 53)(805) -9 --> (805) -9:PUGB0, pass, PEGB3
			8'd53 : rdata = 44'b11000111000000010000000000000000000010110000;
			// PEs: 0 -> 60
			// srcs: (324, 54)(805) -9 --> (805) -9:PUGB0, pass, PEGB4
			8'd54 : rdata = 44'b11000111000000010000000000000000000011000000;
			// PEs: 0 -> 61
			// srcs: (325, 55)(805) -9 --> (805) -9:PUGB0, pass, PEGB5
			8'd55 : rdata = 44'b11000111000000010000000000000000000011010000;
			// PEs: 0 -> 62
			// srcs: (326, 56)(805) -9 --> (805) -9:PUGB0, pass, PEGB6
			8'd56 : rdata = 44'b11000111000000010000000000000000000011100000;
			// PEs: 0 -> 63
			// srcs: (327, 57)(805) -9 --> (805) -9:PUGB0, pass, PEGB7
			8'd57 : rdata = 44'b11000111000000010000000000000000000011110000;
			default : rdata = 44'b00000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 57) begin
	always @(*) begin
		case(address)
			// PEs: 57, 57 -> 57
			// srcs: (1, 0)(71) 5, (272) 3 --> (472) 15:ND0, NW0, *, NI0
			8'd0 : rdata = 44'b00011011000000000100000000010000000000000000;
			// PEs: 57, 57 -> 57
			// srcs: (2, 1)(149) 5, (350) 9 --> (550) 45:ND1, NW1, *, NI1
			8'd1 : rdata = 44'b00011011000000010100000000110100000000000000;
			// PEs: 57, 57 -> 57
			// srcs: (3, 2)(69) 6, (270) 4 --> (470) 24:ND2, NW2, *, NI2
			8'd2 : rdata = 44'b00011011000000100100000001011000000000000000;
			// PEs: 56, 57 -> 58
			// srcs: (8, 3)(471) 8, (472) 15 --> (668) 23:PENB, NI0, +, PENB
			8'd3 : rdata = 44'b00001110111111101010000000000000000100000000;
			// PEs: 56, 57 -> 56
			// srcs: (9, 4)(549) 48, (550) 45 --> (745) 93:PENB, NI1, +, PEGB0
			8'd4 : rdata = 44'b00001110111111101010000000100000000010000000;
			// PEs: 56 -> 
			// srcs: (23, 5)(429) 4 --> (429) 4:PENB, pass, 
			8'd5 : rdata = 44'b11000110111111100000000000000000000000000000;
			// PEs: 56, 57 -> 57
			// srcs: (29, 6)(624) 48, (429) 4 --> (625) 52:PENB, ALU, +, NI0
			8'd6 : rdata = 44'b00001110111111100011111111110000000000000000;
			// PEs: 56, 57 -> 58
			// srcs: (30, 7)(666) 48, (470) 24 --> (667) 72:PENB, NI2, +, PENB
			8'd7 : rdata = 44'b00001110111111101010000001000000000100000000;
			// PEs: 56 -> 
			// srcs: (32, 8)(511) 14 --> (511) 14:PENB, pass, 
			8'd8 : rdata = 44'b11000110111111100000000000000000000000000000;
			// PEs: 56, 57 -> 57
			// srcs: (38, 9)(707) 30, (511) 14 --> (708) 44:PENB, ALU, +, NI1
			8'd9 : rdata = 44'b00001110111111100011111111110100000000000000;
			// PEs: 56 -> 
			// srcs: (44, 10)(545) 36 --> (545) 36:PENB, pass, 
			8'd10 : rdata = 44'b11000110111111100000000000000000000000000000;
			// PEs: 56, 57 -> 56
			// srcs: (50, 11)(740) 24, (545) 36 --> (741) 60:PENB, ALU, +, PEGB0
			8'd11 : rdata = 44'b00001110111111100011111111100000000010000000;
			// PEs: 56 -> 
			// srcs: (52, 12)(564) 0 --> (564) 0:PENB, pass, 
			8'd12 : rdata = 44'b11000110111111100000000000000000000000000000;
			// PEs: 56, 57 -> 56
			// srcs: (58, 13)(759) 57, (564) 0 --> (760) 57:PENB, ALU, +, PEGB0
			8'd13 : rdata = 44'b00001110111111100011111111100000000010000000;
			// PEs: 56, 57 -> 57
			// srcs: (59, 14)(623) 46, (625) 52 --> (626) 98:PENB, NI0, +, NI2
			8'd14 : rdata = 44'b00001110111111101010000000011000000000000000;
			// PEs: 56, 57 -> 57
			// srcs: (69, 15)(706) 11, (708) 44 --> (709) 55:PENB, NI1, +, NI0
			8'd15 : rdata = 44'b00001110111111101010000000110000000000000000;
			// PEs: 56, 57 -> 56
			// srcs: (72, 16)(621) 218, (626) 98 --> (627) 316:PENB, NI2, +, PEGB0
			8'd16 : rdata = 44'b00001110111111101010000001000000000010000000;
			// PEs: 57, 56 -> 56
			// srcs: (82, 17)(709) 55, (714) 89 --> (715) 144:NI0, PENB, +, PEGB0
			8'd17 : rdata = 44'b00001101000000001101111111000000000010000000;
			// PEs: 56 -> 
			// srcs: (100, 18)(749) 195 --> (749) 195:PENB, pass, 
			8'd18 : rdata = 44'b11000110111111100000000000000000000000000000;
			// PEs: 56, 57 -> 57
			// srcs: (106, 19)(744) 92, (749) 195 --> (750) 287:PENB, ALU, +, NI0
			8'd19 : rdata = 44'b00001110111111100011111111110000000000000000;
			// PEs: 56, 62 -> 56
			// srcs: (107, 20)(665) 184, (676) 141 --> (677) 325:PENB, PEGB6, +, PEGB0
			8'd20 : rdata = 44'b00001110111111101110000110000000000010000000;
			// PEs: 56, 57 -> 56
			// srcs: (116, 21)(739) 437, (750) 287 --> (751) 724:PENB, NI0, +, PEGB0
			8'd21 : rdata = 44'b00001110111111101010000000000000000010000000;
			// PEs: 56, 57 -> 58
			// srcs: (241, 22)(805) -9, (69) 6 --> (871) -54:PENB, ND2, *, PENB
			8'd22 : rdata = 44'b00011110111111100110000001000000000100000000;
			// PEs: 56, 57 -> 58
			// srcs: (243, 23)(805) -9, (71) 5 --> (873) -45:PENB, ND0, *, PENB
			8'd23 : rdata = 44'b00011110111111100110000000000000000100000000;
			// PEs: 57, 58 -> 57
			// srcs: (250, 25)(270) 4, (1071) -54 --> (1271) 58:NW2, PEGB2, -, NW2
			8'd24 : rdata = 44'b00010010000000101110000010000010100000000000;
			// PEs: 57, 58 -> 57
			// srcs: (252, 26)(272) 3, (1073) -45 --> (1273) 48:NW0, PEGB2, -, NW0
			8'd25 : rdata = 44'b00010010000000001110000010000010000000000000;
			// PEs: 56, 57 -> 58
			// srcs: (321, 24)(805) -9, (149) 5 --> (951) -45:PENB, ND1, *, PENB
			8'd26 : rdata = 44'b00011110111111100110000000100000000100000000;
			// PEs: 57, 58 -> 57
			// srcs: (330, 27)(350) 9, (1151) -45 --> (1351) 54:NW1, PEGB2, -, NW1
			8'd27 : rdata = 44'b00010010000000011110000010000010010000000000;
			default : rdata = 44'b00000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 58) begin
	always @(*) begin
		case(address)
			// PEs: 58, 58 -> 59
			// srcs: (1, 0)(73) 5, (274) 6 --> (474) 30:ND0, NW0, *, PENB
			8'd0 : rdata = 44'b00011011000000000100000000000000000100000000;
			// PEs: 58, 58 -> 59
			// srcs: (2, 1)(151) 7, (352) 7 --> (552) 49:ND1, NW1, *, PENB
			8'd1 : rdata = 44'b00011011000000010100000000100000000100000000;
			// PEs: 58, 58 -> 
			// srcs: (3, 2)(72) 1, (273) 5 --> (473) 5:ND2, NW2, *, 
			8'd2 : rdata = 44'b00011011000000100100000001000000000000000000;
			// PEs: 57, 58 -> 
			// srcs: (11, 3)(668) 23, (473) 5 --> (669) 28:PENB, ALU, +, 
			8'd3 : rdata = 44'b00001110111111100011111111100000000000000000;
			// PEs: 57, 58 -> 62
			// srcs: (33, 4)(667) 72, (669) 28 --> (670) 100:PENB, ALU, +, PEGB6
			8'd4 : rdata = 44'b00001110111111100011111111100000000011100000;
			// PEs: 58, 57 -> 57
			// srcs: (244, 8)(3) 1, (871) -54 --> (1071) -54:NM0, PENB, *, PEGB1
			8'd5 : rdata = 44'b00011100000000001101111111000000000010010000;
			// PEs: 58, 57 -> 57
			// srcs: (246, 9)(3) 1, (873) -45 --> (1073) -45:NM0, PENB, *, PEGB1
			8'd6 : rdata = 44'b00011100000000001101111111000000000010010000;
			// PEs: 56, 58 -> 58
			// srcs: (247, 5)(805) -9, (72) 1 --> (874) -9:PEGB0, ND2, *, NI0
			8'd7 : rdata = 44'b00011111000000000110000001010000000000000000;
			// PEs: 56, 58 -> 59
			// srcs: (248, 6)(805) -9, (73) 5 --> (875) -45:PEGB0, ND0, *, PENB
			8'd8 : rdata = 44'b00011111000000000110000000000000000100000000;
			// PEs: 58, 58 -> 
			// srcs: (250, 10)(3) 1, (874) -9 --> (1074) -9:NM0, NI0, *, 
			8'd9 : rdata = 44'b00011100000000001010000000000000000000000000;
			// PEs: 58, 58 -> 58
			// srcs: (253, 12)(273) 5, (1074) -9 --> (1274) 14:NW2, ALU, -, NW2
			8'd10 : rdata = 44'b00010010000000100011111111100010100000000000;
			// PEs: 58, 59 -> 58
			// srcs: (257, 13)(274) 6, (1075) -45 --> (1275) 51:NW0, PEGB3, -, NW0
			8'd11 : rdata = 44'b00010010000000001110000011000010000000000000;
			// PEs: 58, 57 -> 57
			// srcs: (324, 11)(3) 1, (951) -45 --> (1151) -45:NM0, PENB, *, PEGB1
			8'd12 : rdata = 44'b00011100000000001101111111000000000010010000;
			// PEs: 56, 58 -> 59
			// srcs: (326, 7)(805) -9, (151) 7 --> (953) -63:PEGB0, ND1, *, PENB
			8'd13 : rdata = 44'b00011111000000000110000000100000000100000000;
			// PEs: 58, 59 -> 58
			// srcs: (335, 14)(352) 7, (1153) -63 --> (1353) 70:NW1, PEGB3, -, NW1
			8'd14 : rdata = 44'b00010010000000011110000011000010010000000000;
			default : rdata = 44'b00000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 59) begin
	always @(*) begin
		case(address)
			// PEs: 59, 59 -> 59
			// srcs: (1, 0)(74) 0, (275) 1 --> (475) 0:ND0, NW0, *, NI0
			8'd0 : rdata = 44'b00011011000000000100000000010000000000000000;
			// PEs: 59, 59 -> 59
			// srcs: (2, 1)(152) 6, (353) 3 --> (553) 18:ND1, NW1, *, NI1
			8'd1 : rdata = 44'b00011011000000010100000000110100000000000000;
			// PEs: 59, 59 -> 59
			// srcs: (3, 2)(75) 1, (276) 1 --> (476) 1:ND2, NW2, *, NI2
			8'd2 : rdata = 44'b00011011000000100100000001011000000000000000;
			// PEs: 58, 59 -> 60
			// srcs: (4, 3)(474) 30, (475) 0 --> (671) 30:PENB, NI0, +, PENB
			8'd3 : rdata = 44'b00001110111111101010000000000000000100000000;
			// PEs: 58, 59 -> 56
			// srcs: (5, 4)(552) 49, (553) 18 --> (747) 67:PENB, NI1, +, PEGB0
			8'd4 : rdata = 44'b00001110111111101010000000100000000010000000;
			// PEs: 59 -> 60
			// srcs: (11, 5)(476) 1 --> (476) 1:NI2, pass, PENB
			8'd5 : rdata = 44'b11000101000000100000000000000000000100000000;
			// PEs: 56, 59 -> 60
			// srcs: (249, 6)(805) -9, (74) 0 --> (876) 0:PEGB0, ND0, *, PENB
			8'd6 : rdata = 44'b00011111000000000110000000000000000100000000;
			// PEs: 56, 59 -> 59
			// srcs: (250, 7)(805) -9, (75) 1 --> (877) -9:PEGB0, ND2, *, NI0
			8'd7 : rdata = 44'b00011111000000000110000001010000000000000000;
			// PEs: 59, 58 -> 58
			// srcs: (251, 9)(3) 1, (875) -45 --> (1075) -45:NM0, PENB, *, PEGB2
			8'd8 : rdata = 44'b00011100000000001101111111000000000010100000;
			// PEs: 59, 59 -> 
			// srcs: (253, 10)(3) 1, (877) -9 --> (1077) -9:NM0, NI0, *, 
			8'd9 : rdata = 44'b00011100000000001010000000000000000000000000;
			// PEs: 59, 59 -> 59
			// srcs: (256, 13)(276) 1, (1077) -9 --> (1277) 10:NW2, ALU, -, NW2
			8'd10 : rdata = 44'b00010010000000100011111111100010100000000000;
			// PEs: 59, 60 -> 59
			// srcs: (258, 12)(275) 1, (1076) 0 --> (1276) 1:NW0, PEGB4, -, NW0
			8'd11 : rdata = 44'b00010010000000001110000100000010000000000000;
			// PEs: 56, 59 -> 60
			// srcs: (327, 8)(805) -9, (152) 6 --> (954) -54:PEGB0, ND1, *, PENB
			8'd12 : rdata = 44'b00011111000000000110000000100000000100000000;
			// PEs: 59, 58 -> 58
			// srcs: (329, 11)(3) 1, (953) -63 --> (1153) -63:NM0, PENB, *, PEGB2
			8'd13 : rdata = 44'b00011100000000001101111111000000000010100000;
			// PEs: 59, 60 -> 59
			// srcs: (336, 14)(353) 3, (1154) -54 --> (1354) 57:NW1, PEGB4, -, NW1
			8'd14 : rdata = 44'b00010010000000011110000100000010010000000000;
			default : rdata = 44'b00000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 60) begin
	always @(*) begin
		case(address)
			// PEs: 60, 60 -> 61
			// srcs: (1, 0)(76) 1, (277) 0 --> (477) 0:ND0, NW0, *, PENB
			8'd0 : rdata = 44'b00011011000000000100000000000000000100000000;
			// PEs: 60, 60 -> 61
			// srcs: (2, 1)(154) 0, (355) 3 --> (555) 0:ND1, NW1, *, PENB
			8'd1 : rdata = 44'b00011011000000010100000000100000000100000000;
			// PEs: 60, 60 -> 61
			// srcs: (3, 2)(78) 2, (279) 5 --> (479) 10:ND2, NW2, *, PENB
			8'd2 : rdata = 44'b00011011000000100100000001000000000100000000;
			// PEs: 59 -> 
			// srcs: (6, 3)(671) 30 --> (671) 30:PENB, pass, 
			8'd3 : rdata = 44'b11000110111111100000000000000000000000000000;
			// PEs: 60, 59 -> 61
			// srcs: (13, 4)(671) 30, (476) 1 --> (672) 31:ALU, PENB, +, PENB
			8'd4 : rdata = 44'b00001001111111111101111111000000000100000000;
			// PEs: 56, 60 -> 60
			// srcs: (251, 5)(805) -9, (76) 1 --> (878) -9:PEGB0, ND0, *, NI0
			8'd5 : rdata = 44'b00011111000000000110000000010000000000000000;
			// PEs: 60, 59 -> 59
			// srcs: (252, 8)(3) 1, (876) 0 --> (1076) 0:NM0, PENB, *, PEGB3
			8'd6 : rdata = 44'b00011100000000001101111111000000000010110000;
			// PEs: 56, 60 -> 60
			// srcs: (253, 6)(805) -9, (78) 2 --> (880) -18:PEGB0, ND2, *, NI1
			8'd7 : rdata = 44'b00011111000000000110000001010100000000000000;
			// PEs: 60, 60 -> 60
			// srcs: (254, 9)(3) 1, (878) -9 --> (1078) -9:NM0, NI0, *, NI2
			8'd8 : rdata = 44'b00011100000000001010000000011000000000000000;
			// PEs: 60, 60 -> 60
			// srcs: (256, 10)(3) 1, (880) -18 --> (1080) -18:NM0, NI1, *, NI0
			8'd9 : rdata = 44'b00011100000000001010000000110000000000000000;
			// PEs: 60, 60 -> 60
			// srcs: (257, 12)(277) 0, (1078) -9 --> (1278) 9:NW0, NI2, -, NW0
			8'd10 : rdata = 44'b00010010000000001010000001000010000000000000;
			// PEs: 60, 60 -> 60
			// srcs: (259, 13)(279) 5, (1080) -18 --> (1280) 23:NW2, NI0, -, NW2
			8'd11 : rdata = 44'b00010010000000101010000000000010100000000000;
			// PEs: 56, 60 -> 61
			// srcs: (329, 7)(805) -9, (154) 0 --> (956) 0:PEGB0, ND1, *, PENB
			8'd12 : rdata = 44'b00011111000000000110000000100000000100000000;
			// PEs: 60, 59 -> 59
			// srcs: (330, 11)(3) 1, (954) -54 --> (1154) -54:NM0, PENB, *, PEGB3
			8'd13 : rdata = 44'b00011100000000001101111111000000000010110000;
			// PEs: 60, 61 -> 60
			// srcs: (338, 14)(355) 3, (1156) 0 --> (1356) 3:NW1, PEGB5, -, NW1
			8'd14 : rdata = 44'b00010010000000011110000101000010010000000000;
			default : rdata = 44'b00000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 61) begin
	always @(*) begin
		case(address)
			// PEs: 61, 61 -> 61
			// srcs: (1, 0)(77) 0, (278) 9 --> (478) 0:ND0, NW0, *, NI0
			8'd0 : rdata = 44'b00011011000000000100000000010000000000000000;
			// PEs: 61, 61 -> 61
			// srcs: (2, 1)(155) 1, (356) 9 --> (556) 9:ND1, NW1, *, NI1
			8'd1 : rdata = 44'b00011011000000010100000000110100000000000000;
			// PEs: 61, 61 -> 56
			// srcs: (3, 2)(85) 9, (286) 8 --> (486) 72:ND2, NW2, *, PEGB0
			8'd2 : rdata = 44'b00011011000000100100000001000000000010000000;
			// PEs: 60, 61 -> 61
			// srcs: (4, 3)(477) 0, (478) 0 --> (673) 0:PENB, NI0, +, NI2
			8'd3 : rdata = 44'b00001110111111101010000000011000000000000000;
			// PEs: 60, 61 -> 62
			// srcs: (5, 4)(555) 0, (556) 9 --> (753) 9:PENB, NI1, +, PENB
			8'd4 : rdata = 44'b00001110111111101010000000100000000100000000;
			// PEs: 61, 60 -> 
			// srcs: (7, 5)(673) 0, (479) 10 --> (674) 10:NI2, PENB, +, 
			8'd5 : rdata = 44'b00001101000000101101111111000000000000000000;
			// PEs: 60, 61 -> 62
			// srcs: (16, 6)(672) 31, (674) 10 --> (675) 41:PENB, ALU, +, PENB
			8'd6 : rdata = 44'b00001110111111100011111111100000000100000000;
			// PEs: 56, 61 -> 62
			// srcs: (252, 7)(805) -9, (77) 0 --> (879) 0:PEGB0, ND0, *, PENB
			8'd7 : rdata = 44'b00011111000000000110000000000000000100000000;
			// PEs: 56, 61 -> 61
			// srcs: (260, 8)(805) -9, (85) 9 --> (887) -81:PEGB0, ND2, *, NI0
			8'd8 : rdata = 44'b00011111000000000110000001010000000000000000;
			// PEs: 61, 62 -> 61
			// srcs: (261, 12)(278) 9, (1079) 0 --> (1279) 9:NW0, PEGB6, -, NW0
			8'd9 : rdata = 44'b00010010000000001110000110000010000000000000;
			// PEs: 61, 61 -> 
			// srcs: (263, 10)(3) 1, (887) -81 --> (1087) -81:NM0, NI0, *, 
			8'd10 : rdata = 44'b00011100000000001010000000000000000000000000;
			// PEs: 61, 61 -> 61
			// srcs: (266, 13)(286) 8, (1087) -81 --> (1287) 89:NW2, ALU, -, NW2
			8'd11 : rdata = 44'b00010010000000100011111111100010100000000000;
			// PEs: 56, 61 -> 62
			// srcs: (330, 9)(805) -9, (155) 1 --> (957) -9:PEGB0, ND1, *, PENB
			8'd12 : rdata = 44'b00011111000000000110000000100000000100000000;
			// PEs: 61, 60 -> 60
			// srcs: (332, 11)(3) 1, (956) 0 --> (1156) 0:NM0, PENB, *, PEGB4
			8'd13 : rdata = 44'b00011100000000001101111111000000000011000000;
			// PEs: 61, 62 -> 61
			// srcs: (339, 14)(356) 9, (1157) -9 --> (1357) 18:NW1, PEGB6, -, NW1
			8'd14 : rdata = 44'b00010010000000011110000110000010010000000000;
			default : rdata = 44'b00000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 62) begin
	always @(*) begin
		case(address)
			// PEs: 62, 62 -> 63
			// srcs: (1, 0)(79) 7, (280) 6 --> (480) 42:ND0, NW0, *, PENB
			8'd0 : rdata = 44'b00011011000000000100000000000000000100000000;
			// PEs: 62, 62 -> 63
			// srcs: (2, 1)(156) 3, (357) 4 --> (557) 12:ND1, NW1, *, PENB
			8'd1 : rdata = 44'b00011011000000010100000000100000000100000000;
			// PEs: 62, 62 -> 56
			// srcs: (3, 2)(88) 4, (289) 8 --> (489) 32:ND2, NW2, *, PEGB0
			8'd2 : rdata = 44'b00011011000000100100000001000000000010000000;
			// PEs: 61, 63 -> 56
			// srcs: (11, 3)(753) 9, (754) 39 --> (755) 48:PENB, PEGB7, +, PEGB0
			8'd3 : rdata = 44'b00001110111111101110000111000000000010000000;
			// PEs: 58, 61 -> 57
			// srcs: (39, 4)(670) 100, (675) 41 --> (676) 141:PEGB2, PENB, +, PEGB1
			8'd4 : rdata = 44'b00001111000001001101111111000000000010010000;
			// PEs: 56, 62 -> 62
			// srcs: (254, 5)(805) -9, (79) 7 --> (881) -63:PEGB0, ND0, *, NI0
			8'd5 : rdata = 44'b00011111000000000110000000010000000000000000;
			// PEs: 62, 61 -> 61
			// srcs: (255, 8)(3) 1, (879) 0 --> (1079) 0:NM0, PENB, *, PEGB5
			8'd6 : rdata = 44'b00011100000000001101111111000000000011010000;
			// PEs: 62, 62 -> 
			// srcs: (257, 9)(3) 1, (881) -63 --> (1081) -63:NM0, NI0, *, 
			8'd7 : rdata = 44'b00011100000000001010000000000000000000000000;
			// PEs: 62, 62 -> 62
			// srcs: (260, 12)(280) 6, (1081) -63 --> (1281) 69:NW0, ALU, -, NW0
			8'd8 : rdata = 44'b00010010000000000011111111100010000000000000;
			// PEs: 56, 62 -> 
			// srcs: (263, 6)(805) -9, (88) 4 --> (890) -36:PEGB0, ND2, *, 
			8'd9 : rdata = 44'b00011111000000000110000001000000000000000000;
			// PEs: 62, 62 -> 
			// srcs: (266, 10)(3) 1, (890) -36 --> (1090) -36:NM0, ALU, *, 
			8'd10 : rdata = 44'b00011100000000000011111111100000000000000000;
			// PEs: 62, 62 -> 62
			// srcs: (269, 13)(289) 8, (1090) -36 --> (1290) 44:NW2, ALU, -, NW2
			8'd11 : rdata = 44'b00010010000000100011111111100010100000000000;
			// PEs: 56, 62 -> 63
			// srcs: (331, 7)(805) -9, (156) 3 --> (958) -27:PEGB0, ND1, *, PENB
			8'd12 : rdata = 44'b00011111000000000110000000100000000100000000;
			// PEs: 62, 61 -> 61
			// srcs: (333, 11)(3) 1, (957) -9 --> (1157) -9:NM0, PENB, *, PEGB5
			8'd13 : rdata = 44'b00011100000000001101111111000000000011010000;
			// PEs: 62, 63 -> 62
			// srcs: (340, 14)(357) 4, (1158) -27 --> (1358) 31:NW1, PEGB7, -, NW1
			8'd14 : rdata = 44'b00010010000000011110000111000010010000000000;
			default : rdata = 44'b00000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 63) begin
	always @(*) begin
		case(address)
			// PEs: 63, 63 -> 63
			// srcs: (1, 0)(80) 5, (281) 4 --> (481) 20:ND0, NW0, *, NI0
			8'd0 : rdata = 44'b00011011000000000100000000010000000000000000;
			// PEs: 63, 63 -> 63
			// srcs: (2, 1)(157) 3, (358) 9 --> (558) 27:ND1, NW1, *, NI1
			8'd1 : rdata = 44'b00011011000000010100000000110100000000000000;
			// PEs: 63, 63 -> 63
			// srcs: (3, 2)(91) 0, (292) 8 --> (492) 0:ND2, NW2, *, NI2
			8'd2 : rdata = 44'b00011011000000100100000001011000000000000000;
			// PEs: 62, 63 -> 56
			// srcs: (4, 3)(480) 42, (481) 20 --> (678) 62:PENB, NI0, +, PENB
			8'd3 : rdata = 44'b00001110111111101010000000000000000100000000;
			// PEs: 62, 63 -> 62
			// srcs: (5, 4)(557) 12, (558) 27 --> (754) 39:PENB, NI1, +, PEGB6
			8'd4 : rdata = 44'b00001110111111101010000000100000000011100000;
			// PEs: 63 -> 56
			// srcs: (12, 5)(492) 0 --> (492) 0:NI2, pass, PENB
			8'd5 : rdata = 44'b11000101000000100000000000000000000100000000;
			// PEs: 56, 63 -> 
			// srcs: (255, 6)(805) -9, (80) 5 --> (882) -45:PEGB0, ND0, *, 
			8'd6 : rdata = 44'b00011111000000000110000000000000000000000000;
			// PEs: 63, 63 -> 
			// srcs: (258, 9)(3) 1, (882) -45 --> (1082) -45:NM0, ALU, *, 
			8'd7 : rdata = 44'b00011100000000000011111111100000000000000000;
			// PEs: 63, 63 -> 63
			// srcs: (261, 13)(281) 4, (1082) -45 --> (1282) 49:NW0, ALU, -, NW0
			8'd8 : rdata = 44'b00010010000000000011111111100010000000000000;
			// PEs: 56, 63 -> 
			// srcs: (266, 7)(805) -9, (91) 0 --> (893) 0:PEGB0, ND2, *, 
			8'd9 : rdata = 44'b00011111000000000110000001000000000000000000;
			// PEs: 63, 63 -> 
			// srcs: (269, 10)(3) 1, (893) 0 --> (1093) 0:NM0, ALU, *, 
			8'd10 : rdata = 44'b00011100000000000011111111100000000000000000;
			// PEs: 63, 63 -> 63
			// srcs: (272, 14)(292) 8, (1093) 0 --> (1293) 8:NW2, ALU, -, NW2
			8'd11 : rdata = 44'b00010010000000100011111111100010100000000000;
			// PEs: 56, 63 -> 63
			// srcs: (332, 8)(805) -9, (157) 3 --> (959) -27:PEGB0, ND1, *, NI0
			8'd12 : rdata = 44'b00011111000000000110000000110000000000000000;
			// PEs: 63, 62 -> 62
			// srcs: (334, 11)(3) 1, (958) -27 --> (1158) -27:NM0, PENB, *, PEGB6
			8'd13 : rdata = 44'b00011100000000001101111111000000000011100000;
			// PEs: 63, 63 -> 
			// srcs: (335, 12)(3) 1, (959) -27 --> (1159) -27:NM0, NI0, *, 
			8'd14 : rdata = 44'b00011100000000001010000000000000000000000000;
			// PEs: 63, 63 -> 63
			// srcs: (338, 15)(358) 9, (1159) -27 --> (1359) 36:NW1, ALU, -, NW1
			8'd15 : rdata = 44'b00010010000000010011111111100010010000000000;
			default : rdata = 44'b00000000000000000000000000000000000000000000;
		endcase
	end
end

endgenerate
/*****************************************************************************/
endmodule
