
`timescale 1ns/1ps
module instruction_memory #(
    parameter integer addrLen = 5,
    parameter integer dataLen = 32,
    parameter integer peId  = 1
)(
    input clk,
    input rstn,
    
    input stall,
    input start,
    input restart,
    
    output reg [dataLen - 1: 0] data_out
);
//--------------------------------------------------------------------------------------
//reg [dataLen - 1: 0] mem  [0: (1 << addrLen) - 1];
reg [addrLen-1:0]        address;
reg enable;
reg [dataLen - 1: 0] rdata;
wire end_of_instruction;
always @(posedge clk or negedge rstn)
    if(~rstn)
        enable <= 1'b0;
    else if(start)
        enable <= 1'b1;
    else if(end_of_instruction)
       enable <= 1'b0;
always @(posedge clk or negedge rstn) begin
    if(~rstn)
        address <= {addrLen{1'b0}};
    else begin
        if(end_of_instruction)
            address <= {addrLen{1'b0}};
        else if(~stall && enable )
            address <= address + {{addrLen-1{1'b0}},1'b1};   
    end     
end
always @(posedge clk or negedge rstn) begin
    if(~rstn)
        data_out <= {1'b1,{dataLen-1{1'b0}}};
    else if((~stall && enable && ~end_of_instruction)||(end_of_instruction && start))
       data_out <= rdata;
end
    
assign end_of_instruction = (data_out[dataLen-1:dataLen-5] == 5'b0);
/****************************************************************************/
generate
if(peId == 0) begin
	always @(*) begin
		case(address)
			// PEs: 7 -> 16
			// srcs: (3, 6)(804) 1395 --> (804) 1395:PENB, pass, PUGB2
			9'd0 : rdata = 43'b1100011011110000000000000000000000000001010;
			// PEs: 7 -> 16
			// srcs: (4, 13)(805) 930 --> (805) 930:PENB, pass, PUGB2
			9'd1 : rdata = 43'b1100011011110000000000000000000000000001010;
			// PEs: 1 -> 24
			// srcs: (6, 0)(624) 84 --> (624) 84:PEGB1, pass, PUGB3
			9'd2 : rdata = 43'b1100011100010000000000000000000000000001011;
			// PEs: 2 -> 24
			// srcs: (7, 1)(654) 11 --> (654) 11:PEGB2, pass, PUGB3
			9'd3 : rdata = 43'b1100011100100000000000000000000000000001011;
			// PEs: 3 -> 32
			// srcs: (8, 2)(684) 1032 --> (684) 1032:PEGB3, pass, PUGB4
			9'd4 : rdata = 43'b1100011100110000000000000000000000000001100;
			// PEs: 4 -> 32
			// srcs: (9, 3)(714) 2116 --> (714) 2116:PEGB4, pass, PUGB4
			9'd5 : rdata = 43'b1100011101000000000000000000000000000001100;
			// PEs: 5 -> 32
			// srcs: (10, 4)(744) 120 --> (744) 120:PEGB5, pass, PUGB4
			9'd6 : rdata = 43'b1100011101010000000000000000000000000001100;
			// PEs: 6 -> 32
			// srcs: (11, 5)(774) 722 --> (774) 722:PEGB6, pass, PUGB4
			9'd7 : rdata = 43'b1100011101100000000000000000000000000001100;
			// PEs: 1 -> 24
			// srcs: (12, 7)(625) 560 --> (625) 560:PEGB1, pass, PUGB3
			9'd8 : rdata = 43'b1100011100010000000000000000000000000001011;
			// PEs: 2 -> 24
			// srcs: (13, 8)(655) 176 --> (655) 176:PEGB2, pass, PUGB3
			9'd9 : rdata = 43'b1100011100100000000000000000000000000001011;
			// PEs: 3 -> 24
			// srcs: (14, 9)(685) 864 --> (685) 864:PEGB3, pass, PUGB3
			9'd10 : rdata = 43'b1100011100110000000000000000000000000001011;
			// PEs: 4 -> 24
			// srcs: (15, 10)(715) 1104 --> (715) 1104:PEGB4, pass, PUGB3
			9'd11 : rdata = 43'b1100011101000000000000000000000000000001011;
			// PEs: 5 -> 24
			// srcs: (16, 11)(745) 1008 --> (745) 1008:PEGB5, pass, PUGB3
			9'd12 : rdata = 43'b1100011101010000000000000000000000000001011;
			// PEs: 6 -> 24
			// srcs: (17, 12)(775) 551 --> (775) 551:PEGB6, pass, PUGB3
			9'd13 : rdata = 43'b1100011101100000000000000000000000000001011;
			// PEs: 1 -> 24
			// srcs: (18, 14)(626) 364 --> (626) 364:PEGB1, pass, PUGB3
			9'd14 : rdata = 43'b1100011100010000000000000000000000000001011;
			// PEs: 2 -> 24
			// srcs: (19, 15)(656) 121 --> (656) 121:PEGB2, pass, PUGB3
			9'd15 : rdata = 43'b1100011100100000000000000000000000000001011;
			// PEs: 3 -> 24
			// srcs: (20, 16)(686) 816 --> (686) 816:PEGB3, pass, PUGB3
			9'd16 : rdata = 43'b1100011100110000000000000000000000000001011;
			// PEs: 4 -> 24
			// srcs: (21, 17)(716) 644 --> (716) 644:PEGB4, pass, PUGB3
			9'd17 : rdata = 43'b1100011101000000000000000000000000000001011;
			// PEs: 5 -> 24
			// srcs: (22, 18)(746) 792 --> (746) 792:PEGB5, pass, PUGB3
			9'd18 : rdata = 43'b1100011101010000000000000000000000000001011;
			// PEs: 6 -> 24
			// srcs: (23, 19)(776) 361 --> (776) 361:PEGB6, pass, PUGB3
			9'd19 : rdata = 43'b1100011101100000000000000000000000000001011;
			// PEs: 7 -> 24
			// srcs: (24, 20)(806) 372 --> (806) 372:PENB, pass, PUGB3
			9'd20 : rdata = 43'b1100011011110000000000000000000000000001011;
			// PEs: 1 -> 32
			// srcs: (25, 21)(627) 238 --> (627) 238:PEGB1, pass, PUGB4
			9'd21 : rdata = 43'b1100011100010000000000000000000000000001100;
			// PEs: 2 -> 32
			// srcs: (26, 22)(657) 66 --> (657) 66:PEGB2, pass, PUGB4
			9'd22 : rdata = 43'b1100011100100000000000000000000000000001100;
			// PEs: 3 -> 32
			// srcs: (27, 23)(687) 168 --> (687) 168:PEGB3, pass, PUGB4
			9'd23 : rdata = 43'b1100011100110000000000000000000000000001100;
			// PEs: 4 -> 32
			// srcs: (28, 24)(717) 598 --> (717) 598:PEGB4, pass, PUGB4
			9'd24 : rdata = 43'b1100011101000000000000000000000000000001100;
			// PEs: 5 -> 32
			// srcs: (29, 25)(747) 864 --> (747) 864:PEGB5, pass, PUGB4
			9'd25 : rdata = 43'b1100011101010000000000000000000000000001100;
			// PEs: 6 -> 32
			// srcs: (30, 26)(777) 703 --> (777) 703:PEGB6, pass, PUGB4
			9'd26 : rdata = 43'b1100011101100000000000000000000000000001100;
			// PEs: 7 -> 40
			// srcs: (31, 27)(807) 310 --> (807) 310:PENB, pass, PUGB5
			9'd27 : rdata = 43'b1100011011110000000000000000000000000001101;
			// PEs: 1 -> 40
			// srcs: (32, 28)(628) 336 --> (628) 336:PEGB1, pass, PUGB5
			9'd28 : rdata = 43'b1100011100010000000000000000000000000001101;
			// PEs: 2 -> 40
			// srcs: (33, 29)(658) 308 --> (658) 308:PEGB2, pass, PUGB5
			9'd29 : rdata = 43'b1100011100100000000000000000000000000001101;
			// PEs: 3 -> 48
			// srcs: (34, 30)(688) 1032 --> (688) 1032:PEGB3, pass, PUGB6
			9'd30 : rdata = 43'b1100011100110000000000000000000000000001110;
			// PEs: 4 -> 48
			// srcs: (35, 31)(718) 1564 --> (718) 1564:PEGB4, pass, PUGB6
			9'd31 : rdata = 43'b1100011101000000000000000000000000000001110;
			// PEs: 5 -> 48
			// srcs: (36, 32)(748) 984 --> (748) 984:PEGB5, pass, PUGB6
			9'd32 : rdata = 43'b1100011101010000000000000000000000000001110;
			// PEs: 6 -> 48
			// srcs: (37, 33)(778) 532 --> (778) 532:PEGB6, pass, PUGB6
			9'd33 : rdata = 43'b1100011101100000000000000000000000000001110;
			// PEs: 7 -> 48
			// srcs: (38, 34)(808) -93 --> (808) -93:PENB, pass, PUGB6
			9'd34 : rdata = 43'b1100011011110000000000000000000000000001110;
			// PEs: 1 -> 56
			// srcs: (39, 35)(629) 630 --> (629) 630:PEGB1, pass, PUGB7
			9'd35 : rdata = 43'b1100011100010000000000000000000000000001111;
			// PEs: 2 -> 56
			// srcs: (40, 36)(659) 22 --> (659) 22:PEGB2, pass, PUGB7
			9'd36 : rdata = 43'b1100011100100000000000000000000000000001111;
			// PEs: 3 -> 56
			// srcs: (41, 37)(689) 600 --> (689) 600:PEGB3, pass, PUGB7
			9'd37 : rdata = 43'b1100011100110000000000000000000000000001111;
			// PEs: 4 -> 56
			// srcs: (42, 38)(719) 1104 --> (719) 1104:PEGB4, pass, PUGB7
			9'd38 : rdata = 43'b1100011101000000000000000000000000000001111;
			// PEs: 5 -> 56
			// srcs: (43, 39)(749) 360 --> (749) 360:PEGB5, pass, PUGB7
			9'd39 : rdata = 43'b1100011101010000000000000000000000000001111;
			// PEs: 6 -> 56
			// srcs: (44, 40)(779) 95 --> (779) 95:PEGB6, pass, PUGB7
			9'd40 : rdata = 43'b1100011101100000000000000000000000000001111;
			// PEs: 7 -> 56
			// srcs: (45, 41)(809) 310 --> (809) 310:PENB, pass, PUGB7
			9'd41 : rdata = 43'b1100011011110000000000000000000000000001111;
			// PEs: 1 -> 32
			// srcs: (46, 42)(630) 252 --> (630) 252:PEGB1, pass, PUGB4
			9'd42 : rdata = 43'b1100011100010000000000000000000000000001100;
			// PEs: 2 -> 32
			// srcs: (47, 43)(660) -22 --> (660) -22:PEGB2, pass, PUGB4
			9'd43 : rdata = 43'b1100011100100000000000000000000000000001100;
			// PEs: 3 -> 32
			// srcs: (48, 44)(690) 192 --> (690) 192:PEGB3, pass, PUGB4
			9'd44 : rdata = 43'b1100011100110000000000000000000000000001100;
			// PEs: 4 -> 32
			// srcs: (49, 45)(720) 1288 --> (720) 1288:PEGB4, pass, PUGB4
			9'd45 : rdata = 43'b1100011101000000000000000000000000000001100;
			// PEs: 5 -> 32
			// srcs: (50, 46)(750) 816 --> (750) 816:PEGB5, pass, PUGB4
			9'd46 : rdata = 43'b1100011101010000000000000000000000000001100;
			// PEs: 6 -> 32
			// srcs: (51, 47)(780) 855 --> (780) 855:PEGB6, pass, PUGB4
			9'd47 : rdata = 43'b1100011101100000000000000000000000000001100;
			// PEs: 7 -> 32
			// srcs: (52, 48)(810) 1178 --> (810) 1178:PENB, pass, PUGB4
			9'd48 : rdata = 43'b1100011011110000000000000000000000000001100;
			// PEs: 1 -> 24
			// srcs: (53, 49)(631) 28 --> (631) 28:PEGB1, pass, PUGB3
			9'd49 : rdata = 43'b1100011100010000000000000000000000000001011;
			// PEs: 2 -> 24
			// srcs: (54, 50)(661) 99 --> (661) 99:PEGB2, pass, PUGB3
			9'd50 : rdata = 43'b1100011100100000000000000000000000000001011;
			// PEs: 3 -> 24
			// srcs: (55, 51)(691) 240 --> (691) 240:PEGB3, pass, PUGB3
			9'd51 : rdata = 43'b1100011100110000000000000000000000000001011;
			// PEs: 4 -> 24
			// srcs: (56, 52)(721) 506 --> (721) 506:PEGB4, pass, PUGB3
			9'd52 : rdata = 43'b1100011101000000000000000000000000000001011;
			// PEs: 5 -> 24
			// srcs: (57, 53)(751) 552 --> (751) 552:PEGB5, pass, PUGB3
			9'd53 : rdata = 43'b1100011101010000000000000000000000000001011;
			// PEs: 6 -> 24
			// srcs: (58, 54)(781) 114 --> (781) 114:PEGB6, pass, PUGB3
			9'd54 : rdata = 43'b1100011101100000000000000000000000000001011;
			// PEs: 7 -> 16
			// srcs: (59, 55)(811) 279 --> (811) 279:PENB, pass, PUGB2
			9'd55 : rdata = 43'b1100011011110000000000000000000000000001010;
			// PEs: 1 -> 40
			// srcs: (60, 56)(632) 112 --> (632) 112:PEGB1, pass, PUGB5
			9'd56 : rdata = 43'b1100011100010000000000000000000000000001101;
			// PEs: 2 -> 40
			// srcs: (61, 57)(662) 264 --> (662) 264:PEGB2, pass, PUGB5
			9'd57 : rdata = 43'b1100011100100000000000000000000000000001101;
			// PEs: 3 -> 40
			// srcs: (62, 58)(692) 456 --> (692) 456:PEGB3, pass, PUGB5
			9'd58 : rdata = 43'b1100011100110000000000000000000000000001101;
			// PEs: 4 -> 40
			// srcs: (63, 59)(722) 1564 --> (722) 1564:PEGB4, pass, PUGB5
			9'd59 : rdata = 43'b1100011101000000000000000000000000000001101;
			// PEs: 5 -> 40
			// srcs: (64, 60)(752) 312 --> (752) 312:PEGB5, pass, PUGB5
			9'd60 : rdata = 43'b1100011101010000000000000000000000000001101;
			// PEs: 6 -> 40
			// srcs: (65, 61)(782) 589 --> (782) 589:PEGB6, pass, PUGB5
			9'd61 : rdata = 43'b1100011101100000000000000000000000000001101;
			// PEs: 7 -> 16
			// srcs: (66, 62)(812) 1457 --> (812) 1457:PENB, pass, PUGB2
			9'd62 : rdata = 43'b1100011011110000000000000000000000000001010;
			// PEs: 1 -> 32
			// srcs: (67, 63)(633) 672 --> (633) 672:PEGB1, pass, PUGB4
			9'd63 : rdata = 43'b1100011100010000000000000000000000000001100;
			// PEs: 2 -> 32
			// srcs: (68, 64)(663) 165 --> (663) 165:PEGB2, pass, PUGB4
			9'd64 : rdata = 43'b1100011100100000000000000000000000000001100;
			// PEs: 3 -> 32
			// srcs: (69, 65)(693) 864 --> (693) 864:PEGB3, pass, PUGB4
			9'd65 : rdata = 43'b1100011100110000000000000000000000000001100;
			// PEs: 4 -> 32
			// srcs: (70, 66)(723) 184 --> (723) 184:PEGB4, pass, PUGB4
			9'd66 : rdata = 43'b1100011101000000000000000000000000000001100;
			// PEs: 5 -> 32
			// srcs: (71, 67)(753) 816 --> (753) 816:PEGB5, pass, PUGB4
			9'd67 : rdata = 43'b1100011101010000000000000000000000000001100;
			// PEs: 6 -> 32
			// srcs: (72, 68)(783) 836 --> (783) 836:PEGB6, pass, PUGB4
			9'd68 : rdata = 43'b1100011101100000000000000000000000000001100;
			// PEs: 7 -> 32
			// srcs: (73, 69)(813) 62 --> (813) 62:PENB, pass, PUGB4
			9'd69 : rdata = 43'b1100011011110000000000000000000000000001100;
			// PEs: 1 -> 40
			// srcs: (74, 70)(634) 448 --> (634) 448:PEGB1, pass, PUGB5
			9'd70 : rdata = 43'b1100011100010000000000000000000000000001101;
			// PEs: 2 -> 40
			// srcs: (75, 71)(664) 528 --> (664) 528:PEGB2, pass, PUGB5
			9'd71 : rdata = 43'b1100011100100000000000000000000000000001101;
			// PEs: 3 -> 40
			// srcs: (76, 72)(694) 960 --> (694) 960:PEGB3, pass, PUGB5
			9'd72 : rdata = 43'b1100011100110000000000000000000000000001101;
			// PEs: 4 -> 40
			// srcs: (77, 73)(724) 874 --> (724) 874:PEGB4, pass, PUGB5
			9'd73 : rdata = 43'b1100011101000000000000000000000000000001101;
			// PEs: 5 -> 40
			// srcs: (78, 74)(754) 1176 --> (754) 1176:PEGB5, pass, PUGB5
			9'd74 : rdata = 43'b1100011101010000000000000000000000000001101;
			// PEs: 6 -> 40
			// srcs: (79, 75)(784) -38 --> (784) -38:PEGB6, pass, PUGB5
			9'd75 : rdata = 43'b1100011101100000000000000000000000000001101;
			// PEs: 7 -> 40
			// srcs: (80, 76)(814) 744 --> (814) 744:PENB, pass, PUGB5
			9'd76 : rdata = 43'b1100011011110000000000000000000000000001101;
			// PEs: 1 -> 48
			// srcs: (81, 77)(635) 434 --> (635) 434:PEGB1, pass, PUGB6
			9'd77 : rdata = 43'b1100011100010000000000000000000000000001110;
			// PEs: 2 -> 48
			// srcs: (82, 78)(665) 429 --> (665) 429:PEGB2, pass, PUGB6
			9'd78 : rdata = 43'b1100011100100000000000000000000000000001110;
			// PEs: 3 -> 48
			// srcs: (83, 79)(695) 336 --> (695) 336:PEGB3, pass, PUGB6
			9'd79 : rdata = 43'b1100011100110000000000000000000000000001110;
			// PEs: 4 -> 48
			// srcs: (84, 80)(725) 184 --> (725) 184:PEGB4, pass, PUGB6
			9'd80 : rdata = 43'b1100011101000000000000000000000000000001110;
			// PEs: 5 -> 48
			// srcs: (85, 81)(755) -24 --> (755) -24:PEGB5, pass, PUGB6
			9'd81 : rdata = 43'b1100011101010000000000000000000000000001110;
			// PEs: 6 -> 48
			// srcs: (86, 82)(785) 304 --> (785) 304:PEGB6, pass, PUGB6
			9'd82 : rdata = 43'b1100011101100000000000000000000000000001110;
			// PEs: 7 -> 56
			// srcs: (87, 83)(815) 1054 --> (815) 1054:PENB, pass, PUGB7
			9'd83 : rdata = 43'b1100011011110000000000000000000000000001111;
			// PEs: 1 -> 56
			// srcs: (88, 84)(636) 140 --> (636) 140:PEGB1, pass, PUGB7
			9'd84 : rdata = 43'b1100011100010000000000000000000000000001111;
			// PEs: 2 -> 56
			// srcs: (89, 85)(666) -22 --> (666) -22:PEGB2, pass, PUGB7
			9'd85 : rdata = 43'b1100011100100000000000000000000000000001111;
			// PEs: 3 -> 24
			// srcs: (90, 86)(696) 792 --> (696) 792:PEGB3, pass, PUGB3
			9'd86 : rdata = 43'b1100011100110000000000000000000000000001011;
			// PEs: 4 -> 24
			// srcs: (91, 87)(726) 1242 --> (726) 1242:PEGB4, pass, PUGB3
			9'd87 : rdata = 43'b1100011101000000000000000000000000000001011;
			// PEs: 5 -> 24
			// srcs: (92, 88)(756) 72 --> (756) 72:PEGB5, pass, PUGB3
			9'd88 : rdata = 43'b1100011101010000000000000000000000000001011;
			// PEs: 6 -> 24
			// srcs: (93, 89)(786) 266 --> (786) 266:PEGB6, pass, PUGB3
			9'd89 : rdata = 43'b1100011101100000000000000000000000000001011;
			// PEs: 7 -> 16
			// srcs: (94, 90)(816) 341 --> (816) 341:PENB, pass, PUGB2
			9'd90 : rdata = 43'b1100011011110000000000000000000000000001010;
			// PEs: 1 -> 24
			// srcs: (95, 91)(637) 84 --> (637) 84:PEGB1, pass, PUGB3
			9'd91 : rdata = 43'b1100011100010000000000000000000000000001011;
			// PEs: 2 -> 24
			// srcs: (96, 92)(667) 0 --> (667) 0:PEGB2, pass, PUGB3
			9'd92 : rdata = 43'b1100011100100000000000000000000000000001011;
			// PEs: 3 -> 24
			// srcs: (97, 93)(697) 1176 --> (697) 1176:PEGB3, pass, PUGB3
			9'd93 : rdata = 43'b1100011100110000000000000000000000000001011;
			// PEs: 4 -> 24
			// srcs: (98, 94)(727) 184 --> (727) 184:PEGB4, pass, PUGB3
			9'd94 : rdata = 43'b1100011101000000000000000000000000000001011;
			// PEs: 5 -> 24
			// srcs: (99, 95)(757) 888 --> (757) 888:PEGB5, pass, PUGB3
			9'd95 : rdata = 43'b1100011101010000000000000000000000000001011;
			// PEs: 6 -> 24
			// srcs: (100, 96)(787) 741 --> (787) 741:PEGB6, pass, PUGB3
			9'd96 : rdata = 43'b1100011101100000000000000000000000000001011;
			// PEs: 7 -> 16
			// srcs: (101, 97)(817) 372 --> (817) 372:PENB, pass, PUGB2
			9'd97 : rdata = 43'b1100011011110000000000000000000000000001010;
			// PEs: 1 -> 32
			// srcs: (102, 98)(638) 28 --> (638) 28:PEGB1, pass, PUGB4
			9'd98 : rdata = 43'b1100011100010000000000000000000000000001100;
			// PEs: 2 -> 32
			// srcs: (103, 99)(668) 264 --> (668) 264:PEGB2, pass, PUGB4
			9'd99 : rdata = 43'b1100011100100000000000000000000000000001100;
			// PEs: 3 -> 32
			// srcs: (104, 100)(698) 432 --> (698) 432:PEGB3, pass, PUGB4
			9'd100 : rdata = 43'b1100011100110000000000000000000000000001100;
			// PEs: 4 -> 32
			// srcs: (105, 101)(728) 966 --> (728) 966:PEGB4, pass, PUGB4
			9'd101 : rdata = 43'b1100011101000000000000000000000000000001100;
			// PEs: 5 -> 32
			// srcs: (106, 102)(758) 936 --> (758) 936:PEGB5, pass, PUGB4
			9'd102 : rdata = 43'b1100011101010000000000000000000000000001100;
			// PEs: 6 -> 32
			// srcs: (107, 103)(788) 399 --> (788) 399:PEGB6, pass, PUGB4
			9'd103 : rdata = 43'b1100011101100000000000000000000000000001100;
			// PEs: 7 -> 32
			// srcs: (108, 104)(818) 837 --> (818) 837:PENB, pass, PUGB4
			9'd104 : rdata = 43'b1100011011110000000000000000000000000001100;
			// PEs: 1 -> 24
			// srcs: (109, 105)(639) 56 --> (639) 56:PEGB1, pass, PUGB3
			9'd105 : rdata = 43'b1100011100010000000000000000000000000001011;
			// PEs: 2 -> 24
			// srcs: (110, 106)(669) 187 --> (669) 187:PEGB2, pass, PUGB3
			9'd106 : rdata = 43'b1100011100100000000000000000000000000001011;
			// PEs: 3 -> 24
			// srcs: (111, 107)(699) 408 --> (699) 408:PEGB3, pass, PUGB3
			9'd107 : rdata = 43'b1100011100110000000000000000000000000001011;
			// PEs: 4 -> 24
			// srcs: (112, 108)(729) 1472 --> (729) 1472:PEGB4, pass, PUGB3
			9'd108 : rdata = 43'b1100011101000000000000000000000000000001011;
			// PEs: 5 -> 24
			// srcs: (113, 109)(759) 840 --> (759) 840:PEGB5, pass, PUGB3
			9'd109 : rdata = 43'b1100011101010000000000000000000000000001011;
			// PEs: 6 -> 24
			// srcs: (114, 110)(789) 532 --> (789) 532:PEGB6, pass, PUGB3
			9'd110 : rdata = 43'b1100011101100000000000000000000000000001011;
			// PEs: 7 -> 32
			// srcs: (115, 111)(819) 868 --> (819) 868:PENB, pass, PUGB4
			9'd111 : rdata = 43'b1100011011110000000000000000000000000001100;
			// PEs: 1 -> 40
			// srcs: (116, 112)(640) -28 --> (640) -28:PEGB1, pass, PUGB5
			9'd112 : rdata = 43'b1100011100010000000000000000000000000001101;
			// PEs: 2 -> 40
			// srcs: (117, 113)(670) 44 --> (670) 44:PEGB2, pass, PUGB5
			9'd113 : rdata = 43'b1100011100100000000000000000000000000001101;
			// PEs: 3 -> 40
			// srcs: (118, 114)(700) 624 --> (700) 624:PEGB3, pass, PUGB5
			9'd114 : rdata = 43'b1100011100110000000000000000000000000001101;
			// PEs: 4 -> 40
			// srcs: (119, 115)(730) 828 --> (730) 828:PEGB4, pass, PUGB5
			9'd115 : rdata = 43'b1100011101000000000000000000000000000001101;
			// PEs: 5 -> 40
			// srcs: (120, 116)(760) 600 --> (760) 600:PEGB5, pass, PUGB5
			9'd116 : rdata = 43'b1100011101010000000000000000000000000001101;
			// PEs: 6 -> 40
			// srcs: (121, 117)(790) 779 --> (790) 779:PEGB6, pass, PUGB5
			9'd117 : rdata = 43'b1100011101100000000000000000000000000001101;
			// PEs: 7 -> 40
			// srcs: (122, 118)(820) 837 --> (820) 837:PENB, pass, PUGB5
			9'd118 : rdata = 43'b1100011011110000000000000000000000000001101;
			// PEs: 1 -> 48
			// srcs: (123, 119)(641) 112 --> (641) 112:PEGB1, pass, PUGB6
			9'd119 : rdata = 43'b1100011100010000000000000000000000000001110;
			// PEs: 2 -> 48
			// srcs: (124, 120)(671) 242 --> (671) 242:PEGB2, pass, PUGB6
			9'd120 : rdata = 43'b1100011100100000000000000000000000000001110;
			// PEs: 3 -> 48
			// srcs: (125, 121)(701) -72 --> (701) -72:PEGB3, pass, PUGB6
			9'd121 : rdata = 43'b1100011100110000000000000000000000000001110;
			// PEs: 4 -> 48
			// srcs: (126, 122)(731) -92 --> (731) -92:PEGB4, pass, PUGB6
			9'd122 : rdata = 43'b1100011101000000000000000000000000000001110;
			// PEs: 5 -> 48
			// srcs: (127, 123)(761) 672 --> (761) 672:PEGB5, pass, PUGB6
			9'd123 : rdata = 43'b1100011101010000000000000000000000000001110;
			// PEs: 6 -> 48
			// srcs: (128, 124)(791) 722 --> (791) 722:PEGB6, pass, PUGB6
			9'd124 : rdata = 43'b1100011101100000000000000000000000000001110;
			// PEs: 7 -> 48
			// srcs: (129, 125)(821) 837 --> (821) 837:PENB, pass, PUGB6
			9'd125 : rdata = 43'b1100011011110000000000000000000000000001110;
			// PEs: 1 -> 56
			// srcs: (130, 126)(642) 238 --> (642) 238:PEGB1, pass, PUGB7
			9'd126 : rdata = 43'b1100011100010000000000000000000000000001111;
			// PEs: 2 -> 56
			// srcs: (131, 127)(672) 506 --> (672) 506:PEGB2, pass, PUGB7
			9'd127 : rdata = 43'b1100011100100000000000000000000000000001111;
			// PEs: 3 -> 56
			// srcs: (132, 128)(702) 864 --> (702) 864:PEGB3, pass, PUGB7
			9'd128 : rdata = 43'b1100011100110000000000000000000000000001111;
			// PEs: 4 -> 56
			// srcs: (133, 129)(732) 1748 --> (732) 1748:PEGB4, pass, PUGB7
			9'd129 : rdata = 43'b1100011101000000000000000000000000000001111;
			// PEs: 5 -> 56
			// srcs: (134, 130)(762) 1056 --> (762) 1056:PEGB5, pass, PUGB7
			9'd130 : rdata = 43'b1100011101010000000000000000000000000001111;
			// PEs: 6 -> 56
			// srcs: (135, 131)(792) 114 --> (792) 114:PEGB6, pass, PUGB7
			9'd131 : rdata = 43'b1100011101100000000000000000000000000001111;
			// PEs: 7 -> 56
			// srcs: (136, 132)(822) 1364 --> (822) 1364:PENB, pass, PUGB7
			9'd132 : rdata = 43'b1100011011110000000000000000000000000001111;
			// PEs: 1 -> 8
			// srcs: (137, 139)(643) 266 --> (643) 266:PEGB1, pass, PUNB
			9'd133 : rdata = 43'b1100011100010000000000000000000001000000000;
			// PEs: 2 -> 8
			// srcs: (138, 140)(673) 143 --> (673) 143:PEGB2, pass, PUNB
			9'd134 : rdata = 43'b1100011100100000000000000000000001000000000;
			// PEs: 3 -> 8
			// srcs: (139, 141)(703) 72 --> (703) 72:PEGB3, pass, PUNB
			9'd135 : rdata = 43'b1100011100110000000000000000000001000000000;
			// PEs: 8 -> 0
			// srcs: (140, 133)(942) 1276 --> (942) 1276:PUGB1, pass, NI0
			9'd136 : rdata = 43'b1100011100011000000001000000000000000000000;
			// PEs: 8 -> 1
			// srcs: (141, 134)(972) 561 --> (972) 561:PUGB1, pass, PENB
			9'd137 : rdata = 43'b1100011100011000000000000000000000100000000;
			// PEs: 4 -> 8
			// srcs: (142, 142)(733) 460 --> (733) 460:PEGB4, pass, PUNB
			9'd138 : rdata = 43'b1100011101000000000000000000000001000000000;
			// PEs: 5 -> 8
			// srcs: (143, 143)(763) -72 --> (763) -72:PEGB5, pass, PUNB
			9'd139 : rdata = 43'b1100011101010000000000000000000001000000000;
			// PEs: 6 -> 8
			// srcs: (144, 144)(793) 95 --> (793) 95:PEGB6, pass, PUNB
			9'd140 : rdata = 43'b1100011101100000000000000000000001000000000;
			// PEs: 7 -> 16
			// srcs: (145, 145)(823) 620 --> (823) 620:PENB, pass, PUGB2
			9'd141 : rdata = 43'b1100011011110000000000000000000000000001010;
			// PEs: 1 -> 8
			// srcs: (146, 146)(644) 210 --> (644) 210:PEGB1, pass, PUNB
			9'd142 : rdata = 43'b1100011100010000000000000000000001000000000;
			// PEs: 0 -> 1
			// srcs: (147, 135)(942) 1276 --> (942) 1276:NI0, pass, PENB
			9'd143 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 8 -> 0
			// srcs: (148, 136)(1002) 42 --> (1002) 42:PUGB1, pass, NI0
			9'd144 : rdata = 43'b1100011100011000000001000000000000000000000;
			// PEs: 8 -> 1
			// srcs: (149, 137)(1032) 594 --> (1032) 594:PUGB1, pass, PENB
			9'd145 : rdata = 43'b1100011100011000000000000000000000100000000;
			// PEs: 2 -> 8
			// srcs: (150, 147)(674) 132 --> (674) 132:PEGB2, pass, PUNB
			9'd146 : rdata = 43'b1100011100100000000000000000000001000000000;
			// PEs: 3 -> 8
			// srcs: (151, 148)(704) 120 --> (704) 120:PEGB3, pass, PUNB
			9'd147 : rdata = 43'b1100011100110000000000000000000001000000000;
			// PEs: 4 -> 8
			// srcs: (152, 149)(734) 46 --> (734) 46:PEGB4, pass, PUNB
			9'd148 : rdata = 43'b1100011101000000000000000000000001000000000;
			// PEs: 5 -> 8
			// srcs: (153, 150)(764) 480 --> (764) 480:PEGB5, pass, PUNB
			9'd149 : rdata = 43'b1100011101010000000000000000000001000000000;
			// PEs: 6 -> 8
			// srcs: (154, 151)(794) 798 --> (794) 798:PEGB6, pass, PUNB
			9'd150 : rdata = 43'b1100011101100000000000000000000001000000000;
			// PEs: 0 -> 1
			// srcs: (155, 138)(1002) 42 --> (1002) 42:NI0, pass, PENB
			9'd151 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 7 -> 8
			// srcs: (156, 152)(824) 713 --> (824) 713:PENB, pass, PUNB
			9'd152 : rdata = 43'b1100011011110000000000000000000001000000000;
			// PEs: 1 -> 8
			// srcs: (157, 153)(645) 98 --> (645) 98:PEGB1, pass, PUNB
			9'd153 : rdata = 43'b1100011100010000000000000000000001000000000;
			// PEs: 2 -> 8
			// srcs: (158, 154)(675) 231 --> (675) 231:PEGB2, pass, PUNB
			9'd154 : rdata = 43'b1100011100100000000000000000000001000000000;
			// PEs: 3 -> 8
			// srcs: (159, 155)(705) 456 --> (705) 456:PEGB3, pass, PUNB
			9'd155 : rdata = 43'b1100011100110000000000000000000001000000000;
			// PEs: 4 -> 8
			// srcs: (160, 156)(735) 1196 --> (735) 1196:PEGB4, pass, PUNB
			9'd156 : rdata = 43'b1100011101000000000000000000000001000000000;
			// PEs: 5 -> 8
			// srcs: (161, 157)(765) 552 --> (765) 552:PEGB5, pass, PUNB
			9'd157 : rdata = 43'b1100011101010000000000000000000001000000000;
			// PEs: 6 -> 8
			// srcs: (162, 158)(795) 209 --> (795) 209:PEGB6, pass, PUNB
			9'd158 : rdata = 43'b1100011101100000000000000000000001000000000;
			// PEs: 7 -> 8
			// srcs: (163, 159)(825) 403 --> (825) 403:PENB, pass, PUNB
			9'd159 : rdata = 43'b1100011011110000000000000000000001000000000;
			// PEs: 1 -> 8
			// srcs: (164, 160)(646) 420 --> (646) 420:PEGB1, pass, PUNB
			9'd160 : rdata = 43'b1100011100010000000000000000000001000000000;
			// PEs: 2 -> 8
			// srcs: (165, 161)(676) 451 --> (676) 451:PEGB2, pass, PUNB
			9'd161 : rdata = 43'b1100011100100000000000000000000001000000000;
			// PEs: 3 -> 8
			// srcs: (166, 162)(706) 576 --> (706) 576:PEGB3, pass, PUNB
			9'd162 : rdata = 43'b1100011100110000000000000000000001000000000;
			// PEs: 4 -> 8
			// srcs: (167, 163)(736) 1196 --> (736) 1196:PEGB4, pass, PUNB
			9'd163 : rdata = 43'b1100011101000000000000000000000001000000000;
			// PEs: 5 -> 8
			// srcs: (168, 164)(766) 504 --> (766) 504:PEGB5, pass, PUNB
			9'd164 : rdata = 43'b1100011101010000000000000000000001000000000;
			// PEs: 6 -> 8
			// srcs: (169, 165)(796) 456 --> (796) 456:PEGB6, pass, PUNB
			9'd165 : rdata = 43'b1100011101100000000000000000000001000000000;
			// PEs: 7 -> 8
			// srcs: (170, 166)(826) 248 --> (826) 248:PENB, pass, PUNB
			9'd166 : rdata = 43'b1100011011110000000000000000000001000000000;
			// PEs: 1 -> 8
			// srcs: (171, 167)(647) 546 --> (647) 546:PEGB1, pass, PUNB
			9'd167 : rdata = 43'b1100011100010000000000000000000001000000000;
			// PEs: 2 -> 8
			// srcs: (172, 168)(677) 121 --> (677) 121:PEGB2, pass, PUNB
			9'd168 : rdata = 43'b1100011100100000000000000000000001000000000;
			// PEs: 3 -> 8
			// srcs: (173, 169)(707) 120 --> (707) 120:PEGB3, pass, PUNB
			9'd169 : rdata = 43'b1100011100110000000000000000000001000000000;
			// PEs: 4 -> 8
			// srcs: (174, 170)(737) 828 --> (737) 828:PEGB4, pass, PUNB
			9'd170 : rdata = 43'b1100011101000000000000000000000001000000000;
			// PEs: 5 -> 8
			// srcs: (175, 171)(767) 672 --> (767) 672:PEGB5, pass, PUNB
			9'd171 : rdata = 43'b1100011101010000000000000000000001000000000;
			// PEs: 6 -> 8
			// srcs: (176, 172)(797) 399 --> (797) 399:PEGB6, pass, PUNB
			9'd172 : rdata = 43'b1100011101100000000000000000000001000000000;
			// PEs: 7 -> 8
			// srcs: (177, 173)(827) 217 --> (827) 217:PENB, pass, PUNB
			9'd173 : rdata = 43'b1100011011110000000000000000000001000000000;
			// PEs: 7 -> 8
			// srcs: (178, 174)(828) 1271 --> (828) 1271:PENB, pass, PUNB
			9'd174 : rdata = 43'b1100011011110000000000000000000001000000000;
			// PEs: 7 -> 8
			// srcs: (179, 175)(829) 992 --> (829) 992:PENB, pass, PUNB
			9'd175 : rdata = 43'b1100011011110000000000000000000001000000000;
			// PEs: 7 -> 8
			// srcs: (180, 176)(830) 806 --> (830) 806:PENB, pass, PUNB
			9'd176 : rdata = 43'b1100011011110000000000000000000001000000000;
			// PEs: 7 -> 8
			// srcs: (181, 177)(831) 744 --> (831) 744:PENB, pass, PUNB
			9'd177 : rdata = 43'b1100011011110000000000000000000001000000000;
			// PEs: 7 -> 8
			// srcs: (182, 178)(832) 341 --> (832) 341:PENB, pass, PUNB
			9'd178 : rdata = 43'b1100011011110000000000000000000001000000000;
			// PEs: 7 -> 8
			// srcs: (183, 179)(833) 465 --> (833) 465:PENB, pass, PUNB
			9'd179 : rdata = 43'b1100011011110000000000000000000001000000000;
			// PEs: 56 -> 0
			// srcs: (184, 180)(1325) 596 --> (1325) 596:PUNB, pass, NI0
			9'd180 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 1 -> 56
			// srcs: (185, 184)(1572) 636 --> (1572) 636:PEGB1, pass, PUGB7
			9'd181 : rdata = 43'b1100011100010000000000000000000000000001111;
			// PEs: 3 -> 8
			// srcs: (186, 185)(1682) 1636 --> (1682) 1636:PEGB3, pass, PUNB
			9'd182 : rdata = 43'b1100011100110000000000000000000001000000000;
			// PEs: 3 -> 24
			// srcs: (187, 186)(1701) 1049 --> (1701) 1049:PEGB3, pass, PUGB3
			9'd183 : rdata = 43'b1100011100110000000000000000000000000001011;
			// PEs: 7 -> 8
			// srcs: (188, 187)(1720) 613 --> (1720) 613:PENB, pass, PUNB
			9'd184 : rdata = 43'b1100011011110000000000000000000001000000000;
			// PEs: 6 -> 32
			// srcs: (189, 188)(1739) 863 --> (1739) 863:PEGB6, pass, PUGB4
			9'd185 : rdata = 43'b1100011101100000000000000000000000000001100;
			// PEs: 2 -> 8
			// srcs: (190, 189)(1758) 1534 --> (1758) 1534:PEGB2, pass, PUNB
			9'd186 : rdata = 43'b1100011100100000000000000000000001000000000;
			// PEs: 6 -> 40
			// srcs: (191, 190)(1777) 1462 --> (1777) 1462:PEGB6, pass, PUGB5
			9'd187 : rdata = 43'b1100011101100000000000000000000000000001101;
			// PEs: 6 -> 8
			// srcs: (192, 193)(1728) 2715 --> (1728) 2715:PEGB6, pass, PUNB
			9'd188 : rdata = 43'b1100011101100000000000000000000001000000000;
			// PEs: 1 -> 32
			// srcs: (199, 191)(1690) 3957 --> (1690) 3957:PEGB1, pass, PUGB4
			9'd189 : rdata = 43'b1100011100010000000000000000000000000001100;
			// PEs: 2 -> 32
			// srcs: (200, 192)(1709) 668 --> (1709) 668:PEGB2, pass, PUGB4
			9'd190 : rdata = 43'b1100011100100000000000000000000000000001100;
			// PEs: 1 -> 8
			// srcs: (201, 195)(1766) 3199 --> (1766) 3199:PEGB1, pass, PUNB
			9'd191 : rdata = 43'b1100011100010000000000000000000001000000000;
			// PEs: 1 -> 32
			// srcs: (208, 194)(1747) 1080 --> (1747) 1080:PEGB1, pass, PUGB4
			9'd192 : rdata = 43'b1100011100010000000000000000000000000001100;
			// PEs: 1 -> 32
			// srcs: (216, 196)(1785) 3847 --> (1785) 3847:PEGB1, pass, PUGB4
			9'd193 : rdata = 43'b1100011100010000000000000000000000000001100;
			// PEs: 16 -> 1
			// srcs: (327, 181)(1326) 1131 --> (1326) 1131:PUGB2, pass, PENB
			9'd194 : rdata = 43'b1100011100101000000000000000000000100000000;
			// PEs: 0 -> 1
			// srcs: (333, 182)(1325) 596 --> (1325) 596:NI0, pass, PENB
			9'd195 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 56 -> 1
			// srcs: (334, 183)(1570) 556 --> (1570) 556:PUNB, pass, PENB
			9'd196 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 56 -> 1
			// srcs: (373, 197)(1331) 2705 --> (1331) 2705:PUNB, pass, PENB
			9'd197 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 1 -> 40
			// srcs: (380, 206)(1335) 4432 --> (1335) 4432:PEGB1, pass, PUGB5
			9'd198 : rdata = 43'b1100011100010000000000000000000000000001101;
			// PEs: 56 -> 1
			// srcs: (470, 198)(1579) 1920 --> (1579) 1920:PUNB, pass, PENB
			9'd199 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 8 -> 0
			// srcs: (471, 199)(1749) 1988 --> (1749) 1988:PUGB1, pass, NI0
			9'd200 : rdata = 43'b1100011100011000000001000000000000000000000;
			// PEs: 16 -> 1
			// srcs: (472, 200)(1750) 917 --> (1750) 917:PUGB2, pass, PENB
			9'd201 : rdata = 43'b1100011100101000000000000000000000100000000;
			// PEs: 0 -> 1
			// srcs: (478, 201)(1749) 1988 --> (1749) 1988:NI0, pass, PENB
			9'd202 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 1 -> 48
			// srcs: (479, 207)(1582) 4313 --> (1582) 4313:PEGB1, pass, PUGB6
			9'd203 : rdata = 43'b1100011100010000000000000000000000000001110;
			// PEs: 1 -> 56
			// srcs: (485, 208)(1753) 2905 --> (1753) 2905:PEGB1, pass, PUGB7
			9'd204 : rdata = 43'b1100011100010000000000000000000000000001111;
			// PEs: 24 -> 0
			// srcs: (558, 202)(1238) 945 --> (1238) 945:PUGB3, pass, NI0
			9'd205 : rdata = 43'b1100011100111000000001000000000000000000000;
			// PEs: 48 -> 1
			// srcs: (559, 203)(1239) 6472 --> (1239) 6472:PUGB6, pass, PENB
			9'd206 : rdata = 43'b1100011101101000000000000000000000100000000;
			// PEs: 0 -> 1
			// srcs: (565, 204)(1238) 945 --> (1238) 945:NI0, pass, PENB
			9'd207 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 1 -> 32
			// srcs: (572, 205)(1241) 7417 --> (1241) 7417:PEGB1, pass, PUGB4
			9'd208 : rdata = 43'b1100011100010000000000000000000000000001100;
			// PEs: 16 -> 0
			// srcs: (1012, 209)(1791) 3445 --> (1791) 3445:PUGB2, pass, NI0
			9'd209 : rdata = 43'b1100011100101000000001000000000000000000000;
			// PEs: 32 -> 1
			// srcs: (1013, 210)(1792) 9011 --> (1792) 9011:PUGB4, pass, PENB
			9'd210 : rdata = 43'b1100011101001000000000000000000000100000000;
			// PEs: 0 -> 1
			// srcs: (1019, 211)(1791) 3445 --> (1791) 3445:NI0, pass, PENB
			9'd211 : rdata = 43'b1100010100000000000000000000000000100000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 1) begin
	always @(*) begin
		case(address)
			// PEs: 1, 1 -> 0
			// srcs: (1, 0)(24) 6, (4) 14 --> (624) 84:NW0, ND0, *, PEGB0
			9'd0 : rdata = 43'b0001101000000011000000000000000000010000000;
			// PEs: 1, 1 -> 0
			// srcs: (2, 1)(25) 40, (4) 14 --> (625) 560:NW1, ND0, *, PEGB0
			9'd1 : rdata = 43'b0001101000001011000000000000000000010000000;
			// PEs: 1, 1 -> 0
			// srcs: (3, 2)(26) 26, (4) 14 --> (626) 364:NW2, ND0, *, PEGB0
			9'd2 : rdata = 43'b0001101000010011000000000000000000010000000;
			// PEs: 1, 1 -> 0
			// srcs: (4, 3)(27) 17, (4) 14 --> (627) 238:NW3, ND0, *, PEGB0
			9'd3 : rdata = 43'b0001101000011011000000000000000000010000000;
			// PEs: 1, 1 -> 0
			// srcs: (5, 4)(28) 24, (4) 14 --> (628) 336:NW4, ND0, *, PEGB0
			9'd4 : rdata = 43'b0001101000100011000000000000000000010000000;
			// PEs: 1, 1 -> 0
			// srcs: (6, 5)(29) 45, (4) 14 --> (629) 630:NW5, ND0, *, PEGB0
			9'd5 : rdata = 43'b0001101000101011000000000000000000010000000;
			// PEs: 1, 1 -> 0
			// srcs: (7, 6)(30) 18, (4) 14 --> (630) 252:NW6, ND0, *, PEGB0
			9'd6 : rdata = 43'b0001101000110011000000000000000000010000000;
			// PEs: 1, 1 -> 0
			// srcs: (8, 7)(31) 2, (4) 14 --> (631) 28:NW7, ND0, *, PEGB0
			9'd7 : rdata = 43'b0001101000111011000000000000000000010000000;
			// PEs: 1, 1 -> 0
			// srcs: (9, 8)(32) 8, (4) 14 --> (632) 112:NW8, ND0, *, PEGB0
			9'd8 : rdata = 43'b0001101001000011000000000000000000010000000;
			// PEs: 1, 1 -> 0
			// srcs: (10, 9)(33) 48, (4) 14 --> (633) 672:NW9, ND0, *, PEGB0
			9'd9 : rdata = 43'b0001101001001011000000000000000000010000000;
			// PEs: 1, 1 -> 0
			// srcs: (11, 10)(34) 32, (4) 14 --> (634) 448:NW10, ND0, *, PEGB0
			9'd10 : rdata = 43'b0001101001010011000000000000000000010000000;
			// PEs: 1, 1 -> 0
			// srcs: (12, 11)(35) 31, (4) 14 --> (635) 434:NW11, ND0, *, PEGB0
			9'd11 : rdata = 43'b0001101001011011000000000000000000010000000;
			// PEs: 1, 1 -> 0
			// srcs: (13, 12)(36) 10, (4) 14 --> (636) 140:NW12, ND0, *, PEGB0
			9'd12 : rdata = 43'b0001101001100011000000000000000000010000000;
			// PEs: 1, 1 -> 0
			// srcs: (14, 13)(37) 6, (4) 14 --> (637) 84:NW13, ND0, *, PEGB0
			9'd13 : rdata = 43'b0001101001101011000000000000000000010000000;
			// PEs: 1, 1 -> 0
			// srcs: (15, 14)(38) 2, (4) 14 --> (638) 28:NW14, ND0, *, PEGB0
			9'd14 : rdata = 43'b0001101001110011000000000000000000010000000;
			// PEs: 1, 1 -> 0
			// srcs: (16, 15)(39) 4, (4) 14 --> (639) 56:NW15, ND0, *, PEGB0
			9'd15 : rdata = 43'b0001101001111011000000000000000000010000000;
			// PEs: 1, 1 -> 0
			// srcs: (17, 16)(40) -2, (4) 14 --> (640) -28:NW16, ND0, *, PEGB0
			9'd16 : rdata = 43'b0001101010000011000000000000000000010000000;
			// PEs: 1, 1 -> 0
			// srcs: (18, 17)(41) 8, (4) 14 --> (641) 112:NW17, ND0, *, PEGB0
			9'd17 : rdata = 43'b0001101010001011000000000000000000010000000;
			// PEs: 1, 1 -> 0
			// srcs: (19, 18)(42) 17, (4) 14 --> (642) 238:NW18, ND0, *, PEGB0
			9'd18 : rdata = 43'b0001101010010011000000000000000000010000000;
			// PEs: 1, 1 -> 0
			// srcs: (20, 19)(43) 19, (4) 14 --> (643) 266:NW19, ND0, *, PEGB0
			9'd19 : rdata = 43'b0001101010011011000000000000000000010000000;
			// PEs: 1, 1 -> 0
			// srcs: (21, 20)(44) 15, (4) 14 --> (644) 210:NW20, ND0, *, PEGB0
			9'd20 : rdata = 43'b0001101010100011000000000000000000010000000;
			// PEs: 1, 1 -> 0
			// srcs: (22, 21)(45) 7, (4) 14 --> (645) 98:NW21, ND0, *, PEGB0
			9'd21 : rdata = 43'b0001101010101011000000000000000000010000000;
			// PEs: 1, 1 -> 0
			// srcs: (23, 22)(46) 30, (4) 14 --> (646) 420:NW22, ND0, *, PEGB0
			9'd22 : rdata = 43'b0001101010110011000000000000000000010000000;
			// PEs: 1, 1 -> 0
			// srcs: (24, 23)(47) 39, (4) 14 --> (647) 546:NW23, ND0, *, PEGB0
			9'd23 : rdata = 43'b0001101010111011000000000000000000010000000;
			// PEs: 1, 1 -> 1
			// srcs: (25, 24)(48) 32, (4) 14 --> (648) 448:NW24, ND0, *, NI0
			9'd24 : rdata = 43'b0001101011000011000001000000000000000000000;
			// PEs: 1, 1 -> 1
			// srcs: (26, 25)(49) 2, (4) 14 --> (649) 28:NW25, ND0, *, NI1
			9'd25 : rdata = 43'b0001101011001011000001000010000000000000000;
			// PEs: 1, 1 -> 5
			// srcs: (27, 26)(50) 27, (4) 14 --> (650) 378:NW26, ND0, *, PEGB5
			9'd26 : rdata = 43'b0001101011010011000000000000000000011010000;
			// PEs: 1, 1 -> 1
			// srcs: (28, 27)(51) 24, (4) 14 --> (651) 336:NW27, ND0, *, NI2
			9'd27 : rdata = 43'b0001101011011011000001000100000000000000000;
			// PEs: 1, 1 -> 1
			// srcs: (29, 28)(52) 32, (4) 14 --> (652) 448:NW28, ND0, *, NI3
			9'd28 : rdata = 43'b0001101011100011000001000110000000000000000;
			// PEs: 1, 1 -> 1
			// srcs: (30, 29)(53) 33, (4) 14 --> (653) 462:NW29, ND0, *, NI4
			9'd29 : rdata = 43'b0001101011101011000001001000000000000000000;
			// PEs: 1, 2 -> 1
			// srcs: (31, 34)(648) 448, (678) 429 --> (1680) 877:NI0, PEGB2, +, NI5
			9'd30 : rdata = 43'b0000110100000111001001001010000000000000000;
			// PEs: 1, 2 -> 2
			// srcs: (32, 35)(649) 28, (679) 352 --> (1699) 380:NI1, PEGB2, +, PENB
			9'd31 : rdata = 43'b0000110100001111001000000000000000100000000;
			// PEs: 1, 2 -> 1
			// srcs: (34, 36)(651) 336, (681) -22 --> (1737) 314:NI2, PEGB2, +, NI0
			9'd32 : rdata = 43'b0000110100010111001001000000000000000000000;
			// PEs: 1, 2 -> 1
			// srcs: (35, 37)(652) 448, (682) 253 --> (1756) 701:NI3, PEGB2, +, NI1
			9'd33 : rdata = 43'b0000110100011111001001000010000000000000000;
			// PEs: 1, 2 -> 1
			// srcs: (36, 38)(653) 462, (683) 165 --> (1775) 627:NI4, PEGB2, +, NI2
			9'd34 : rdata = 43'b0000110100100111001001000100000000000000000;
			// PEs: 1, 2 -> 1
			// srcs: (39, 42)(1680) 877, (1681) 3080 --> (1690) 3957:NI5, PEGB2, +, NI3
			9'd35 : rdata = 43'b0000110100101111001001000110000000000000000;
			// PEs: 1, 4 -> 1
			// srcs: (40, 43)(1737) 314, (1738) 766 --> (1747) 1080:NI0, PEGB4, +, NI4
			9'd36 : rdata = 43'b0000110100000111010001001000000000000000000;
			// PEs: 1, 4 -> 1
			// srcs: (41, 44)(1756) 701, (1757) 2498 --> (1766) 3199:NI1, PEGB4, +, NI0
			9'd37 : rdata = 43'b0000110100001111010001000000000000000000000;
			// PEs: 1, 4 -> 1
			// srcs: (42, 45)(1775) 627, (1776) 3220 --> (1785) 3847:NI2, PEGB4, +, NI1
			9'd38 : rdata = 43'b0000110100010111010001000010000000000000000;
			// PEs: 0 -> 
			// srcs: (143, 30)(972) 561 --> (972) 561:PENB, pass, 
			9'd39 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 0, 1 -> 1
			// srcs: (149, 31)(942) 1276, (972) 561 --> (1571) 1837:PENB, ALU, +, NI2
			9'd40 : rdata = 43'b0000111011110001111111000100000000000000000;
			// PEs: 0 -> 
			// srcs: (151, 32)(1032) 594 --> (1032) 594:PENB, pass, 
			9'd41 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 0, 1 -> 0
			// srcs: (157, 33)(1002) 42, (1032) 594 --> (1572) 636:PENB, ALU, +, PEGB0
			9'd42 : rdata = 43'b0000111011110001111110000000000000010000000;
			// PEs: 1 -> 0
			// srcs: (194, 46)(1690) 3957 --> (1690) 3957:NI3, pass, PEGB0
			9'd43 : rdata = 43'b1100010100011000000000000000000000010000000;
			// PEs: 1 -> 0
			// srcs: (195, 48)(1766) 3199 --> (1766) 3199:NI0, pass, PEGB0
			9'd44 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 1 -> 0
			// srcs: (203, 47)(1747) 1080 --> (1747) 1080:NI4, pass, PEGB0
			9'd45 : rdata = 43'b1100010100100000000000000000000000010000000;
			// PEs: 1 -> 0
			// srcs: (211, 49)(1785) 3847 --> (1785) 3847:NI1, pass, PEGB0
			9'd46 : rdata = 43'b1100010100001000000000000000000000010000000;
			// PEs: 0 -> 
			// srcs: (329, 39)(1326) 1131 --> (1326) 1131:PENB, pass, 
			9'd47 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 0, 1 -> 1
			// srcs: (335, 40)(1325) 596, (1326) 1131 --> (1332) 1727:PENB, ALU, +, NI0
			9'd48 : rdata = 43'b0000111011110001111111000000000000000000000;
			// PEs: 0, 1 -> 1
			// srcs: (336, 41)(1570) 556, (1571) 1837 --> (1578) 2393:PENB, NI2, +, NI1
			9'd49 : rdata = 43'b0000111011110101000101000010000000000000000;
			// PEs: 0, 1 -> 0
			// srcs: (375, 50)(1331) 2705, (1332) 1727 --> (1335) 4432:PENB, NI0, +, PEGB0
			9'd50 : rdata = 43'b0000111011110101000000000000000000010000000;
			// PEs: 1, 0 -> 0
			// srcs: (473, 51)(1578) 2393, (1579) 1920 --> (1582) 4313:NI1, PENB, +, PEGB0
			9'd51 : rdata = 43'b0000110100001110111100000000000000010000000;
			// PEs: 0 -> 
			// srcs: (474, 52)(1750) 917 --> (1750) 917:PENB, pass, 
			9'd52 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 0, 1 -> 0
			// srcs: (480, 53)(1749) 1988, (1750) 917 --> (1753) 2905:PENB, ALU, +, PEGB0
			9'd53 : rdata = 43'b0000111011110001111110000000000000010000000;
			// PEs: 0 -> 
			// srcs: (561, 54)(1239) 6472 --> (1239) 6472:PENB, pass, 
			9'd54 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 0, 1 -> 0
			// srcs: (567, 55)(1238) 945, (1239) 6472 --> (1241) 7417:PENB, ALU, +, PEGB0
			9'd55 : rdata = 43'b0000111011110001111110000000000000010000000;
			// PEs: 0 -> 
			// srcs: (1015, 56)(1792) 9011 --> (1792) 9011:PENB, pass, 
			9'd56 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 0, 1 -> 1
			// srcs: (1021, 57)(1791) 3445, (1792) 9011 --> (1793) 12456:PENB, ALU, +, NW30
			9'd57 : rdata = 43'b0000111011110001111110000001111100000000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 2) begin
	always @(*) begin
		case(address)
			// PEs: 2, 2 -> 0
			// srcs: (1, 0)(54) 1, (5) 11 --> (654) 11:NW0, ND0, *, PEGB0
			9'd0 : rdata = 43'b0001101000000011000000000000000000010000000;
			// PEs: 2, 2 -> 0
			// srcs: (2, 1)(55) 16, (5) 11 --> (655) 176:NW1, ND0, *, PEGB0
			9'd1 : rdata = 43'b0001101000001011000000000000000000010000000;
			// PEs: 2, 2 -> 0
			// srcs: (3, 2)(56) 11, (5) 11 --> (656) 121:NW2, ND0, *, PEGB0
			9'd2 : rdata = 43'b0001101000010011000000000000000000010000000;
			// PEs: 2, 2 -> 0
			// srcs: (4, 3)(57) 6, (5) 11 --> (657) 66:NW3, ND0, *, PEGB0
			9'd3 : rdata = 43'b0001101000011011000000000000000000010000000;
			// PEs: 2, 2 -> 0
			// srcs: (5, 4)(58) 28, (5) 11 --> (658) 308:NW4, ND0, *, PEGB0
			9'd4 : rdata = 43'b0001101000100011000000000000000000010000000;
			// PEs: 2, 2 -> 0
			// srcs: (6, 5)(59) 2, (5) 11 --> (659) 22:NW5, ND0, *, PEGB0
			9'd5 : rdata = 43'b0001101000101011000000000000000000010000000;
			// PEs: 2, 2 -> 0
			// srcs: (7, 6)(60) -2, (5) 11 --> (660) -22:NW6, ND0, *, PEGB0
			9'd6 : rdata = 43'b0001101000110011000000000000000000010000000;
			// PEs: 2, 2 -> 0
			// srcs: (8, 7)(61) 9, (5) 11 --> (661) 99:NW7, ND0, *, PEGB0
			9'd7 : rdata = 43'b0001101000111011000000000000000000010000000;
			// PEs: 2, 2 -> 0
			// srcs: (9, 8)(62) 24, (5) 11 --> (662) 264:NW8, ND0, *, PEGB0
			9'd8 : rdata = 43'b0001101001000011000000000000000000010000000;
			// PEs: 2, 2 -> 0
			// srcs: (10, 9)(63) 15, (5) 11 --> (663) 165:NW9, ND0, *, PEGB0
			9'd9 : rdata = 43'b0001101001001011000000000000000000010000000;
			// PEs: 2, 2 -> 0
			// srcs: (11, 10)(64) 48, (5) 11 --> (664) 528:NW10, ND0, *, PEGB0
			9'd10 : rdata = 43'b0001101001010011000000000000000000010000000;
			// PEs: 2, 2 -> 0
			// srcs: (12, 11)(65) 39, (5) 11 --> (665) 429:NW11, ND0, *, PEGB0
			9'd11 : rdata = 43'b0001101001011011000000000000000000010000000;
			// PEs: 2, 2 -> 0
			// srcs: (13, 12)(66) -2, (5) 11 --> (666) -22:NW12, ND0, *, PEGB0
			9'd12 : rdata = 43'b0001101001100011000000000000000000010000000;
			// PEs: 2, 2 -> 0
			// srcs: (14, 13)(67) 0, (5) 11 --> (667) 0:NW13, ND0, *, PEGB0
			9'd13 : rdata = 43'b0001101001101011000000000000000000010000000;
			// PEs: 2, 2 -> 0
			// srcs: (15, 14)(68) 24, (5) 11 --> (668) 264:NW14, ND0, *, PEGB0
			9'd14 : rdata = 43'b0001101001110011000000000000000000010000000;
			// PEs: 2, 2 -> 0
			// srcs: (16, 15)(69) 17, (5) 11 --> (669) 187:NW15, ND0, *, PEGB0
			9'd15 : rdata = 43'b0001101001111011000000000000000000010000000;
			// PEs: 2, 2 -> 0
			// srcs: (17, 16)(70) 4, (5) 11 --> (670) 44:NW16, ND0, *, PEGB0
			9'd16 : rdata = 43'b0001101010000011000000000000000000010000000;
			// PEs: 2, 2 -> 0
			// srcs: (18, 17)(71) 22, (5) 11 --> (671) 242:NW17, ND0, *, PEGB0
			9'd17 : rdata = 43'b0001101010001011000000000000000000010000000;
			// PEs: 2, 2 -> 0
			// srcs: (19, 18)(72) 46, (5) 11 --> (672) 506:NW18, ND0, *, PEGB0
			9'd18 : rdata = 43'b0001101010010011000000000000000000010000000;
			// PEs: 2, 2 -> 0
			// srcs: (20, 19)(73) 13, (5) 11 --> (673) 143:NW19, ND0, *, PEGB0
			9'd19 : rdata = 43'b0001101010011011000000000000000000010000000;
			// PEs: 2, 2 -> 0
			// srcs: (21, 20)(74) 12, (5) 11 --> (674) 132:NW20, ND0, *, PEGB0
			9'd20 : rdata = 43'b0001101010100011000000000000000000010000000;
			// PEs: 2, 2 -> 0
			// srcs: (22, 21)(75) 21, (5) 11 --> (675) 231:NW21, ND0, *, PEGB0
			9'd21 : rdata = 43'b0001101010101011000000000000000000010000000;
			// PEs: 2, 2 -> 0
			// srcs: (23, 22)(76) 41, (5) 11 --> (676) 451:NW22, ND0, *, PEGB0
			9'd22 : rdata = 43'b0001101010110011000000000000000000010000000;
			// PEs: 2, 2 -> 0
			// srcs: (24, 23)(77) 11, (5) 11 --> (677) 121:NW23, ND0, *, PEGB0
			9'd23 : rdata = 43'b0001101010111011000000000000000000010000000;
			// PEs: 2, 2 -> 1
			// srcs: (25, 24)(78) 39, (5) 11 --> (678) 429:NW24, ND0, *, PEGB1
			9'd24 : rdata = 43'b0001101011000011000000000000000000010010000;
			// PEs: 2, 2 -> 1
			// srcs: (26, 25)(79) 32, (5) 11 --> (679) 352:NW25, ND0, *, PEGB1
			9'd25 : rdata = 43'b0001101011001011000000000000000000010010000;
			// PEs: 2, 2 -> 5
			// srcs: (27, 26)(80) 43, (5) 11 --> (680) 473:NW26, ND0, *, PEGB5
			9'd26 : rdata = 43'b0001101011010011000000000000000000011010000;
			// PEs: 2, 2 -> 1
			// srcs: (28, 27)(81) -2, (5) 11 --> (681) -22:NW27, ND0, *, PEGB1
			9'd27 : rdata = 43'b0001101011011011000000000000000000010010000;
			// PEs: 2, 2 -> 1
			// srcs: (29, 28)(82) 23, (5) 11 --> (682) 253:NW28, ND0, *, PEGB1
			9'd28 : rdata = 43'b0001101011100011000000000000000000010010000;
			// PEs: 2, 2 -> 1
			// srcs: (30, 29)(83) 15, (5) 11 --> (683) 165:NW29, ND0, *, PEGB1
			9'd29 : rdata = 43'b0001101011101011000000000000000000010010000;
			// PEs: 4 -> 2
			// srcs: (31, 30)(738) 2024 --> (738) 2024:PEGB4, pass, NI0
			9'd30 : rdata = 43'b1100011101000000000001000000000000000000000;
			// PEs: 4 -> 2
			// srcs: (32, 32)(739) 0 --> (739) 0:PEGB4, pass, NI1
			9'd31 : rdata = 43'b1100011101000000000001000010000000000000000;
			// PEs: 3, 2 -> 1
			// srcs: (33, 31)(708) 1056, (738) 2024 --> (1681) 3080:PEGB3, NI0, +, PEGB1
			9'd32 : rdata = 43'b0000111100110101000000000000000000010010000;
			// PEs: 6 -> 2
			// srcs: (34, 34)(802) 646 --> (802) 646:PEGB6, pass, NI0
			9'd33 : rdata = 43'b1100011101100000000001000000000000000000000;
			// PEs: 3, 2 -> 2
			// srcs: (36, 33)(709) 288, (739) 0 --> (1700) 288:PEGB3, NI1, +, NI2
			9'd34 : rdata = 43'b0000111100110101000011000100000000000000000;
			// PEs: 5, 2 -> 0
			// srcs: (37, 35)(772) 888, (802) 646 --> (1758) 1534:PEGB5, NI0, +, PEGB0
			9'd35 : rdata = 43'b0000111101010101000000000000000000010000000;
			// PEs: 1, 2 -> 0
			// srcs: (39, 36)(1699) 380, (1700) 288 --> (1709) 668:PENB, NI2, +, PEGB0
			9'd36 : rdata = 43'b0000111011110101000100000000000000010000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 3) begin
	always @(*) begin
		case(address)
			// PEs: 3, 3 -> 0
			// srcs: (1, 0)(84) 43, (6) 24 --> (684) 1032:NW0, ND0, *, PEGB0
			9'd0 : rdata = 43'b0001101000000011000000000000000000010000000;
			// PEs: 3, 3 -> 0
			// srcs: (2, 1)(85) 36, (6) 24 --> (685) 864:NW1, ND0, *, PEGB0
			9'd1 : rdata = 43'b0001101000001011000000000000000000010000000;
			// PEs: 3, 3 -> 0
			// srcs: (3, 2)(86) 34, (6) 24 --> (686) 816:NW2, ND0, *, PEGB0
			9'd2 : rdata = 43'b0001101000010011000000000000000000010000000;
			// PEs: 3, 3 -> 0
			// srcs: (4, 3)(87) 7, (6) 24 --> (687) 168:NW3, ND0, *, PEGB0
			9'd3 : rdata = 43'b0001101000011011000000000000000000010000000;
			// PEs: 3, 3 -> 0
			// srcs: (5, 4)(88) 43, (6) 24 --> (688) 1032:NW4, ND0, *, PEGB0
			9'd4 : rdata = 43'b0001101000100011000000000000000000010000000;
			// PEs: 3, 3 -> 0
			// srcs: (6, 5)(89) 25, (6) 24 --> (689) 600:NW5, ND0, *, PEGB0
			9'd5 : rdata = 43'b0001101000101011000000000000000000010000000;
			// PEs: 3, 3 -> 0
			// srcs: (7, 6)(90) 8, (6) 24 --> (690) 192:NW6, ND0, *, PEGB0
			9'd6 : rdata = 43'b0001101000110011000000000000000000010000000;
			// PEs: 3, 3 -> 0
			// srcs: (8, 7)(91) 10, (6) 24 --> (691) 240:NW7, ND0, *, PEGB0
			9'd7 : rdata = 43'b0001101000111011000000000000000000010000000;
			// PEs: 3, 3 -> 0
			// srcs: (9, 8)(92) 19, (6) 24 --> (692) 456:NW8, ND0, *, PEGB0
			9'd8 : rdata = 43'b0001101001000011000000000000000000010000000;
			// PEs: 3, 3 -> 0
			// srcs: (10, 9)(93) 36, (6) 24 --> (693) 864:NW9, ND0, *, PEGB0
			9'd9 : rdata = 43'b0001101001001011000000000000000000010000000;
			// PEs: 3, 3 -> 0
			// srcs: (11, 10)(94) 40, (6) 24 --> (694) 960:NW10, ND0, *, PEGB0
			9'd10 : rdata = 43'b0001101001010011000000000000000000010000000;
			// PEs: 3, 3 -> 0
			// srcs: (12, 11)(95) 14, (6) 24 --> (695) 336:NW11, ND0, *, PEGB0
			9'd11 : rdata = 43'b0001101001011011000000000000000000010000000;
			// PEs: 3, 3 -> 0
			// srcs: (13, 12)(96) 33, (6) 24 --> (696) 792:NW12, ND0, *, PEGB0
			9'd12 : rdata = 43'b0001101001100011000000000000000000010000000;
			// PEs: 3, 3 -> 0
			// srcs: (14, 13)(97) 49, (6) 24 --> (697) 1176:NW13, ND0, *, PEGB0
			9'd13 : rdata = 43'b0001101001101011000000000000000000010000000;
			// PEs: 3, 3 -> 0
			// srcs: (15, 14)(98) 18, (6) 24 --> (698) 432:NW14, ND0, *, PEGB0
			9'd14 : rdata = 43'b0001101001110011000000000000000000010000000;
			// PEs: 3, 3 -> 0
			// srcs: (16, 15)(99) 17, (6) 24 --> (699) 408:NW15, ND0, *, PEGB0
			9'd15 : rdata = 43'b0001101001111011000000000000000000010000000;
			// PEs: 3, 3 -> 0
			// srcs: (17, 16)(100) 26, (6) 24 --> (700) 624:NW16, ND0, *, PEGB0
			9'd16 : rdata = 43'b0001101010000011000000000000000000010000000;
			// PEs: 3, 3 -> 0
			// srcs: (18, 17)(101) -3, (6) 24 --> (701) -72:NW17, ND0, *, PEGB0
			9'd17 : rdata = 43'b0001101010001011000000000000000000010000000;
			// PEs: 3, 3 -> 0
			// srcs: (19, 18)(102) 36, (6) 24 --> (702) 864:NW18, ND0, *, PEGB0
			9'd18 : rdata = 43'b0001101010010011000000000000000000010000000;
			// PEs: 3, 3 -> 0
			// srcs: (20, 19)(103) 3, (6) 24 --> (703) 72:NW19, ND0, *, PEGB0
			9'd19 : rdata = 43'b0001101010011011000000000000000000010000000;
			// PEs: 3, 3 -> 0
			// srcs: (21, 20)(104) 5, (6) 24 --> (704) 120:NW20, ND0, *, PEGB0
			9'd20 : rdata = 43'b0001101010100011000000000000000000010000000;
			// PEs: 3, 3 -> 0
			// srcs: (22, 21)(105) 19, (6) 24 --> (705) 456:NW21, ND0, *, PEGB0
			9'd21 : rdata = 43'b0001101010101011000000000000000000010000000;
			// PEs: 3, 3 -> 0
			// srcs: (23, 22)(106) 24, (6) 24 --> (706) 576:NW22, ND0, *, PEGB0
			9'd22 : rdata = 43'b0001101010110011000000000000000000010000000;
			// PEs: 3, 3 -> 0
			// srcs: (24, 23)(107) 5, (6) 24 --> (707) 120:NW23, ND0, *, PEGB0
			9'd23 : rdata = 43'b0001101010111011000000000000000000010000000;
			// PEs: 3, 3 -> 2
			// srcs: (25, 24)(108) 44, (6) 24 --> (708) 1056:NW24, ND0, *, PEGB2
			9'd24 : rdata = 43'b0001101011000011000000000000000000010100000;
			// PEs: 3, 3 -> 2
			// srcs: (26, 25)(109) 12, (6) 24 --> (709) 288:NW25, ND0, *, PEGB2
			9'd25 : rdata = 43'b0001101011001011000000000000000000010100000;
			// PEs: 3, 3 -> 6
			// srcs: (27, 26)(110) 47, (6) 24 --> (710) 1128:NW26, ND0, *, PEGB6
			9'd26 : rdata = 43'b0001101011010011000000000000000000011100000;
			// PEs: 3, 3 -> 4
			// srcs: (28, 27)(111) 7, (6) 24 --> (711) 168:NW27, ND0, *, PENB
			9'd27 : rdata = 43'b0001101011011011000000000000000000100000000;
			// PEs: 3, 3 -> 4
			// srcs: (29, 28)(112) 37, (6) 24 --> (712) 888:NW28, ND0, *, PENB
			9'd28 : rdata = 43'b0001101011100011000000000000000000100000000;
			// PEs: 3, 3 -> 4
			// srcs: (30, 29)(113) 46, (6) 24 --> (713) 1104:NW29, ND0, *, PENB
			9'd29 : rdata = 43'b0001101011101011000000000000000000100000000;
			// PEs: 6 -> 3
			// srcs: (31, 30)(798) 532 --> (798) 532:PEGB6, pass, NI0
			9'd30 : rdata = 43'b1100011101100000000001000000000000000000000;
			// PEs: 6 -> 3
			// srcs: (32, 32)(799) 665 --> (799) 665:PEGB6, pass, NI1
			9'd31 : rdata = 43'b1100011101100000000001000010000000000000000;
			// PEs: 5, 3 -> 0
			// srcs: (33, 31)(768) 1104, (798) 532 --> (1682) 1636:PEGB5, NI0, +, PEGB0
			9'd32 : rdata = 43'b0000111101010101000000000000000000010000000;
			// PEs: 5, 3 -> 0
			// srcs: (36, 33)(769) 384, (799) 665 --> (1701) 1049:PEGB5, NI1, +, PEGB0
			9'd33 : rdata = 43'b0000111101010101000010000000000000010000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 4) begin
	always @(*) begin
		case(address)
			// PEs: 4, 4 -> 0
			// srcs: (1, 0)(114) 46, (7) 46 --> (714) 2116:NW0, ND0, *, PEGB0
			9'd0 : rdata = 43'b0001101000000011000000000000000000010000000;
			// PEs: 4, 4 -> 0
			// srcs: (2, 1)(115) 24, (7) 46 --> (715) 1104:NW1, ND0, *, PEGB0
			9'd1 : rdata = 43'b0001101000001011000000000000000000010000000;
			// PEs: 4, 4 -> 0
			// srcs: (3, 2)(116) 14, (7) 46 --> (716) 644:NW2, ND0, *, PEGB0
			9'd2 : rdata = 43'b0001101000010011000000000000000000010000000;
			// PEs: 4, 4 -> 0
			// srcs: (4, 3)(117) 13, (7) 46 --> (717) 598:NW3, ND0, *, PEGB0
			9'd3 : rdata = 43'b0001101000011011000000000000000000010000000;
			// PEs: 4, 4 -> 0
			// srcs: (5, 4)(118) 34, (7) 46 --> (718) 1564:NW4, ND0, *, PEGB0
			9'd4 : rdata = 43'b0001101000100011000000000000000000010000000;
			// PEs: 4, 4 -> 0
			// srcs: (6, 5)(119) 24, (7) 46 --> (719) 1104:NW5, ND0, *, PEGB0
			9'd5 : rdata = 43'b0001101000101011000000000000000000010000000;
			// PEs: 4, 4 -> 0
			// srcs: (7, 6)(120) 28, (7) 46 --> (720) 1288:NW6, ND0, *, PEGB0
			9'd6 : rdata = 43'b0001101000110011000000000000000000010000000;
			// PEs: 4, 4 -> 0
			// srcs: (8, 7)(121) 11, (7) 46 --> (721) 506:NW7, ND0, *, PEGB0
			9'd7 : rdata = 43'b0001101000111011000000000000000000010000000;
			// PEs: 4, 4 -> 0
			// srcs: (9, 8)(122) 34, (7) 46 --> (722) 1564:NW8, ND0, *, PEGB0
			9'd8 : rdata = 43'b0001101001000011000000000000000000010000000;
			// PEs: 4, 4 -> 0
			// srcs: (10, 9)(123) 4, (7) 46 --> (723) 184:NW9, ND0, *, PEGB0
			9'd9 : rdata = 43'b0001101001001011000000000000000000010000000;
			// PEs: 4, 4 -> 0
			// srcs: (11, 10)(124) 19, (7) 46 --> (724) 874:NW10, ND0, *, PEGB0
			9'd10 : rdata = 43'b0001101001010011000000000000000000010000000;
			// PEs: 4, 4 -> 0
			// srcs: (12, 11)(125) 4, (7) 46 --> (725) 184:NW11, ND0, *, PEGB0
			9'd11 : rdata = 43'b0001101001011011000000000000000000010000000;
			// PEs: 4, 4 -> 0
			// srcs: (13, 12)(126) 27, (7) 46 --> (726) 1242:NW12, ND0, *, PEGB0
			9'd12 : rdata = 43'b0001101001100011000000000000000000010000000;
			// PEs: 4, 4 -> 0
			// srcs: (14, 13)(127) 4, (7) 46 --> (727) 184:NW13, ND0, *, PEGB0
			9'd13 : rdata = 43'b0001101001101011000000000000000000010000000;
			// PEs: 4, 4 -> 0
			// srcs: (15, 14)(128) 21, (7) 46 --> (728) 966:NW14, ND0, *, PEGB0
			9'd14 : rdata = 43'b0001101001110011000000000000000000010000000;
			// PEs: 4, 4 -> 0
			// srcs: (16, 15)(129) 32, (7) 46 --> (729) 1472:NW15, ND0, *, PEGB0
			9'd15 : rdata = 43'b0001101001111011000000000000000000010000000;
			// PEs: 4, 4 -> 0
			// srcs: (17, 16)(130) 18, (7) 46 --> (730) 828:NW16, ND0, *, PEGB0
			9'd16 : rdata = 43'b0001101010000011000000000000000000010000000;
			// PEs: 4, 4 -> 0
			// srcs: (18, 17)(131) -2, (7) 46 --> (731) -92:NW17, ND0, *, PEGB0
			9'd17 : rdata = 43'b0001101010001011000000000000000000010000000;
			// PEs: 4, 4 -> 0
			// srcs: (19, 18)(132) 38, (7) 46 --> (732) 1748:NW18, ND0, *, PEGB0
			9'd18 : rdata = 43'b0001101010010011000000000000000000010000000;
			// PEs: 4, 4 -> 0
			// srcs: (20, 19)(133) 10, (7) 46 --> (733) 460:NW19, ND0, *, PEGB0
			9'd19 : rdata = 43'b0001101010011011000000000000000000010000000;
			// PEs: 4, 4 -> 0
			// srcs: (21, 20)(134) 1, (7) 46 --> (734) 46:NW20, ND0, *, PEGB0
			9'd20 : rdata = 43'b0001101010100011000000000000000000010000000;
			// PEs: 4, 4 -> 0
			// srcs: (22, 21)(135) 26, (7) 46 --> (735) 1196:NW21, ND0, *, PEGB0
			9'd21 : rdata = 43'b0001101010101011000000000000000000010000000;
			// PEs: 4, 4 -> 0
			// srcs: (23, 22)(136) 26, (7) 46 --> (736) 1196:NW22, ND0, *, PEGB0
			9'd22 : rdata = 43'b0001101010110011000000000000000000010000000;
			// PEs: 4, 4 -> 0
			// srcs: (24, 23)(137) 18, (7) 46 --> (737) 828:NW23, ND0, *, PEGB0
			9'd23 : rdata = 43'b0001101010111011000000000000000000010000000;
			// PEs: 4, 4 -> 2
			// srcs: (25, 24)(138) 44, (7) 46 --> (738) 2024:NW24, ND0, *, PEGB2
			9'd24 : rdata = 43'b0001101011000011000000000000000000010100000;
			// PEs: 4, 4 -> 2
			// srcs: (26, 25)(139) 0, (7) 46 --> (739) 0:NW25, ND0, *, PEGB2
			9'd25 : rdata = 43'b0001101011001011000000000000000000010100000;
			// PEs: 4, 4 -> 6
			// srcs: (27, 26)(140) 16, (7) 46 --> (740) 736:NW26, ND0, *, PEGB6
			9'd26 : rdata = 43'b0001101011010011000000000000000000011100000;
			// PEs: 4, 4 -> 4
			// srcs: (28, 27)(141) 13, (7) 46 --> (741) 598:NW27, ND0, *, NI0
			9'd27 : rdata = 43'b0001101011011011000001000000000000000000000;
			// PEs: 4, 4 -> 4
			// srcs: (29, 28)(142) 35, (7) 46 --> (742) 1610:NW28, ND0, *, NI1
			9'd28 : rdata = 43'b0001101011100011000001000010000000000000000;
			// PEs: 4, 4 -> 4
			// srcs: (30, 29)(143) 46, (7) 46 --> (743) 2116:NW29, ND0, *, NI2
			9'd29 : rdata = 43'b0001101011101011000001000100000000000000000;
			// PEs: 3, 4 -> 1
			// srcs: (31, 30)(711) 168, (741) 598 --> (1738) 766:PENB, NI0, +, PEGB1
			9'd30 : rdata = 43'b0000111011110101000000000000000000010010000;
			// PEs: 3, 4 -> 1
			// srcs: (32, 31)(712) 888, (742) 1610 --> (1757) 2498:PENB, NI1, +, PEGB1
			9'd31 : rdata = 43'b0000111011110101000010000000000000010010000;
			// PEs: 3, 4 -> 1
			// srcs: (33, 32)(713) 1104, (743) 2116 --> (1776) 3220:PENB, NI2, +, PEGB1
			9'd32 : rdata = 43'b0000111011110101000100000000000000010010000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 5) begin
	always @(*) begin
		case(address)
			// PEs: 5, 5 -> 0
			// srcs: (1, 0)(144) 5, (8) 24 --> (744) 120:NW0, ND0, *, PEGB0
			9'd0 : rdata = 43'b0001101000000011000000000000000000010000000;
			// PEs: 5, 5 -> 0
			// srcs: (2, 1)(145) 42, (8) 24 --> (745) 1008:NW1, ND0, *, PEGB0
			9'd1 : rdata = 43'b0001101000001011000000000000000000010000000;
			// PEs: 5, 5 -> 0
			// srcs: (3, 2)(146) 33, (8) 24 --> (746) 792:NW2, ND0, *, PEGB0
			9'd2 : rdata = 43'b0001101000010011000000000000000000010000000;
			// PEs: 5, 5 -> 0
			// srcs: (4, 3)(147) 36, (8) 24 --> (747) 864:NW3, ND0, *, PEGB0
			9'd3 : rdata = 43'b0001101000011011000000000000000000010000000;
			// PEs: 5, 5 -> 0
			// srcs: (5, 4)(148) 41, (8) 24 --> (748) 984:NW4, ND0, *, PEGB0
			9'd4 : rdata = 43'b0001101000100011000000000000000000010000000;
			// PEs: 5, 5 -> 0
			// srcs: (6, 5)(149) 15, (8) 24 --> (749) 360:NW5, ND0, *, PEGB0
			9'd5 : rdata = 43'b0001101000101011000000000000000000010000000;
			// PEs: 5, 5 -> 0
			// srcs: (7, 6)(150) 34, (8) 24 --> (750) 816:NW6, ND0, *, PEGB0
			9'd6 : rdata = 43'b0001101000110011000000000000000000010000000;
			// PEs: 5, 5 -> 0
			// srcs: (8, 7)(151) 23, (8) 24 --> (751) 552:NW7, ND0, *, PEGB0
			9'd7 : rdata = 43'b0001101000111011000000000000000000010000000;
			// PEs: 5, 5 -> 0
			// srcs: (9, 8)(152) 13, (8) 24 --> (752) 312:NW8, ND0, *, PEGB0
			9'd8 : rdata = 43'b0001101001000011000000000000000000010000000;
			// PEs: 5, 5 -> 0
			// srcs: (10, 9)(153) 34, (8) 24 --> (753) 816:NW9, ND0, *, PEGB0
			9'd9 : rdata = 43'b0001101001001011000000000000000000010000000;
			// PEs: 5, 5 -> 0
			// srcs: (11, 10)(154) 49, (8) 24 --> (754) 1176:NW10, ND0, *, PEGB0
			9'd10 : rdata = 43'b0001101001010011000000000000000000010000000;
			// PEs: 5, 5 -> 0
			// srcs: (12, 11)(155) -1, (8) 24 --> (755) -24:NW11, ND0, *, PEGB0
			9'd11 : rdata = 43'b0001101001011011000000000000000000010000000;
			// PEs: 5, 5 -> 0
			// srcs: (13, 12)(156) 3, (8) 24 --> (756) 72:NW12, ND0, *, PEGB0
			9'd12 : rdata = 43'b0001101001100011000000000000000000010000000;
			// PEs: 5, 5 -> 0
			// srcs: (14, 13)(157) 37, (8) 24 --> (757) 888:NW13, ND0, *, PEGB0
			9'd13 : rdata = 43'b0001101001101011000000000000000000010000000;
			// PEs: 5, 5 -> 0
			// srcs: (15, 14)(158) 39, (8) 24 --> (758) 936:NW14, ND0, *, PEGB0
			9'd14 : rdata = 43'b0001101001110011000000000000000000010000000;
			// PEs: 5, 5 -> 0
			// srcs: (16, 15)(159) 35, (8) 24 --> (759) 840:NW15, ND0, *, PEGB0
			9'd15 : rdata = 43'b0001101001111011000000000000000000010000000;
			// PEs: 5, 5 -> 0
			// srcs: (17, 16)(160) 25, (8) 24 --> (760) 600:NW16, ND0, *, PEGB0
			9'd16 : rdata = 43'b0001101010000011000000000000000000010000000;
			// PEs: 5, 5 -> 0
			// srcs: (18, 17)(161) 28, (8) 24 --> (761) 672:NW17, ND0, *, PEGB0
			9'd17 : rdata = 43'b0001101010001011000000000000000000010000000;
			// PEs: 5, 5 -> 0
			// srcs: (19, 18)(162) 44, (8) 24 --> (762) 1056:NW18, ND0, *, PEGB0
			9'd18 : rdata = 43'b0001101010010011000000000000000000010000000;
			// PEs: 5, 5 -> 0
			// srcs: (20, 19)(163) -3, (8) 24 --> (763) -72:NW19, ND0, *, PEGB0
			9'd19 : rdata = 43'b0001101010011011000000000000000000010000000;
			// PEs: 5, 5 -> 0
			// srcs: (21, 20)(164) 20, (8) 24 --> (764) 480:NW20, ND0, *, PEGB0
			9'd20 : rdata = 43'b0001101010100011000000000000000000010000000;
			// PEs: 5, 5 -> 0
			// srcs: (22, 21)(165) 23, (8) 24 --> (765) 552:NW21, ND0, *, PEGB0
			9'd21 : rdata = 43'b0001101010101011000000000000000000010000000;
			// PEs: 5, 5 -> 0
			// srcs: (23, 22)(166) 21, (8) 24 --> (766) 504:NW22, ND0, *, PEGB0
			9'd22 : rdata = 43'b0001101010110011000000000000000000010000000;
			// PEs: 5, 5 -> 0
			// srcs: (24, 23)(167) 28, (8) 24 --> (767) 672:NW23, ND0, *, PEGB0
			9'd23 : rdata = 43'b0001101010111011000000000000000000010000000;
			// PEs: 5, 5 -> 3
			// srcs: (25, 24)(168) 46, (8) 24 --> (768) 1104:NW24, ND0, *, PEGB3
			9'd24 : rdata = 43'b0001101011000011000000000000000000010110000;
			// PEs: 5, 5 -> 3
			// srcs: (26, 25)(169) 16, (8) 24 --> (769) 384:NW25, ND0, *, PEGB3
			9'd25 : rdata = 43'b0001101011001011000000000000000000010110000;
			// PEs: 5, 5 -> 7
			// srcs: (27, 26)(170) 20, (8) 24 --> (770) 480:NW26, ND0, *, PEGB7
			9'd26 : rdata = 43'b0001101011010011000000000000000000011110000;
			// PEs: 5, 5 -> 6
			// srcs: (28, 27)(171) 32, (8) 24 --> (771) 768:NW27, ND0, *, PENB
			9'd27 : rdata = 43'b0001101011011011000000000000000000100000000;
			// PEs: 5, 5 -> 2
			// srcs: (29, 28)(172) 37, (8) 24 --> (772) 888:NW28, ND0, *, PEGB2
			9'd28 : rdata = 43'b0001101011100011000000000000000000010100000;
			// PEs: 5, 5 -> 6
			// srcs: (30, 29)(173) 34, (8) 24 --> (773) 816:NW29, ND0, *, PENB
			9'd29 : rdata = 43'b0001101011101011000000000000000000100000000;
			// PEs: 2 -> 
			// srcs: (32, 30)(680) 473 --> (680) 473:PEGB2, pass, 
			9'd30 : rdata = 43'b1100011100100000000000000000000000000000000;
			// PEs: 1, 5 -> 6
			// srcs: (35, 31)(650) 378, (680) 473 --> (1718) 851:PEGB1, ALU, +, PENB
			9'd31 : rdata = 43'b0000111100010001111110000000000000100000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 6) begin
	always @(*) begin
		case(address)
			// PEs: 6, 6 -> 0
			// srcs: (1, 0)(174) 38, (9) 19 --> (774) 722:NW0, ND0, *, PEGB0
			9'd0 : rdata = 43'b0001101000000011000000000000000000010000000;
			// PEs: 6, 6 -> 0
			// srcs: (2, 1)(175) 29, (9) 19 --> (775) 551:NW1, ND0, *, PEGB0
			9'd1 : rdata = 43'b0001101000001011000000000000000000010000000;
			// PEs: 6, 6 -> 0
			// srcs: (3, 2)(176) 19, (9) 19 --> (776) 361:NW2, ND0, *, PEGB0
			9'd2 : rdata = 43'b0001101000010011000000000000000000010000000;
			// PEs: 6, 6 -> 0
			// srcs: (4, 3)(177) 37, (9) 19 --> (777) 703:NW3, ND0, *, PEGB0
			9'd3 : rdata = 43'b0001101000011011000000000000000000010000000;
			// PEs: 6, 6 -> 0
			// srcs: (5, 4)(178) 28, (9) 19 --> (778) 532:NW4, ND0, *, PEGB0
			9'd4 : rdata = 43'b0001101000100011000000000000000000010000000;
			// PEs: 6, 6 -> 0
			// srcs: (6, 5)(179) 5, (9) 19 --> (779) 95:NW5, ND0, *, PEGB0
			9'd5 : rdata = 43'b0001101000101011000000000000000000010000000;
			// PEs: 6, 6 -> 0
			// srcs: (7, 6)(180) 45, (9) 19 --> (780) 855:NW6, ND0, *, PEGB0
			9'd6 : rdata = 43'b0001101000110011000000000000000000010000000;
			// PEs: 6, 6 -> 0
			// srcs: (8, 7)(181) 6, (9) 19 --> (781) 114:NW7, ND0, *, PEGB0
			9'd7 : rdata = 43'b0001101000111011000000000000000000010000000;
			// PEs: 6, 6 -> 0
			// srcs: (9, 8)(182) 31, (9) 19 --> (782) 589:NW8, ND0, *, PEGB0
			9'd8 : rdata = 43'b0001101001000011000000000000000000010000000;
			// PEs: 6, 6 -> 0
			// srcs: (10, 9)(183) 44, (9) 19 --> (783) 836:NW9, ND0, *, PEGB0
			9'd9 : rdata = 43'b0001101001001011000000000000000000010000000;
			// PEs: 6, 6 -> 0
			// srcs: (11, 10)(184) -2, (9) 19 --> (784) -38:NW10, ND0, *, PEGB0
			9'd10 : rdata = 43'b0001101001010011000000000000000000010000000;
			// PEs: 6, 6 -> 0
			// srcs: (12, 11)(185) 16, (9) 19 --> (785) 304:NW11, ND0, *, PEGB0
			9'd11 : rdata = 43'b0001101001011011000000000000000000010000000;
			// PEs: 6, 6 -> 0
			// srcs: (13, 12)(186) 14, (9) 19 --> (786) 266:NW12, ND0, *, PEGB0
			9'd12 : rdata = 43'b0001101001100011000000000000000000010000000;
			// PEs: 6, 6 -> 0
			// srcs: (14, 13)(187) 39, (9) 19 --> (787) 741:NW13, ND0, *, PEGB0
			9'd13 : rdata = 43'b0001101001101011000000000000000000010000000;
			// PEs: 6, 6 -> 0
			// srcs: (15, 14)(188) 21, (9) 19 --> (788) 399:NW14, ND0, *, PEGB0
			9'd14 : rdata = 43'b0001101001110011000000000000000000010000000;
			// PEs: 6, 6 -> 0
			// srcs: (16, 15)(189) 28, (9) 19 --> (789) 532:NW15, ND0, *, PEGB0
			9'd15 : rdata = 43'b0001101001111011000000000000000000010000000;
			// PEs: 6, 6 -> 0
			// srcs: (17, 16)(190) 41, (9) 19 --> (790) 779:NW16, ND0, *, PEGB0
			9'd16 : rdata = 43'b0001101010000011000000000000000000010000000;
			// PEs: 6, 6 -> 0
			// srcs: (18, 17)(191) 38, (9) 19 --> (791) 722:NW17, ND0, *, PEGB0
			9'd17 : rdata = 43'b0001101010001011000000000000000000010000000;
			// PEs: 6, 6 -> 0
			// srcs: (19, 18)(192) 6, (9) 19 --> (792) 114:NW18, ND0, *, PEGB0
			9'd18 : rdata = 43'b0001101010010011000000000000000000010000000;
			// PEs: 6, 6 -> 0
			// srcs: (20, 19)(193) 5, (9) 19 --> (793) 95:NW19, ND0, *, PEGB0
			9'd19 : rdata = 43'b0001101010011011000000000000000000010000000;
			// PEs: 6, 6 -> 0
			// srcs: (21, 20)(194) 42, (9) 19 --> (794) 798:NW20, ND0, *, PEGB0
			9'd20 : rdata = 43'b0001101010100011000000000000000000010000000;
			// PEs: 6, 6 -> 0
			// srcs: (22, 21)(195) 11, (9) 19 --> (795) 209:NW21, ND0, *, PEGB0
			9'd21 : rdata = 43'b0001101010101011000000000000000000010000000;
			// PEs: 6, 6 -> 0
			// srcs: (23, 22)(196) 24, (9) 19 --> (796) 456:NW22, ND0, *, PEGB0
			9'd22 : rdata = 43'b0001101010110011000000000000000000010000000;
			// PEs: 6, 6 -> 0
			// srcs: (24, 23)(197) 21, (9) 19 --> (797) 399:NW23, ND0, *, PEGB0
			9'd23 : rdata = 43'b0001101010111011000000000000000000010000000;
			// PEs: 6, 6 -> 3
			// srcs: (25, 24)(198) 28, (9) 19 --> (798) 532:NW24, ND0, *, PEGB3
			9'd24 : rdata = 43'b0001101011000011000000000000000000010110000;
			// PEs: 6, 6 -> 3
			// srcs: (26, 25)(199) 35, (9) 19 --> (799) 665:NW25, ND0, *, PEGB3
			9'd25 : rdata = 43'b0001101011001011000000000000000000010110000;
			// PEs: 6, 6 -> 7
			// srcs: (27, 26)(200) 7, (9) 19 --> (800) 133:NW26, ND0, *, PENB
			9'd26 : rdata = 43'b0001101011010011000000000000000000100000000;
			// PEs: 6, 6 -> 6
			// srcs: (28, 27)(201) 5, (9) 19 --> (801) 95:NW27, ND0, *, NI0
			9'd27 : rdata = 43'b0001101011011011000001000000000000000000000;
			// PEs: 6, 6 -> 2
			// srcs: (29, 28)(202) 34, (9) 19 --> (802) 646:NW28, ND0, *, PEGB2
			9'd28 : rdata = 43'b0001101011100011000000000000000000010100000;
			// PEs: 6, 6 -> 6
			// srcs: (30, 29)(203) 34, (9) 19 --> (803) 646:NW29, ND0, *, NI1
			9'd29 : rdata = 43'b0001101011101011000001000010000000000000000;
			// PEs: 5, 6 -> 0
			// srcs: (31, 32)(771) 768, (801) 95 --> (1739) 863:PENB, NI0, +, PEGB0
			9'd30 : rdata = 43'b0000111011110101000000000000000000010000000;
			// PEs: 4 -> 6
			// srcs: (32, 30)(740) 736 --> (740) 736:PEGB4, pass, NI0
			9'd31 : rdata = 43'b1100011101000000000001000000000000000000000;
			// PEs: 5, 6 -> 0
			// srcs: (33, 33)(773) 816, (803) 646 --> (1777) 1462:PENB, NI1, +, PEGB0
			9'd32 : rdata = 43'b0000111011110101000010000000000000010000000;
			// PEs: 3, 6 -> 
			// srcs: (35, 31)(710) 1128, (740) 736 --> (1719) 1864:PEGB3, NI0, +, 
			9'd33 : rdata = 43'b0000111100110101000000000000000000000000000;
			// PEs: 5, 6 -> 0
			// srcs: (38, 34)(1718) 851, (1719) 1864 --> (1728) 2715:PENB, ALU, +, PEGB0
			9'd34 : rdata = 43'b0000111011110001111110000000000000010000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 7) begin
	always @(*) begin
		case(address)
			// PEs: 7, 7 -> 0
			// srcs: (1, 0)(204) 45, (10) 31 --> (804) 1395:NW0, ND0, *, PENB
			9'd0 : rdata = 43'b0001101000000011000000000000000000100000000;
			// PEs: 7, 7 -> 0
			// srcs: (2, 1)(205) 30, (10) 31 --> (805) 930:NW1, ND0, *, PENB
			9'd1 : rdata = 43'b0001101000001011000000000000000000100000000;
			// PEs: 7, 7 -> 0
			// srcs: (3, 2)(206) 12, (10) 31 --> (806) 372:NW2, ND0, *, PENB
			9'd2 : rdata = 43'b0001101000010011000000000000000000100000000;
			// PEs: 7, 7 -> 0
			// srcs: (4, 3)(207) 10, (10) 31 --> (807) 310:NW3, ND0, *, PENB
			9'd3 : rdata = 43'b0001101000011011000000000000000000100000000;
			// PEs: 7, 7 -> 0
			// srcs: (5, 4)(208) -3, (10) 31 --> (808) -93:NW4, ND0, *, PENB
			9'd4 : rdata = 43'b0001101000100011000000000000000000100000000;
			// PEs: 7, 7 -> 0
			// srcs: (6, 5)(209) 10, (10) 31 --> (809) 310:NW5, ND0, *, PENB
			9'd5 : rdata = 43'b0001101000101011000000000000000000100000000;
			// PEs: 7, 7 -> 0
			// srcs: (7, 6)(210) 38, (10) 31 --> (810) 1178:NW6, ND0, *, PENB
			9'd6 : rdata = 43'b0001101000110011000000000000000000100000000;
			// PEs: 7, 7 -> 0
			// srcs: (8, 7)(211) 9, (10) 31 --> (811) 279:NW7, ND0, *, PENB
			9'd7 : rdata = 43'b0001101000111011000000000000000000100000000;
			// PEs: 7, 7 -> 0
			// srcs: (9, 8)(212) 47, (10) 31 --> (812) 1457:NW8, ND0, *, PENB
			9'd8 : rdata = 43'b0001101001000011000000000000000000100000000;
			// PEs: 7, 7 -> 0
			// srcs: (10, 9)(213) 2, (10) 31 --> (813) 62:NW9, ND0, *, PENB
			9'd9 : rdata = 43'b0001101001001011000000000000000000100000000;
			// PEs: 7, 7 -> 0
			// srcs: (11, 10)(214) 24, (10) 31 --> (814) 744:NW10, ND0, *, PENB
			9'd10 : rdata = 43'b0001101001010011000000000000000000100000000;
			// PEs: 7, 7 -> 0
			// srcs: (12, 11)(215) 34, (10) 31 --> (815) 1054:NW11, ND0, *, PENB
			9'd11 : rdata = 43'b0001101001011011000000000000000000100000000;
			// PEs: 7, 7 -> 0
			// srcs: (13, 12)(216) 11, (10) 31 --> (816) 341:NW12, ND0, *, PENB
			9'd12 : rdata = 43'b0001101001100011000000000000000000100000000;
			// PEs: 7, 7 -> 0
			// srcs: (14, 13)(217) 12, (10) 31 --> (817) 372:NW13, ND0, *, PENB
			9'd13 : rdata = 43'b0001101001101011000000000000000000100000000;
			// PEs: 7, 7 -> 0
			// srcs: (15, 14)(218) 27, (10) 31 --> (818) 837:NW14, ND0, *, PENB
			9'd14 : rdata = 43'b0001101001110011000000000000000000100000000;
			// PEs: 7, 7 -> 0
			// srcs: (16, 15)(219) 28, (10) 31 --> (819) 868:NW15, ND0, *, PENB
			9'd15 : rdata = 43'b0001101001111011000000000000000000100000000;
			// PEs: 7, 7 -> 0
			// srcs: (17, 16)(220) 27, (10) 31 --> (820) 837:NW16, ND0, *, PENB
			9'd16 : rdata = 43'b0001101010000011000000000000000000100000000;
			// PEs: 7, 7 -> 0
			// srcs: (18, 17)(221) 27, (10) 31 --> (821) 837:NW17, ND0, *, PENB
			9'd17 : rdata = 43'b0001101010001011000000000000000000100000000;
			// PEs: 7, 7 -> 0
			// srcs: (19, 18)(222) 44, (10) 31 --> (822) 1364:NW18, ND0, *, PENB
			9'd18 : rdata = 43'b0001101010010011000000000000000000100000000;
			// PEs: 7, 7 -> 0
			// srcs: (20, 19)(223) 20, (10) 31 --> (823) 620:NW19, ND0, *, PENB
			9'd19 : rdata = 43'b0001101010011011000000000000000000100000000;
			// PEs: 7, 7 -> 0
			// srcs: (21, 20)(224) 23, (10) 31 --> (824) 713:NW20, ND0, *, PENB
			9'd20 : rdata = 43'b0001101010100011000000000000000000100000000;
			// PEs: 7, 7 -> 0
			// srcs: (22, 21)(225) 13, (10) 31 --> (825) 403:NW21, ND0, *, PENB
			9'd21 : rdata = 43'b0001101010101011000000000000000000100000000;
			// PEs: 7, 7 -> 0
			// srcs: (23, 22)(226) 8, (10) 31 --> (826) 248:NW22, ND0, *, PENB
			9'd22 : rdata = 43'b0001101010110011000000000000000000100000000;
			// PEs: 7, 7 -> 0
			// srcs: (24, 23)(227) 7, (10) 31 --> (827) 217:NW23, ND0, *, PENB
			9'd23 : rdata = 43'b0001101010111011000000000000000000100000000;
			// PEs: 7, 7 -> 0
			// srcs: (25, 24)(228) 41, (10) 31 --> (828) 1271:NW24, ND0, *, PENB
			9'd24 : rdata = 43'b0001101011000011000000000000000000100000000;
			// PEs: 7, 7 -> 0
			// srcs: (26, 25)(229) 32, (10) 31 --> (829) 992:NW25, ND0, *, PENB
			9'd25 : rdata = 43'b0001101011001011000000000000000000100000000;
			// PEs: 7, 7 -> 0
			// srcs: (27, 26)(230) 26, (10) 31 --> (830) 806:NW26, ND0, *, PENB
			9'd26 : rdata = 43'b0001101011010011000000000000000000100000000;
			// PEs: 7, 7 -> 0
			// srcs: (28, 27)(231) 24, (10) 31 --> (831) 744:NW27, ND0, *, PENB
			9'd27 : rdata = 43'b0001101011011011000000000000000000100000000;
			// PEs: 7, 7 -> 0
			// srcs: (29, 28)(232) 11, (10) 31 --> (832) 341:NW28, ND0, *, PENB
			9'd28 : rdata = 43'b0001101011100011000000000000000000100000000;
			// PEs: 7, 7 -> 0
			// srcs: (30, 29)(233) 15, (10) 31 --> (833) 465:NW29, ND0, *, PENB
			9'd29 : rdata = 43'b0001101011101011000000000000000000100000000;
			// PEs: 5, 6 -> 0
			// srcs: (33, 30)(770) 480, (800) 133 --> (1720) 613:PEGB5, PENB, +, PENB
			9'd30 : rdata = 43'b0000111101010110111100000000000000100000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 8) begin
	always @(*) begin
		case(address)
			// PEs: 9 -> 16
			// srcs: (6, 0)(834) 992 --> (834) 992:PEGB1, pass, PUNB
			9'd0 : rdata = 43'b1100011100010000000000000000000001000000000;
			// PEs: 10 -> 32
			// srcs: (7, 1)(864) 1216 --> (864) 1216:PEGB2, pass, PUGB4
			9'd1 : rdata = 43'b1100011100100000000000000000000000000001100;
			// PEs: 11 -> 32
			// srcs: (8, 2)(894) -22 --> (894) -22:PEGB3, pass, PUGB4
			9'd2 : rdata = 43'b1100011100110000000000000000000000000001100;
			// PEs: 12 -> 32
			// srcs: (9, 3)(924) 667 --> (924) 667:PEGB4, pass, PUGB4
			9'd3 : rdata = 43'b1100011101000000000000000000000000000001100;
			// PEs: 13 -> 32
			// srcs: (10, 4)(954) 1551 --> (954) 1551:PEGB5, pass, PUGB4
			9'd4 : rdata = 43'b1100011101010000000000000000000000000001100;
			// PEs: 14 -> 32
			// srcs: (11, 5)(984) 92 --> (984) 92:PEGB6, pass, PUGB4
			9'd5 : rdata = 43'b1100011101100000000000000000000000000001100;
			// PEs: 15 -> 32
			// srcs: (12, 6)(1014) 462 --> (1014) 462:PENB, pass, PUGB4
			9'd6 : rdata = 43'b1100011011110000000000000000000000000001100;
			// PEs: 9 -> 16
			// srcs: (13, 7)(835) 32 --> (835) 32:PEGB1, pass, PUNB
			9'd7 : rdata = 43'b1100011100010000000000000000000001000000000;
			// PEs: 10 -> 16
			// srcs: (14, 8)(865) 1312 --> (865) 1312:PEGB2, pass, PUNB
			9'd8 : rdata = 43'b1100011100100000000000000000000001000000000;
			// PEs: 11 -> 16
			// srcs: (15, 9)(895) -23 --> (895) -23:PEGB3, pass, PUNB
			9'd9 : rdata = 43'b1100011100110000000000000000000001000000000;
			// PEs: 12 -> 16
			// srcs: (16, 10)(925) 638 --> (925) 638:PEGB4, pass, PUNB
			9'd10 : rdata = 43'b1100011101000000000000000000000001000000000;
			// PEs: 13 -> 16
			// srcs: (17, 11)(955) 462 --> (955) 462:PEGB5, pass, PUNB
			9'd11 : rdata = 43'b1100011101010000000000000000000001000000000;
			// PEs: 14 -> 16
			// srcs: (18, 12)(985) 52 --> (985) 52:PEGB6, pass, PUNB
			9'd12 : rdata = 43'b1100011101100000000000000000000001000000000;
			// PEs: 15 -> 16
			// srcs: (19, 13)(1015) 44 --> (1015) 44:PENB, pass, PUNB
			9'd13 : rdata = 43'b1100011011110000000000000000000001000000000;
			// PEs: 9 -> 24
			// srcs: (20, 14)(836) 672 --> (836) 672:PEGB1, pass, PUGB3
			9'd14 : rdata = 43'b1100011100010000000000000000000000000001011;
			// PEs: 10 -> 24
			// srcs: (21, 15)(866) 416 --> (866) 416:PEGB2, pass, PUGB3
			9'd15 : rdata = 43'b1100011100100000000000000000000000000001011;
			// PEs: 11 -> 24
			// srcs: (22, 16)(896) -5 --> (896) -5:PEGB3, pass, PUGB3
			9'd16 : rdata = 43'b1100011100110000000000000000000000000001011;
			// PEs: 12 -> 40
			// srcs: (23, 17)(926) 116 --> (926) 116:PEGB4, pass, PUGB5
			9'd17 : rdata = 43'b1100011101000000000000000000000000000001101;
			// PEs: 13 -> 40
			// srcs: (24, 18)(956) 165 --> (956) 165:PEGB5, pass, PUGB5
			9'd18 : rdata = 43'b1100011101010000000000000000000000000001101;
			// PEs: 14 -> 40
			// srcs: (25, 19)(986) 56 --> (986) 56:PEGB6, pass, PUGB5
			9'd19 : rdata = 43'b1100011101100000000000000000000000000001101;
			// PEs: 15 -> 40
			// srcs: (26, 20)(1016) -22 --> (1016) -22:PENB, pass, PUGB5
			9'd20 : rdata = 43'b1100011011110000000000000000000000000001101;
			// PEs: 9 -> 40
			// srcs: (27, 21)(837) 1440 --> (837) 1440:PEGB1, pass, PUGB5
			9'd21 : rdata = 43'b1100011100010000000000000000000000000001101;
			// PEs: 10 -> 40
			// srcs: (28, 22)(867) 896 --> (867) 896:PEGB2, pass, PUGB5
			9'd22 : rdata = 43'b1100011100100000000000000000000000000001101;
			// PEs: 11 -> 40
			// srcs: (29, 23)(897) -9 --> (897) -9:PEGB3, pass, PUGB5
			9'd23 : rdata = 43'b1100011100110000000000000000000000000001101;
			// PEs: 12 -> 40
			// srcs: (30, 24)(927) 29 --> (927) 29:PEGB4, pass, PUGB5
			9'd24 : rdata = 43'b1100011101000000000000000000000000000001101;
			// PEs: 13 -> 40
			// srcs: (31, 25)(957) 1320 --> (957) 1320:PEGB5, pass, PUGB5
			9'd25 : rdata = 43'b1100011101010000000000000000000000000001101;
			// PEs: 14 -> 40
			// srcs: (32, 26)(987) 94 --> (987) 94:PEGB6, pass, PUGB5
			9'd26 : rdata = 43'b1100011101100000000000000000000000000001101;
			// PEs: 15 -> 40
			// srcs: (33, 27)(1017) 968 --> (1017) 968:PENB, pass, PUGB5
			9'd27 : rdata = 43'b1100011011110000000000000000000000000001101;
			// PEs: 9 -> 48
			// srcs: (34, 28)(838) 256 --> (838) 256:PEGB1, pass, PUGB6
			9'd28 : rdata = 43'b1100011100010000000000000000000000000001110;
			// PEs: 10 -> 48
			// srcs: (35, 29)(868) 32 --> (868) 32:PEGB2, pass, PUGB6
			9'd29 : rdata = 43'b1100011100100000000000000000000000000001110;
			// PEs: 11 -> 48
			// srcs: (36, 30)(898) -9 --> (898) -9:PEGB3, pass, PUGB6
			9'd30 : rdata = 43'b1100011100110000000000000000000000000001110;
			// PEs: 12 -> 48
			// srcs: (37, 31)(928) 29 --> (928) 29:PEGB4, pass, PUGB6
			9'd31 : rdata = 43'b1100011101000000000000000000000000000001110;
			// PEs: 13 -> 48
			// srcs: (38, 32)(958) 759 --> (958) 759:PEGB5, pass, PUGB6
			9'd32 : rdata = 43'b1100011101010000000000000000000000000001110;
			// PEs: 14 -> 48
			// srcs: (39, 33)(988) 18 --> (988) 18:PEGB6, pass, PUGB6
			9'd33 : rdata = 43'b1100011101100000000000000000000000000001110;
			// PEs: 15 -> 48
			// srcs: (40, 34)(1018) 440 --> (1018) 440:PENB, pass, PUGB6
			9'd34 : rdata = 43'b1100011011110000000000000000000000000001110;
			// PEs: 9 -> 56
			// srcs: (41, 35)(839) 736 --> (839) 736:PEGB1, pass, PUGB7
			9'd35 : rdata = 43'b1100011100010000000000000000000000000001111;
			// PEs: 10 -> 56
			// srcs: (42, 36)(869) 704 --> (869) 704:PEGB2, pass, PUGB7
			9'd36 : rdata = 43'b1100011100100000000000000000000000000001111;
			// PEs: 11 -> 56
			// srcs: (43, 37)(899) -4 --> (899) -4:PEGB3, pass, PUGB7
			9'd37 : rdata = 43'b1100011100110000000000000000000000000001111;
			// PEs: 12 -> 56
			// srcs: (44, 38)(929) 1015 --> (929) 1015:PEGB4, pass, PUGB7
			9'd38 : rdata = 43'b1100011101000000000000000000000000000001111;
			// PEs: 13 -> 56
			// srcs: (45, 39)(959) 990 --> (959) 990:PEGB5, pass, PUGB7
			9'd39 : rdata = 43'b1100011101010000000000000000000000000001111;
			// PEs: 14 -> 56
			// srcs: (46, 40)(989) 90 --> (989) 90:PEGB6, pass, PUGB7
			9'd40 : rdata = 43'b1100011101100000000000000000000000000001111;
			// PEs: 15 -> 56
			// srcs: (47, 41)(1019) 506 --> (1019) 506:PENB, pass, PUGB7
			9'd41 : rdata = 43'b1100011011110000000000000000000000000001111;
			// PEs: 9 -> 32
			// srcs: (48, 42)(840) 64 --> (840) 64:PEGB1, pass, PUGB4
			9'd42 : rdata = 43'b1100011100010000000000000000000000000001100;
			// PEs: 10 -> 32
			// srcs: (49, 43)(870) 1024 --> (870) 1024:PEGB2, pass, PUGB4
			9'd43 : rdata = 43'b1100011100100000000000000000000000000001100;
			// PEs: 11 -> 32
			// srcs: (50, 44)(900) 2 --> (900) 2:PEGB3, pass, PUGB4
			9'd44 : rdata = 43'b1100011100110000000000000000000000000001100;
			// PEs: 12 -> 32
			// srcs: (51, 45)(930) 1305 --> (930) 1305:PEGB4, pass, PUGB4
			9'd45 : rdata = 43'b1100011101000000000000000000000000000001100;
			// PEs: 13 -> 32
			// srcs: (52, 46)(960) -33 --> (960) -33:PEGB5, pass, PUGB4
			9'd46 : rdata = 43'b1100011101010000000000000000000000000001100;
			// PEs: 14 -> 32
			// srcs: (53, 47)(990) 82 --> (990) 82:PEGB6, pass, PUGB4
			9'd47 : rdata = 43'b1100011101100000000000000000000000000001100;
			// PEs: 15 -> 32
			// srcs: (54, 48)(1020) -22 --> (1020) -22:PENB, pass, PUGB4
			9'd48 : rdata = 43'b1100011011110000000000000000000000000001100;
			// PEs: 9 -> 16
			// srcs: (55, 49)(841) -96 --> (841) -96:PEGB1, pass, PUNB
			9'd49 : rdata = 43'b1100011100010000000000000000000001000000000;
			// PEs: 10 -> 16
			// srcs: (56, 50)(871) 928 --> (871) 928:PEGB2, pass, PUNB
			9'd50 : rdata = 43'b1100011100100000000000000000000001000000000;
			// PEs: 11 -> 16
			// srcs: (57, 51)(901) -47 --> (901) -47:PEGB3, pass, PUNB
			9'd51 : rdata = 43'b1100011100110000000000000000000001000000000;
			// PEs: 12 -> 16
			// srcs: (58, 52)(931) 464 --> (931) 464:PEGB4, pass, PUNB
			9'd52 : rdata = 43'b1100011101000000000000000000000001000000000;
			// PEs: 13 -> 16
			// srcs: (59, 53)(961) 363 --> (961) 363:PEGB5, pass, PUNB
			9'd53 : rdata = 43'b1100011101010000000000000000000001000000000;
			// PEs: 14 -> 16
			// srcs: (60, 54)(991) 50 --> (991) 50:PEGB6, pass, PUNB
			9'd54 : rdata = 43'b1100011101100000000000000000000001000000000;
			// PEs: 15 -> 16
			// srcs: (61, 55)(1021) 880 --> (1021) 880:PENB, pass, PUNB
			9'd55 : rdata = 43'b1100011011110000000000000000000001000000000;
			// PEs: 9 -> 16
			// srcs: (62, 56)(842) 416 --> (842) 416:PEGB1, pass, PUNB
			9'd56 : rdata = 43'b1100011100010000000000000000000001000000000;
			// PEs: 10 -> 16
			// srcs: (63, 57)(872) 1024 --> (872) 1024:PEGB2, pass, PUNB
			9'd57 : rdata = 43'b1100011100100000000000000000000001000000000;
			// PEs: 11 -> 16
			// srcs: (64, 58)(902) -45 --> (902) -45:PEGB3, pass, PUNB
			9'd58 : rdata = 43'b1100011100110000000000000000000001000000000;
			// PEs: 12 -> 16
			// srcs: (65, 59)(932) 580 --> (932) 580:PEGB4, pass, PUNB
			9'd59 : rdata = 43'b1100011101000000000000000000000001000000000;
			// PEs: 13 -> 16
			// srcs: (66, 60)(962) 99 --> (962) 99:PEGB5, pass, PUNB
			9'd60 : rdata = 43'b1100011101010000000000000000000001000000000;
			// PEs: 14 -> 16
			// srcs: (67, 61)(992) 50 --> (992) 50:PEGB6, pass, PUNB
			9'd61 : rdata = 43'b1100011101100000000000000000000001000000000;
			// PEs: 15 -> 16
			// srcs: (68, 62)(1022) 66 --> (1022) 66:PENB, pass, PUNB
			9'd62 : rdata = 43'b1100011011110000000000000000000001000000000;
			// PEs: 9 -> 32
			// srcs: (69, 63)(843) 1344 --> (843) 1344:PEGB1, pass, PUGB4
			9'd63 : rdata = 43'b1100011100010000000000000000000000000001100;
			// PEs: 10 -> 32
			// srcs: (70, 64)(873) 352 --> (873) 352:PEGB2, pass, PUGB4
			9'd64 : rdata = 43'b1100011100100000000000000000000000000001100;
			// PEs: 11 -> 32
			// srcs: (71, 65)(903) -37 --> (903) -37:PEGB3, pass, PUGB4
			9'd65 : rdata = 43'b1100011100110000000000000000000000000001100;
			// PEs: 12 -> 32
			// srcs: (72, 66)(933) 406 --> (933) 406:PEGB4, pass, PUGB4
			9'd66 : rdata = 43'b1100011101000000000000000000000000000001100;
			// PEs: 13 -> 32
			// srcs: (73, 67)(963) 33 --> (963) 33:PEGB5, pass, PUGB4
			9'd67 : rdata = 43'b1100011101010000000000000000000000000001100;
			// PEs: 14 -> 32
			// srcs: (74, 68)(993) 74 --> (993) 74:PEGB6, pass, PUGB4
			9'd68 : rdata = 43'b1100011101100000000000000000000000000001100;
			// PEs: 15 -> 32
			// srcs: (75, 69)(1023) 616 --> (1023) 616:PENB, pass, PUGB4
			9'd69 : rdata = 43'b1100011011110000000000000000000000000001100;
			// PEs: 9 -> 40
			// srcs: (76, 70)(844) 160 --> (844) 160:PEGB1, pass, PUGB5
			9'd70 : rdata = 43'b1100011100010000000000000000000000000001101;
			// PEs: 10 -> 40
			// srcs: (77, 71)(874) 1568 --> (874) 1568:PEGB2, pass, PUGB5
			9'd71 : rdata = 43'b1100011100100000000000000000000000000001101;
			// PEs: 11 -> 40
			// srcs: (78, 72)(904) -4 --> (904) -4:PEGB3, pass, PUGB5
			9'd72 : rdata = 43'b1100011100110000000000000000000000000001101;
			// PEs: 12 -> 48
			// srcs: (79, 73)(934) 1131 --> (934) 1131:PEGB4, pass, PUGB6
			9'd73 : rdata = 43'b1100011101000000000000000000000000000001110;
			// PEs: 13 -> 48
			// srcs: (80, 74)(964) 726 --> (964) 726:PEGB5, pass, PUGB6
			9'd74 : rdata = 43'b1100011101010000000000000000000000000001110;
			// PEs: 14 -> 48
			// srcs: (81, 75)(994) 22 --> (994) 22:PEGB6, pass, PUGB6
			9'd75 : rdata = 43'b1100011101100000000000000000000000000001110;
			// PEs: 15 -> 48
			// srcs: (82, 76)(1024) 836 --> (1024) 836:PENB, pass, PUGB6
			9'd76 : rdata = 43'b1100011011110000000000000000000000000001110;
			// PEs: 9 -> 56
			// srcs: (83, 77)(845) 672 --> (845) 672:PEGB1, pass, PUGB7
			9'd77 : rdata = 43'b1100011100010000000000000000000000000001111;
			// PEs: 10 -> 56
			// srcs: (84, 78)(875) 1536 --> (875) 1536:PEGB2, pass, PUGB7
			9'd78 : rdata = 43'b1100011100100000000000000000000000000001111;
			// PEs: 11 -> 56
			// srcs: (85, 79)(905) -35 --> (905) -35:PEGB3, pass, PUGB7
			9'd79 : rdata = 43'b1100011100110000000000000000000000000001111;
			// PEs: 12 -> 56
			// srcs: (86, 80)(935) 1044 --> (935) 1044:PEGB4, pass, PUGB7
			9'd80 : rdata = 43'b1100011101000000000000000000000000000001111;
			// PEs: 13 -> 56
			// srcs: (87, 81)(965) -99 --> (965) -99:PEGB5, pass, PUGB7
			9'd81 : rdata = 43'b1100011101010000000000000000000000000001111;
			// PEs: 14 -> 56
			// srcs: (88, 82)(995) 60 --> (995) 60:PEGB6, pass, PUGB7
			9'd82 : rdata = 43'b1100011101100000000000000000000000000001111;
			// PEs: 15 -> 56
			// srcs: (89, 83)(1025) 308 --> (1025) 308:PENB, pass, PUGB7
			9'd83 : rdata = 43'b1100011011110000000000000000000000000001111;
			// PEs: 9 -> 16
			// srcs: (90, 84)(846) 448 --> (846) 448:PEGB1, pass, PUNB
			9'd84 : rdata = 43'b1100011100010000000000000000000001000000000;
			// PEs: 10 -> 16
			// srcs: (91, 85)(876) 704 --> (876) 704:PEGB2, pass, PUNB
			9'd85 : rdata = 43'b1100011100100000000000000000000001000000000;
			// PEs: 11 -> 16
			// srcs: (92, 86)(906) -28 --> (906) -28:PEGB3, pass, PUNB
			9'd86 : rdata = 43'b1100011100110000000000000000000001000000000;
			// PEs: 12 -> 16
			// srcs: (93, 87)(936) 290 --> (936) 290:PEGB4, pass, PUNB
			9'd87 : rdata = 43'b1100011101000000000000000000000001000000000;
			// PEs: 13 -> 16
			// srcs: (94, 88)(966) 1518 --> (966) 1518:PEGB5, pass, PUNB
			9'd88 : rdata = 43'b1100011101010000000000000000000001000000000;
			// PEs: 14 -> 16
			// srcs: (95, 89)(996) 64 --> (996) 64:PEGB6, pass, PUNB
			9'd89 : rdata = 43'b1100011101100000000000000000000001000000000;
			// PEs: 15 -> 16
			// srcs: (96, 90)(1026) -22 --> (1026) -22:PENB, pass, PUNB
			9'd90 : rdata = 43'b1100011011110000000000000000000001000000000;
			// PEs: 9 -> 16
			// srcs: (97, 91)(847) 1568 --> (847) 1568:PEGB1, pass, PUNB
			9'd91 : rdata = 43'b1100011100010000000000000000000001000000000;
			// PEs: 10 -> 16
			// srcs: (98, 92)(877) 1024 --> (877) 1024:PEGB2, pass, PUNB
			9'd92 : rdata = 43'b1100011100100000000000000000000001000000000;
			// PEs: 11 -> 16
			// srcs: (99, 93)(907) -13 --> (907) -13:PEGB3, pass, PUNB
			9'd93 : rdata = 43'b1100011100110000000000000000000001000000000;
			// PEs: 12 -> 16
			// srcs: (100, 94)(937) 551 --> (937) 551:PEGB4, pass, PUNB
			9'd94 : rdata = 43'b1100011101000000000000000000000001000000000;
			// PEs: 13 -> 16
			// srcs: (101, 95)(967) 1485 --> (967) 1485:PEGB5, pass, PUNB
			9'd95 : rdata = 43'b1100011101010000000000000000000001000000000;
			// PEs: 14 -> 16
			// srcs: (102, 96)(997) 78 --> (997) 78:PEGB6, pass, PUNB
			9'd96 : rdata = 43'b1100011101100000000000000000000001000000000;
			// PEs: 15 -> 16
			// srcs: (103, 97)(1027) 792 --> (1027) 792:PENB, pass, PUNB
			9'd97 : rdata = 43'b1100011011110000000000000000000001000000000;
			// PEs: 9 -> 32
			// srcs: (104, 98)(848) 864 --> (848) 864:PEGB1, pass, PUGB4
			9'd98 : rdata = 43'b1100011100010000000000000000000000000001100;
			// PEs: 10 -> 32
			// srcs: (105, 99)(878) 608 --> (878) 608:PEGB2, pass, PUGB4
			9'd99 : rdata = 43'b1100011100100000000000000000000000000001100;
			// PEs: 11 -> 32
			// srcs: (106, 100)(908) -20 --> (908) -20:PEGB3, pass, PUGB4
			9'd100 : rdata = 43'b1100011100110000000000000000000000000001100;
			// PEs: 12 -> 32
			// srcs: (107, 101)(938) -87 --> (938) -87:PEGB4, pass, PUGB4
			9'd101 : rdata = 43'b1100011101000000000000000000000000000001100;
			// PEs: 13 -> 32
			// srcs: (108, 102)(968) 231 --> (968) 231:PEGB5, pass, PUGB4
			9'd102 : rdata = 43'b1100011101010000000000000000000000000001100;
			// PEs: 14 -> 32
			// srcs: (109, 103)(998) 0 --> (998) 0:PEGB6, pass, PUGB4
			9'd103 : rdata = 43'b1100011101100000000000000000000000000001100;
			// PEs: 15 -> 32
			// srcs: (110, 104)(1028) 990 --> (1028) 990:PENB, pass, PUGB4
			9'd104 : rdata = 43'b1100011011110000000000000000000000000001100;
			// PEs: 9 -> 32
			// srcs: (111, 105)(849) 320 --> (849) 320:PEGB1, pass, PUGB4
			9'd105 : rdata = 43'b1100011100010000000000000000000000000001100;
			// PEs: 10 -> 32
			// srcs: (112, 106)(879) 128 --> (879) 128:PEGB2, pass, PUGB4
			9'd106 : rdata = 43'b1100011100100000000000000000000000000001100;
			// PEs: 11 -> 32
			// srcs: (113, 107)(909) -37 --> (909) -37:PEGB3, pass, PUGB4
			9'd107 : rdata = 43'b1100011100110000000000000000000000000001100;
			// PEs: 12 -> 32
			// srcs: (114, 108)(939) 783 --> (939) 783:PEGB4, pass, PUGB4
			9'd108 : rdata = 43'b1100011101000000000000000000000000000001100;
			// PEs: 13 -> 32
			// srcs: (115, 109)(969) 858 --> (969) 858:PEGB5, pass, PUGB4
			9'd109 : rdata = 43'b1100011101010000000000000000000000000001100;
			// PEs: 14 -> 32
			// srcs: (116, 110)(999) 44 --> (999) 44:PEGB6, pass, PUGB4
			9'd110 : rdata = 43'b1100011101100000000000000000000000000001100;
			// PEs: 15 -> 32
			// srcs: (117, 111)(1029) -22 --> (1029) -22:PENB, pass, PUGB4
			9'd111 : rdata = 43'b1100011011110000000000000000000000000001100;
			// PEs: 9 -> 40
			// srcs: (118, 112)(850) 480 --> (850) 480:PEGB1, pass, PUGB5
			9'd112 : rdata = 43'b1100011100010000000000000000000000000001101;
			// PEs: 10 -> 40
			// srcs: (119, 113)(880) 704 --> (880) 704:PEGB2, pass, PUGB5
			9'd113 : rdata = 43'b1100011100100000000000000000000000000001101;
			// PEs: 11 -> 40
			// srcs: (120, 114)(910) -2 --> (910) -2:PEGB3, pass, PUGB5
			9'd114 : rdata = 43'b1100011100110000000000000000000000000001101;
			// PEs: 12 -> 40
			// srcs: (121, 115)(940) 348 --> (940) 348:PEGB4, pass, PUGB5
			9'd115 : rdata = 43'b1100011101000000000000000000000000000001101;
			// PEs: 13 -> 40
			// srcs: (122, 116)(970) 891 --> (970) 891:PEGB5, pass, PUGB5
			9'd116 : rdata = 43'b1100011101010000000000000000000000000001101;
			// PEs: 14 -> 40
			// srcs: (123, 117)(1000) 52 --> (1000) 52:PEGB6, pass, PUGB5
			9'd117 : rdata = 43'b1100011101100000000000000000000000000001101;
			// PEs: 15 -> 40
			// srcs: (124, 118)(1030) 462 --> (1030) 462:PENB, pass, PUGB5
			9'd118 : rdata = 43'b1100011011110000000000000000000000000001101;
			// PEs: 9 -> 48
			// srcs: (125, 119)(851) 320 --> (851) 320:PEGB1, pass, PUGB6
			9'd119 : rdata = 43'b1100011100010000000000000000000000000001110;
			// PEs: 10 -> 48
			// srcs: (126, 120)(881) 224 --> (881) 224:PEGB2, pass, PUGB6
			9'd120 : rdata = 43'b1100011100100000000000000000000000000001110;
			// PEs: 11 -> 48
			// srcs: (127, 121)(911) -14 --> (911) -14:PEGB3, pass, PUGB6
			9'd121 : rdata = 43'b1100011100110000000000000000000000000001110;
			// PEs: 12 -> 48
			// srcs: (128, 122)(941) 1334 --> (941) 1334:PEGB4, pass, PUGB6
			9'd122 : rdata = 43'b1100011101000000000000000000000000000001110;
			// PEs: 13 -> 48
			// srcs: (129, 123)(971) 1584 --> (971) 1584:PEGB5, pass, PUGB6
			9'd123 : rdata = 43'b1100011101010000000000000000000000000001110;
			// PEs: 14 -> 48
			// srcs: (130, 124)(1001) 30 --> (1001) 30:PEGB6, pass, PUGB6
			9'd124 : rdata = 43'b1100011101100000000000000000000000000001110;
			// PEs: 15 -> 48
			// srcs: (131, 125)(1031) -44 --> (1031) -44:PENB, pass, PUGB6
			9'd125 : rdata = 43'b1100011011110000000000000000000000000001110;
			// PEs: 9 -> 56
			// srcs: (132, 126)(852) 256 --> (852) 256:PEGB1, pass, PUGB7
			9'd126 : rdata = 43'b1100011100010000000000000000000000000001111;
			// PEs: 10 -> 56
			// srcs: (133, 127)(882) 576 --> (882) 576:PEGB2, pass, PUGB7
			9'd127 : rdata = 43'b1100011100100000000000000000000000000001111;
			// PEs: 11 -> 56
			// srcs: (134, 128)(912) -20 --> (912) -20:PEGB3, pass, PUGB7
			9'd128 : rdata = 43'b1100011100110000000000000000000000000001111;
			// PEs: 12 -> 0
			// srcs: (135, 129)(942) 1276 --> (942) 1276:PEGB4, pass, PUGB0
			9'd129 : rdata = 43'b1100011101000000000000000000000000000001000;
			// PEs: 13 -> 0
			// srcs: (136, 130)(972) 561 --> (972) 561:PEGB5, pass, PUGB0
			9'd130 : rdata = 43'b1100011101010000000000000000000000000001000;
			// PEs: 14 -> 0
			// srcs: (137, 131)(1002) 42 --> (1002) 42:PEGB6, pass, PUGB0
			9'd131 : rdata = 43'b1100011101100000000000000000000000000001000;
			// PEs: 15 -> 0
			// srcs: (138, 132)(1032) 594 --> (1032) 594:PENB, pass, PUGB0
			9'd132 : rdata = 43'b1100011011110000000000000000000000000001000;
			// PEs: 0 -> 8
			// srcs: (139, 133)(643) 266 --> (643) 266:PUNB, pass, NI0
			9'd133 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 0 -> 10
			// srcs: (140, 134)(673) 143 --> (673) 143:PUNB, pass, PEGB2
			9'd134 : rdata = 43'b1100011011111000000000000000000000010100000;
			// PEs: 9 -> 16
			// srcs: (141, 142)(853) 160 --> (853) 160:PEGB1, pass, PUNB
			9'd135 : rdata = 43'b1100011100010000000000000000000001000000000;
			// PEs: 10 -> 16
			// srcs: (142, 143)(883) -96 --> (883) -96:PEGB2, pass, PUNB
			9'd136 : rdata = 43'b1100011100100000000000000000000001000000000;
			// PEs: 11 -> 16
			// srcs: (143, 144)(913) -30 --> (913) -30:PEGB3, pass, PUNB
			9'd137 : rdata = 43'b1100011100110000000000000000000001000000000;
			// PEs: 12 -> 16
			// srcs: (144, 145)(943) 203 --> (943) 203:PEGB4, pass, PUNB
			9'd138 : rdata = 43'b1100011101000000000000000000000001000000000;
			// PEs: 13 -> 16
			// srcs: (145, 146)(973) 363 --> (973) 363:PEGB5, pass, PUNB
			9'd139 : rdata = 43'b1100011101010000000000000000000001000000000;
			// PEs: 14 -> 16
			// srcs: (146, 147)(1003) 94 --> (1003) 94:PEGB6, pass, PUNB
			9'd140 : rdata = 43'b1100011101100000000000000000000001000000000;
			// PEs: 15 -> 16
			// srcs: (147, 148)(1033) 638 --> (1033) 638:PENB, pass, PUNB
			9'd141 : rdata = 43'b1100011011110000000000000000000001000000000;
			// PEs: 16 -> 8
			// srcs: (148, 149)(1123) 851 --> (1123) 851:PUGB2, pass, NI1
			9'd142 : rdata = 43'b1100011100101000000001000010000000000000000;
			// PEs: 8 -> 10
			// srcs: (149, 135)(643) 266 --> (643) 266:NI0, pass, PEGB2
			9'd143 : rdata = 43'b1100010100000000000000000000000000010100000;
			// PEs: 0 -> 8
			// srcs: (150, 136)(703) 72 --> (703) 72:PUNB, pass, NI0
			9'd144 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 0 -> 10
			// srcs: (151, 137)(733) 460 --> (733) 460:PUNB, pass, PEGB2
			9'd145 : rdata = 43'b1100011011111000000000000000000000010100000;
			// PEs: 16 -> 9
			// srcs: (152, 150)(1153) 377 --> (1153) 377:PUGB2, pass, PENB
			9'd146 : rdata = 43'b1100011100101000000000000000000000100000000;
			// PEs: 10 -> 16
			// srcs: (153, 165)(884) 640 --> (884) 640:PEGB2, pass, PUNB
			9'd147 : rdata = 43'b1100011100100000000000000000000001000000000;
			// PEs: 11 -> 16
			// srcs: (154, 166)(914) -19 --> (914) -19:PEGB3, pass, PUNB
			9'd148 : rdata = 43'b1100011100110000000000000000000001000000000;
			// PEs: 12 -> 16
			// srcs: (155, 167)(944) 580 --> (944) 580:PEGB4, pass, PUNB
			9'd149 : rdata = 43'b1100011101000000000000000000000001000000000;
			// PEs: 13 -> 16
			// srcs: (156, 168)(974) 759 --> (974) 759:PEGB5, pass, PUNB
			9'd150 : rdata = 43'b1100011101010000000000000000000001000000000;
			// PEs: 14 -> 16
			// srcs: (157, 169)(1004) 32 --> (1004) 32:PEGB6, pass, PUNB
			9'd151 : rdata = 43'b1100011101100000000000000000000001000000000;
			// PEs: 8 -> 9
			// srcs: (158, 151)(1123) 851 --> (1123) 851:NI1, pass, PENB
			9'd152 : rdata = 43'b1100010100001000000000000000000000100000000;
			// PEs: 16 -> 8
			// srcs: (159, 152)(1183) 72 --> (1183) 72:PUGB2, pass, NI1
			9'd153 : rdata = 43'b1100011100101000000001000010000000000000000;
			// PEs: 8 -> 10
			// srcs: (160, 138)(703) 72 --> (703) 72:NI0, pass, PEGB2
			9'd154 : rdata = 43'b1100010100000000000000000000000000010100000;
			// PEs: 0 -> 8
			// srcs: (161, 139)(763) -72 --> (763) -72:PUNB, pass, NI0
			9'd155 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 0 -> 10
			// srcs: (162, 140)(793) 95 --> (793) 95:PUNB, pass, PEGB2
			9'd156 : rdata = 43'b1100011011111000000000000000000000010100000;
			// PEs: 16 -> 9
			// srcs: (163, 153)(1213) 775 --> (1213) 775:PUGB2, pass, PENB
			9'd157 : rdata = 43'b1100011100101000000000000000000000100000000;
			// PEs: 15 -> 16
			// srcs: (164, 170)(1034) 220 --> (1034) 220:PENB, pass, PUNB
			9'd158 : rdata = 43'b1100011011110000000000000000000001000000000;
			// PEs: 10 -> 16
			// srcs: (165, 181)(885) 128 --> (885) 128:PEGB2, pass, PUNB
			9'd159 : rdata = 43'b1100011100100000000000000000000001000000000;
			// PEs: 11 -> 16
			// srcs: (166, 182)(915) -2 --> (915) -2:PEGB3, pass, PUNB
			9'd160 : rdata = 43'b1100011100110000000000000000000001000000000;
			// PEs: 12 -> 16
			// srcs: (167, 183)(945) 87 --> (945) 87:PEGB4, pass, PUNB
			9'd161 : rdata = 43'b1100011101000000000000000000000001000000000;
			// PEs: 13 -> 16
			// srcs: (168, 184)(975) 1089 --> (975) 1089:PEGB5, pass, PUNB
			9'd162 : rdata = 43'b1100011101010000000000000000000001000000000;
			// PEs: 8 -> 9
			// srcs: (169, 154)(1183) 72 --> (1183) 72:NI1, pass, PENB
			9'd163 : rdata = 43'b1100010100001000000000000000000000100000000;
			// PEs: 0 -> 8
			// srcs: (170, 155)(644) 210 --> (644) 210:PUNB, pass, NI1
			9'd164 : rdata = 43'b1100011011111000000001000010000000000000000;
			// PEs: 8 -> 10
			// srcs: (171, 141)(763) -72 --> (763) -72:NI0, pass, PEGB2
			9'd165 : rdata = 43'b1100010100000000000000000000000000010100000;
			// PEs: 0 -> 9
			// srcs: (172, 156)(674) 132 --> (674) 132:PUNB, pass, PENB
			9'd166 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 14 -> 16
			// srcs: (173, 185)(1005) 44 --> (1005) 44:PEGB6, pass, PUNB
			9'd167 : rdata = 43'b1100011101100000000000000000000001000000000;
			// PEs: 15 -> 16
			// srcs: (174, 186)(1035) 330 --> (1035) 330:PENB, pass, PUNB
			9'd168 : rdata = 43'b1100011011110000000000000000000001000000000;
			// PEs: 10 -> 16
			// srcs: (175, 197)(886) 1024 --> (886) 1024:PEGB2, pass, PUNB
			9'd169 : rdata = 43'b1100011100100000000000000000000001000000000;
			// PEs: 11 -> 16
			// srcs: (176, 198)(916) -23 --> (916) -23:PEGB3, pass, PUNB
			9'd170 : rdata = 43'b1100011100110000000000000000000001000000000;
			// PEs: 12 -> 16
			// srcs: (177, 199)(946) 1421 --> (946) 1421:PEGB4, pass, PUNB
			9'd171 : rdata = 43'b1100011101000000000000000000000001000000000;
			// PEs: 8 -> 9
			// srcs: (178, 157)(644) 210 --> (644) 210:NI1, pass, PENB
			9'd172 : rdata = 43'b1100010100001000000000000000000000100000000;
			// PEs: 0 -> 8
			// srcs: (179, 158)(704) 120 --> (704) 120:PUNB, pass, NI0
			9'd173 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 0 -> 9
			// srcs: (180, 159)(734) 46 --> (734) 46:PUNB, pass, PENB
			9'd174 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 13 -> 16
			// srcs: (181, 200)(976) 891 --> (976) 891:PEGB5, pass, PUNB
			9'd175 : rdata = 43'b1100011101010000000000000000000001000000000;
			// PEs: 14 -> 16
			// srcs: (182, 201)(1006) 70 --> (1006) 70:PEGB6, pass, PUNB
			9'd176 : rdata = 43'b1100011101100000000000000000000001000000000;
			// PEs: 15 -> 16
			// srcs: (183, 202)(1036) 0 --> (1036) 0:PENB, pass, PUNB
			9'd177 : rdata = 43'b1100011011110000000000000000000001000000000;
			// PEs: 10 -> 16
			// srcs: (184, 213)(887) 128 --> (887) 128:PEGB2, pass, PUNB
			9'd178 : rdata = 43'b1100011100100000000000000000000001000000000;
			// PEs: 11 -> 16
			// srcs: (185, 214)(917) -39 --> (917) -39:PEGB3, pass, PUNB
			9'd179 : rdata = 43'b1100011100110000000000000000000001000000000;
			// PEs: 8 -> 9
			// srcs: (186, 160)(704) 120 --> (704) 120:NI0, pass, PENB
			9'd180 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 8
			// srcs: (187, 161)(764) 480 --> (764) 480:PUNB, pass, NI0
			9'd181 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 0 -> 9
			// srcs: (188, 162)(794) 798 --> (794) 798:PUNB, pass, PENB
			9'd182 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 0 -> 12
			// srcs: (189, 164)(824) 713 --> (824) 713:PUNB, pass, PEGB4
			9'd183 : rdata = 43'b1100011011111000000000000000000000011000000;
			// PEs: 12 -> 16
			// srcs: (190, 215)(947) 1015 --> (947) 1015:PEGB4, pass, PUNB
			9'd184 : rdata = 43'b1100011101000000000000000000000001000000000;
			// PEs: 13 -> 16
			// srcs: (191, 216)(977) 132 --> (977) 132:PEGB5, pass, PUNB
			9'd185 : rdata = 43'b1100011101010000000000000000000001000000000;
			// PEs: 14 -> 16
			// srcs: (192, 217)(1007) 72 --> (1007) 72:PEGB6, pass, PUNB
			9'd186 : rdata = 43'b1100011101100000000000000000000001000000000;
			// PEs: 15 -> 16
			// srcs: (193, 218)(1037) 220 --> (1037) 220:PENB, pass, PUNB
			9'd187 : rdata = 43'b1100011011110000000000000000000001000000000;
			// PEs: 8 -> 9
			// srcs: (194, 163)(764) 480 --> (764) 480:NI0, pass, PENB
			9'd188 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 8
			// srcs: (195, 171)(645) 98 --> (645) 98:PUNB, pass, NI0
			9'd189 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 0 -> 9
			// srcs: (196, 172)(675) 231 --> (675) 231:PUNB, pass, PENB
			9'd190 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 10 -> 16
			// srcs: (197, 228)(1587) 23 --> (1587) 23:PEGB2, pass, PUNB
			9'd191 : rdata = 43'b1100011100100000000000000000000001000000000;
			// PEs: 11 -> 16
			// srcs: (198, 233)(1686) 724 --> (1686) 724:PEGB3, pass, PUNB
			9'd192 : rdata = 43'b1100011100110000000000000000000001000000000;
			// PEs: 11 -> 16
			// srcs: (199, 235)(1705) 358 --> (1705) 358:PEGB3, pass, PUNB
			9'd193 : rdata = 43'b1100011100110000000000000000000001000000000;
			// PEs: 13 -> 16
			// srcs: (200, 237)(1724) 482 --> (1724) 482:PEGB5, pass, PUNB
			9'd194 : rdata = 43'b1100011101010000000000000000000001000000000;
			// PEs: 15 -> 16
			// srcs: (201, 239)(1743) 560 --> (1743) 560:PENB, pass, PUNB
			9'd195 : rdata = 43'b1100011011110000000000000000000001000000000;
			// PEs: 8 -> 9
			// srcs: (202, 173)(645) 98 --> (645) 98:NI0, pass, PENB
			9'd196 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 8
			// srcs: (203, 174)(705) 456 --> (705) 456:PUNB, pass, NI0
			9'd197 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 0 -> 9
			// srcs: (204, 175)(735) 1196 --> (735) 1196:PUNB, pass, PENB
			9'd198 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 15 -> 16
			// srcs: (205, 241)(1762) 102 --> (1762) 102:PENB, pass, PUNB
			9'd199 : rdata = 43'b1100011011110000000000000000000001000000000;
			// PEs: 15 -> 16
			// srcs: (206, 243)(1781) 536 --> (1781) 536:PENB, pass, PUNB
			9'd200 : rdata = 43'b1100011011110000000000000000000001000000000;
			// PEs: 9 -> 0
			// srcs: (207, 256)(1749) 1988 --> (1749) 1988:PEGB1, pass, PUGB0
			9'd201 : rdata = 43'b1100011100010000000000000000000000000001000;
			// PEs: 8 -> 9
			// srcs: (210, 176)(705) 456 --> (705) 456:NI0, pass, PENB
			9'd202 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 8
			// srcs: (211, 177)(765) 552 --> (765) 552:PUNB, pass, NI0
			9'd203 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 0 -> 9
			// srcs: (212, 178)(795) 209 --> (795) 209:PUNB, pass, PENB
			9'd204 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 0 -> 10
			// srcs: (213, 180)(825) 403 --> (825) 403:PUNB, pass, PEGB2
			9'd205 : rdata = 43'b1100011011111000000000000000000000010100000;
			// PEs: 10 -> 16
			// srcs: (214, 247)(1595) 941 --> (1595) 941:PEGB2, pass, PUNB
			9'd206 : rdata = 43'b1100011100100000000000000000000001000000000;
			// PEs: 8 -> 9
			// srcs: (218, 179)(765) 552 --> (765) 552:NI0, pass, PENB
			9'd207 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 8
			// srcs: (219, 187)(646) 420 --> (646) 420:PUNB, pass, NI0
			9'd208 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 0 -> 9
			// srcs: (220, 188)(676) 451 --> (676) 451:PUNB, pass, PENB
			9'd209 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 8 -> 9
			// srcs: (226, 189)(646) 420 --> (646) 420:NI0, pass, PENB
			9'd210 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 8
			// srcs: (227, 190)(706) 576 --> (706) 576:PUNB, pass, NI0
			9'd211 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 0 -> 9
			// srcs: (228, 191)(736) 1196 --> (736) 1196:PUNB, pass, PENB
			9'd212 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 8 -> 9
			// srcs: (234, 192)(706) 576 --> (706) 576:NI0, pass, PENB
			9'd213 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 8
			// srcs: (235, 193)(766) 504 --> (766) 504:PUNB, pass, NI0
			9'd214 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 0 -> 9
			// srcs: (236, 194)(796) 456 --> (796) 456:PUNB, pass, PENB
			9'd215 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 0 -> 10
			// srcs: (237, 196)(826) 248 --> (826) 248:PUNB, pass, PEGB2
			9'd216 : rdata = 43'b1100011011111000000000000000000000010100000;
			// PEs: 8 -> 9
			// srcs: (242, 195)(766) 504 --> (766) 504:NI0, pass, PENB
			9'd217 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 8
			// srcs: (243, 203)(647) 546 --> (647) 546:PUNB, pass, NI0
			9'd218 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 0 -> 9
			// srcs: (244, 204)(677) 121 --> (677) 121:PUNB, pass, PENB
			9'd219 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 8 -> 9
			// srcs: (250, 205)(647) 546 --> (647) 546:NI0, pass, PENB
			9'd220 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 8
			// srcs: (251, 206)(707) 120 --> (707) 120:PUNB, pass, NI0
			9'd221 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 0 -> 9
			// srcs: (252, 207)(737) 828 --> (737) 828:PUNB, pass, PENB
			9'd222 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 8 -> 9
			// srcs: (258, 208)(707) 120 --> (707) 120:NI0, pass, PENB
			9'd223 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 8
			// srcs: (259, 209)(767) 672 --> (767) 672:PUNB, pass, NI0
			9'd224 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 0 -> 9
			// srcs: (260, 210)(797) 399 --> (797) 399:PUNB, pass, PENB
			9'd225 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 8 -> 9
			// srcs: (266, 211)(767) 672 --> (767) 672:NI0, pass, PENB
			9'd226 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 9
			// srcs: (267, 212)(827) 217 --> (827) 217:PUNB, pass, PENB
			9'd227 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 0 -> 9
			// srcs: (268, 219)(828) 1271 --> (828) 1271:PUNB, pass, PENB
			9'd228 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 0 -> 10
			// srcs: (269, 220)(829) 992 --> (829) 992:PUNB, pass, PEGB2
			9'd229 : rdata = 43'b1100011011111000000000000000000000010100000;
			// PEs: 0 -> 9
			// srcs: (270, 221)(830) 806 --> (830) 806:PUNB, pass, PENB
			9'd230 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 0 -> 9
			// srcs: (271, 222)(831) 744 --> (831) 744:PUNB, pass, PENB
			9'd231 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 0 -> 10
			// srcs: (272, 223)(832) 341 --> (832) 341:PUNB, pass, PEGB2
			9'd232 : rdata = 43'b1100011011111000000000000000000000010100000;
			// PEs: 0 -> 9
			// srcs: (273, 224)(833) 465 --> (833) 465:PUNB, pass, PENB
			9'd233 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 32 -> 8
			// srcs: (274, 225)(1344) 60 --> (1344) 60:PUGB4, pass, NI0
			9'd234 : rdata = 43'b1100011101001000000001000000000000000000000;
			// PEs: 24 -> 9
			// srcs: (275, 226)(1345) 1815 --> (1345) 1815:PUGB3, pass, PENB
			9'd235 : rdata = 43'b1100011100111000000000000000000000100000000;
			// PEs: 9 -> 32
			// srcs: (278, 238)(1740) 2120 --> (1740) 2120:PEGB1, pass, PUGB4
			9'd236 : rdata = 43'b1100011100010000000000000000000000000001100;
			// PEs: 10 -> 24
			// srcs: (279, 234)(1702) 1312 --> (1702) 1312:PEGB2, pass, PUGB3
			9'd237 : rdata = 43'b1100011100100000000000000000000000000001011;
			// PEs: 9 -> 40
			// srcs: (280, 242)(1778) 1585 --> (1778) 1585:PEGB1, pass, PUGB5
			9'd238 : rdata = 43'b1100011100010000000000000000000000000001101;
			// PEs: 8 -> 9
			// srcs: (281, 227)(1344) 60 --> (1344) 60:NI0, pass, PENB
			9'd239 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 9 -> 40
			// srcs: (288, 251)(1351) 1875 --> (1351) 1875:PEGB1, pass, PUGB5
			9'd240 : rdata = 43'b1100011100010000000000000000000000000001101;
			// PEs: 16 -> 8
			// srcs: (325, 229)(1629) 374 --> (1629) 374:PUGB2, pass, NI0
			9'd241 : rdata = 43'b1100011100101000000001000000000000000000000;
			// PEs: 24 -> 9
			// srcs: (494, 230)(1630) 1473 --> (1630) 1473:PUGB3, pass, PENB
			9'd242 : rdata = 43'b1100011100111000000000000000000000100000000;
			// PEs: 8 -> 9
			// srcs: (501, 231)(1629) 374 --> (1629) 374:NI0, pass, PENB
			9'd243 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 9
			// srcs: (502, 232)(1682) 1636 --> (1682) 1636:PUNB, pass, PENB
			9'd244 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 0 -> 9
			// srcs: (503, 236)(1720) 613 --> (1720) 613:PUNB, pass, PENB
			9'd245 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 0 -> 9
			// srcs: (504, 240)(1758) 1534 --> (1758) 1534:PUNB, pass, PENB
			9'd246 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 32 -> 8
			// srcs: (505, 244)(1291) 1070 --> (1291) 1070:PUGB4, pass, NI0
			9'd247 : rdata = 43'b1100011101001000000001000000000000000000000;
			// PEs: 40 -> 9
			// srcs: (506, 245)(1292) 3317 --> (1292) 3317:PUGB5, pass, PENB
			9'd248 : rdata = 43'b1100011101011000000000000000000000100000000;
			// PEs: 9 -> 16
			// srcs: (508, 252)(1636) 1847 --> (1636) 1847:PEGB1, pass, PUNB
			9'd249 : rdata = 43'b1100011100010000000000000000000001000000000;
			// PEs: 9 -> 32
			// srcs: (509, 248)(1691) 4091 --> (1691) 4091:PEGB1, pass, PUGB4
			9'd250 : rdata = 43'b1100011100010000000000000000000000000001100;
			// PEs: 15 -> 16
			// srcs: (510, 253)(1692) 1410 --> (1692) 1410:PENB, pass, PUNB
			9'd251 : rdata = 43'b1100011011110000000000000000000001000000000;
			// PEs: 11 -> 16
			// srcs: (511, 254)(1711) 1614 --> (1711) 1614:PEGB3, pass, PUNB
			9'd252 : rdata = 43'b1100011100110000000000000000000001000000000;
			// PEs: 8 -> 9
			// srcs: (512, 246)(1291) 1070 --> (1291) 1070:NI0, pass, PENB
			9'd253 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 9
			// srcs: (513, 249)(1728) 2715 --> (1728) 2715:PUNB, pass, PENB
			9'd254 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 0 -> 9
			// srcs: (514, 250)(1766) 3199 --> (1766) 3199:PUNB, pass, PENB
			9'd255 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 11 -> 16
			// srcs: (522, 255)(1730) 2549 --> (1730) 2549:PEGB3, pass, PUNB
			9'd256 : rdata = 43'b1100011100110000000000000000000001000000000;
			// PEs: 10 -> 16
			// srcs: (523, 257)(1768) 3151 --> (1768) 3151:PEGB2, pass, PUNB
			9'd257 : rdata = 43'b1100011100100000000000000000000001000000000;
			// PEs: 13 -> 16
			// srcs: (524, 258)(1787) 2303 --> (1787) 2303:PEGB5, pass, PUNB
			9'd258 : rdata = 43'b1100011101010000000000000000000001000000000;
			// PEs: 10 -> 16
			// srcs: (525, 269)(1599) 2075 --> (1599) 2075:PEGB2, pass, PUNB
			9'd259 : rdata = 43'b1100011100100000000000000000000001000000000;
			// PEs: 9 -> 32
			// srcs: (526, 270)(1619) 3843 --> (1619) 3843:PEGB1, pass, PUGB4
			9'd260 : rdata = 43'b1100011100010000000000000000000000000001100;
			// PEs: 10 -> 32
			// srcs: (534, 271)(1638) 3081 --> (1638) 3081:PEGB2, pass, PUGB4
			9'd261 : rdata = 43'b1100011100100000000000000000000000000001100;
			// PEs: 9 -> 16
			// srcs: (535, 274)(1733) 5670 --> (1733) 5670:PEGB1, pass, PUNB
			9'd262 : rdata = 43'b1100011100010000000000000000000001000000000;
			// PEs: 10 -> 32
			// srcs: (542, 272)(1657) 4043 --> (1657) 4043:PEGB2, pass, PUGB4
			9'd263 : rdata = 43'b1100011100100000000000000000000000000001100;
			// PEs: 9 -> 16
			// srcs: (543, 275)(1771) 6226 --> (1771) 6226:PEGB1, pass, PUNB
			9'd264 : rdata = 43'b1100011100010000000000000000000001000000000;
			// PEs: 9 -> 32
			// srcs: (550, 273)(1676) 3447 --> (1676) 3447:PEGB1, pass, PUGB4
			9'd265 : rdata = 43'b1100011100010000000000000000000000000001100;
			// PEs: 40 -> 9
			// srcs: (607, 259)(1295) 2557 --> (1295) 2557:PUGB5, pass, PENB
			9'd266 : rdata = 43'b1100011101011000000000000000000000100000000;
			// PEs: 9 -> 32
			// srcs: (614, 276)(1298) 6944 --> (1298) 6944:PEGB1, pass, PUGB4
			9'd267 : rdata = 43'b1100011100010000000000000000000000000001100;
			// PEs: 24 -> 8
			// srcs: (848, 260)(1314) 3020 --> (1314) 3020:PUGB3, pass, NI0
			9'd268 : rdata = 43'b1100011100111000000001000000000000000000000;
			// PEs: 48 -> 9
			// srcs: (849, 261)(1315) 4919 --> (1315) 4919:PUGB6, pass, PENB
			9'd269 : rdata = 43'b1100011101101000000000000000000000100000000;
			// PEs: 8 -> 9
			// srcs: (855, 262)(1314) 3020 --> (1314) 3020:NI0, pass, PENB
			9'd270 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 24 -> 8
			// srcs: (856, 263)(1390) 1954 --> (1390) 1954:PUGB3, pass, NI0
			9'd271 : rdata = 43'b1100011100111000000001000000000000000000000;
			// PEs: 48 -> 9
			// srcs: (857, 264)(1391) 5170 --> (1391) 5170:PUGB6, pass, PENB
			9'd272 : rdata = 43'b1100011101101000000000000000000000100000000;
			// PEs: 9 -> 32
			// srcs: (862, 277)(1317) 7939 --> (1317) 7939:PEGB1, pass, PUGB4
			9'd273 : rdata = 43'b1100011100010000000000000000000000000001100;
			// PEs: 8 -> 9
			// srcs: (863, 265)(1390) 1954 --> (1390) 1954:NI0, pass, PENB
			9'd274 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 24 -> 8
			// srcs: (864, 266)(1428) 1960 --> (1428) 1960:PUGB3, pass, NI0
			9'd275 : rdata = 43'b1100011100111000000001000000000000000000000;
			// PEs: 40 -> 9
			// srcs: (865, 267)(1429) 4852 --> (1429) 4852:PUGB5, pass, PENB
			9'd276 : rdata = 43'b1100011101011000000000000000000000100000000;
			// PEs: 8 -> 9
			// srcs: (871, 268)(1428) 1960 --> (1428) 1960:NI0, pass, PENB
			9'd277 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 16 -> 9
			// srcs: (872, 278)(1392) 2905 --> (1392) 2905:PUGB2, pass, PENB
			9'd278 : rdata = 43'b1100011100101000000000000000000000100000000;
			// PEs: 9 -> 40
			// srcs: (878, 279)(1431) 6812 --> (1431) 6812:PEGB1, pass, PUGB5
			9'd279 : rdata = 43'b1100011100010000000000000000000000000001101;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 9) begin
	always @(*) begin
		case(address)
			// PEs: 9, 9 -> 8
			// srcs: (1, 0)(234) 31, (11) 32 --> (834) 992:NW0, ND0, *, PEGB0
			9'd0 : rdata = 43'b0001101000000011000000000000000000010000000;
			// PEs: 9, 9 -> 8
			// srcs: (2, 1)(235) 1, (11) 32 --> (835) 32:NW1, ND0, *, PEGB0
			9'd1 : rdata = 43'b0001101000001011000000000000000000010000000;
			// PEs: 9, 9 -> 8
			// srcs: (3, 2)(236) 21, (11) 32 --> (836) 672:NW2, ND0, *, PEGB0
			9'd2 : rdata = 43'b0001101000010011000000000000000000010000000;
			// PEs: 9, 9 -> 8
			// srcs: (4, 3)(237) 45, (11) 32 --> (837) 1440:NW3, ND0, *, PEGB0
			9'd3 : rdata = 43'b0001101000011011000000000000000000010000000;
			// PEs: 9, 9 -> 8
			// srcs: (5, 4)(238) 8, (11) 32 --> (838) 256:NW4, ND0, *, PEGB0
			9'd4 : rdata = 43'b0001101000100011000000000000000000010000000;
			// PEs: 9, 9 -> 8
			// srcs: (6, 5)(239) 23, (11) 32 --> (839) 736:NW5, ND0, *, PEGB0
			9'd5 : rdata = 43'b0001101000101011000000000000000000010000000;
			// PEs: 9, 9 -> 8
			// srcs: (7, 6)(240) 2, (11) 32 --> (840) 64:NW6, ND0, *, PEGB0
			9'd6 : rdata = 43'b0001101000110011000000000000000000010000000;
			// PEs: 9, 9 -> 8
			// srcs: (8, 7)(241) -3, (11) 32 --> (841) -96:NW7, ND0, *, PEGB0
			9'd7 : rdata = 43'b0001101000111011000000000000000000010000000;
			// PEs: 9, 9 -> 8
			// srcs: (9, 8)(242) 13, (11) 32 --> (842) 416:NW8, ND0, *, PEGB0
			9'd8 : rdata = 43'b0001101001000011000000000000000000010000000;
			// PEs: 9, 9 -> 8
			// srcs: (10, 9)(243) 42, (11) 32 --> (843) 1344:NW9, ND0, *, PEGB0
			9'd9 : rdata = 43'b0001101001001011000000000000000000010000000;
			// PEs: 9, 9 -> 8
			// srcs: (11, 10)(244) 5, (11) 32 --> (844) 160:NW10, ND0, *, PEGB0
			9'd10 : rdata = 43'b0001101001010011000000000000000000010000000;
			// PEs: 9, 9 -> 8
			// srcs: (12, 11)(245) 21, (11) 32 --> (845) 672:NW11, ND0, *, PEGB0
			9'd11 : rdata = 43'b0001101001011011000000000000000000010000000;
			// PEs: 9, 9 -> 8
			// srcs: (13, 12)(246) 14, (11) 32 --> (846) 448:NW12, ND0, *, PEGB0
			9'd12 : rdata = 43'b0001101001100011000000000000000000010000000;
			// PEs: 9, 9 -> 8
			// srcs: (14, 13)(247) 49, (11) 32 --> (847) 1568:NW13, ND0, *, PEGB0
			9'd13 : rdata = 43'b0001101001101011000000000000000000010000000;
			// PEs: 9, 9 -> 8
			// srcs: (15, 14)(248) 27, (11) 32 --> (848) 864:NW14, ND0, *, PEGB0
			9'd14 : rdata = 43'b0001101001110011000000000000000000010000000;
			// PEs: 9, 9 -> 8
			// srcs: (16, 15)(249) 10, (11) 32 --> (849) 320:NW15, ND0, *, PEGB0
			9'd15 : rdata = 43'b0001101001111011000000000000000000010000000;
			// PEs: 9, 9 -> 8
			// srcs: (17, 16)(250) 15, (11) 32 --> (850) 480:NW16, ND0, *, PEGB0
			9'd16 : rdata = 43'b0001101010000011000000000000000000010000000;
			// PEs: 9, 9 -> 8
			// srcs: (18, 17)(251) 10, (11) 32 --> (851) 320:NW17, ND0, *, PEGB0
			9'd17 : rdata = 43'b0001101010001011000000000000000000010000000;
			// PEs: 9, 9 -> 8
			// srcs: (19, 18)(252) 8, (11) 32 --> (852) 256:NW18, ND0, *, PEGB0
			9'd18 : rdata = 43'b0001101010010011000000000000000000010000000;
			// PEs: 9, 9 -> 8
			// srcs: (20, 19)(253) 5, (11) 32 --> (853) 160:NW19, ND0, *, PEGB0
			9'd19 : rdata = 43'b0001101010011011000000000000000000010000000;
			// PEs: 9, 9 -> 12
			// srcs: (21, 20)(254) 42, (11) 32 --> (854) 1344:NW20, ND0, *, PEGB4
			9'd20 : rdata = 43'b0001101010100011000000000000000000011000000;
			// PEs: 9, 9 -> 10
			// srcs: (22, 21)(255) -2, (11) 32 --> (855) -64:NW21, ND0, *, PENB
			9'd21 : rdata = 43'b0001101010101011000000000000000000100000000;
			// PEs: 9, 9 -> 10
			// srcs: (23, 22)(256) 6, (11) 32 --> (856) 192:NW22, ND0, *, PENB
			9'd22 : rdata = 43'b0001101010110011000000000000000000100000000;
			// PEs: 9, 9 -> 9
			// srcs: (24, 23)(257) 17, (11) 32 --> (857) 544:NW23, ND0, *, NI0
			9'd23 : rdata = 43'b0001101010111011000001000000000000000000000;
			// PEs: 9, 9 -> 9
			// srcs: (25, 24)(258) 37, (11) 32 --> (858) 1184:NW24, ND0, *, NI1
			9'd24 : rdata = 43'b0001101011000011000001000010000000000000000;
			// PEs: 9, 9 -> 10
			// srcs: (26, 25)(259) 10, (11) 32 --> (859) 320:NW25, ND0, *, PENB
			9'd25 : rdata = 43'b0001101011001011000000000000000000100000000;
			// PEs: 9, 9 -> 9
			// srcs: (27, 26)(260) 48, (11) 32 --> (860) 1536:NW26, ND0, *, NI2
			9'd26 : rdata = 43'b0001101011010011000001000100000000000000000;
			// PEs: 9, 9 -> 9
			// srcs: (28, 27)(261) 43, (11) 32 --> (861) 1376:NW27, ND0, *, NI3
			9'd27 : rdata = 43'b0001101011011011000001000110000000000000000;
			// PEs: 9, 9 -> 10
			// srcs: (29, 28)(262) 36, (11) 32 --> (862) 1152:NW28, ND0, *, PENB
			9'd28 : rdata = 43'b0001101011100011000000000000000000100000000;
			// PEs: 9, 9 -> 9
			// srcs: (30, 29)(263) 35, (11) 32 --> (863) 1120:NW29, ND0, *, NI4
			9'd29 : rdata = 43'b0001101011101011000001001000000000000000000;
			// PEs: 11 -> 9
			// srcs: (31, 60)(918) -2 --> (918) -2:PEGB3, pass, NI5
			9'd30 : rdata = 43'b1100011100110000000001001010000000000000000;
			// PEs: 11 -> 9
			// srcs: (32, 62)(919) -21 --> (919) -21:PEGB3, pass, NI6
			9'd31 : rdata = 43'b1100011100110000000001001100000000000000000;
			// PEs: 10, 9 -> 15
			// srcs: (33, 61)(888) -32, (918) -2 --> (1684) -34:PEGB2, NI5, +, PEGB7
			9'd32 : rdata = 43'b0000111100100101001010000000000000011110000;
			// PEs: 11 -> 9
			// srcs: (34, 66)(921) -10 --> (921) -10:PEGB3, pass, NI5
			9'd33 : rdata = 43'b1100011100110000000001001010000000000000000;
			// PEs: 11 -> 9
			// srcs: (35, 68)(922) -26 --> (922) -26:PEGB3, pass, NI7
			9'd34 : rdata = 43'b1100011100110000000001001110000000000000000;
			// PEs: 10, 9 -> 11
			// srcs: (36, 63)(889) 576, (919) -21 --> (1703) 555:PEGB2, NI6, +, PEGB3
			9'd35 : rdata = 43'b0000111100100101001100000000000000010110000;
			// PEs: 10, 9 -> 9
			// srcs: (39, 67)(891) 544, (921) -10 --> (1741) 534:PEGB2, NI5, +, NI6
			9'd36 : rdata = 43'b0000111100100101001011001100000000000000000;
			// PEs: 10, 9 -> 9
			// srcs: (42, 69)(892) 1088, (922) -26 --> (1760) 1062:PEGB2, NI7, +, NI5
			9'd37 : rdata = 43'b0000111100100101001111001010000000000000000;
			// PEs: 9, 13 -> 8
			// srcs: (45, 83)(1741) 534, (1742) 1454 --> (1749) 1988:NI6, PEGB5, +, PEGB0
			9'd38 : rdata = 43'b0000110100110111010100000000000000010000000;
			// PEs: 8 -> 
			// srcs: (154, 30)(1153) 377 --> (1153) 377:PENB, pass, 
			9'd39 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 8, 9 -> 9
			// srcs: (160, 31)(1123) 851, (1153) 377 --> (1593) 1228:PENB, ALU, +, NI6
			9'd40 : rdata = 43'b0000111011110001111111001100000000000000000;
			// PEs: 8 -> 
			// srcs: (165, 32)(1213) 775 --> (1213) 775:PENB, pass, 
			9'd41 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 8, 9 -> 9
			// srcs: (171, 33)(1183) 72, (1213) 775 --> (1594) 847:PENB, ALU, +, NI7
			9'd42 : rdata = 43'b0000111011110001111111001110000000000000000;
			// PEs: 8 -> 
			// srcs: (174, 34)(674) 132 --> (674) 132:PENB, pass, 
			9'd43 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 8, 9 -> 9
			// srcs: (180, 35)(644) 210, (674) 132 --> (1604) 342:PENB, ALU, +, NI8
			9'd44 : rdata = 43'b0000111011110001111111010000000000000000000;
			// PEs: 8 -> 
			// srcs: (182, 36)(734) 46 --> (734) 46:PENB, pass, 
			9'd45 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 8, 9 -> 9
			// srcs: (188, 37)(704) 120, (734) 46 --> (1605) 166:PENB, ALU, +, NI9
			9'd46 : rdata = 43'b0000111011110001111111010010000000000000000;
			// PEs: 8 -> 9
			// srcs: (190, 38)(794) 798 --> (794) 798:PENB, pass, NI10
			9'd47 : rdata = 43'b1100011011110000000001010100000000000000000;
			// PEs: 9 -> 9
			// srcs: (191, 108)(1604) 342 --> (1604) 342:NI8, pass, NI8
			9'd48 : rdata = 43'b1100010101000000000001010000000000000000000;
			// PEs: 9, 9 -> 9
			// srcs: (191, 73)(1604) 342, (1605) 166 --> (1614) 508:ALU, NI9, +, NI11
			9'd49 : rdata = 43'b0000100111111101010011010110000000000000000;
			// PEs: 8, 9 -> 9
			// srcs: (196, 39)(764) 480, (794) 798 --> (1606) 1278:PENB, NI10, +, NI8
			9'd50 : rdata = 43'b0000111011110101010101010000000000000000000;
			// PEs: 8 -> 9
			// srcs: (198, 40)(675) 231 --> (675) 231:PENB, pass, NI9
			9'd51 : rdata = 43'b1100011011110000000001010010000000000000000;
			// PEs: 9, 12 -> 9
			// srcs: (202, 74)(1606) 1278, (1607) 2057 --> (1615) 3335:NI8, PEGB4, +, NI10
			9'd52 : rdata = 43'b0000110101000111010001010100000000000000000;
			// PEs: 8, 9 -> 9
			// srcs: (204, 41)(645) 98, (675) 231 --> (1623) 329:PENB, NI9, +, NI8
			9'd53 : rdata = 43'b0000111011110101010011010000000000000000000;
			// PEs: 9 -> 9
			// srcs: (205, 109)(1614) 508 --> (1614) 508:NI11, pass, NI11
			9'd54 : rdata = 43'b1100010101011000000001010110000000000000000;
			// PEs: 9, 9 -> 9
			// srcs: (205, 90)(1614) 508, (1615) 3335 --> (1619) 3843:ALU, NI10, +, NI9
			9'd55 : rdata = 43'b0000100111111101010101010010000000000000000;
			// PEs: 8 -> 
			// srcs: (206, 42)(735) 1196 --> (735) 1196:PENB, pass, 
			9'd56 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 8, 9 -> 9
			// srcs: (212, 43)(705) 456, (735) 1196 --> (1624) 1652:PENB, ALU, +, NI10
			9'd57 : rdata = 43'b0000111011110001111111010100000000000000000;
			// PEs: 8 -> 9
			// srcs: (214, 44)(795) 209 --> (795) 209:PENB, pass, NI11
			9'd58 : rdata = 43'b1100011011110000000001010110000000000000000;
			// PEs: 9 -> 9
			// srcs: (215, 110)(1623) 329 --> (1623) 329:NI8, pass, NI8
			9'd59 : rdata = 43'b1100010101000000000001010000000000000000000;
			// PEs: 9, 9 -> 9
			// srcs: (215, 75)(1623) 329, (1624) 1652 --> (1633) 1981:ALU, NI10, +, NI12
			9'd60 : rdata = 43'b0000100111111101010101011000000000000000000;
			// PEs: 8, 9 -> 10
			// srcs: (220, 45)(765) 552, (795) 209 --> (1625) 761:PENB, NI11, +, PENB
			9'd61 : rdata = 43'b0000111011110101010110000000000000100000000;
			// PEs: 8 -> 
			// srcs: (222, 46)(676) 451 --> (676) 451:PENB, pass, 
			9'd62 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 8, 9 -> 9
			// srcs: (228, 47)(646) 420, (676) 451 --> (1642) 871:PENB, ALU, +, NI8
			9'd63 : rdata = 43'b0000111011110001111111010000000000000000000;
			// PEs: 8 -> 
			// srcs: (230, 48)(736) 1196 --> (736) 1196:PENB, pass, 
			9'd64 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 8, 9 -> 9
			// srcs: (236, 49)(706) 576, (736) 1196 --> (1643) 1772:PENB, ALU, +, NI10
			9'd65 : rdata = 43'b0000111011110001111111010100000000000000000;
			// PEs: 8 -> 9
			// srcs: (238, 50)(796) 456 --> (796) 456:PENB, pass, NI11
			9'd66 : rdata = 43'b1100011011110000000001010110000000000000000;
			// PEs: 9 -> 9
			// srcs: (239, 111)(1642) 871 --> (1642) 871:NI8, pass, NI8
			9'd67 : rdata = 43'b1100010101000000000001010000000000000000000;
			// PEs: 9, 9 -> 9
			// srcs: (239, 78)(1642) 871, (1643) 1772 --> (1652) 2643:ALU, NI10, +, NI13
			9'd68 : rdata = 43'b0000100111111101010101011010000000000000000;
			// PEs: 8, 9 -> 10
			// srcs: (244, 51)(766) 504, (796) 456 --> (1644) 960:PENB, NI11, +, PENB
			9'd69 : rdata = 43'b0000111011110101010110000000000000100000000;
			// PEs: 8 -> 
			// srcs: (246, 52)(677) 121 --> (677) 121:PENB, pass, 
			9'd70 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 8, 9 -> 9
			// srcs: (252, 53)(647) 546, (677) 121 --> (1661) 667:PENB, ALU, +, NI8
			9'd71 : rdata = 43'b0000111011110001111111010000000000000000000;
			// PEs: 8 -> 
			// srcs: (254, 54)(737) 828 --> (737) 828:PENB, pass, 
			9'd72 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 8, 9 -> 9
			// srcs: (260, 55)(707) 120, (737) 828 --> (1662) 948:PENB, ALU, +, NI10
			9'd73 : rdata = 43'b0000111011110001111111010100000000000000000;
			// PEs: 8 -> 9
			// srcs: (262, 56)(797) 399 --> (797) 399:PENB, pass, NI11
			9'd74 : rdata = 43'b1100011011110000000001010110000000000000000;
			// PEs: 9 -> 9
			// srcs: (263, 112)(1661) 667 --> (1661) 667:NI8, pass, NI8
			9'd75 : rdata = 43'b1100010101000000000001010000000000000000000;
			// PEs: 9, 9 -> 9
			// srcs: (263, 79)(1661) 667, (1662) 948 --> (1671) 1615:ALU, NI10, +, NI14
			9'd76 : rdata = 43'b0000100111111101010101011100000000000000000;
			// PEs: 8, 9 -> 9
			// srcs: (268, 57)(767) 672, (797) 399 --> (1663) 1071:PENB, NI11, +, NI8
			9'd77 : rdata = 43'b0000111011110101010111010000000000000000000;
			// PEs: 8, 9 -> 10
			// srcs: (269, 58)(827) 217, (857) 544 --> (1664) 761:PENB, NI0, +, PENB
			9'd78 : rdata = 43'b0000111011110101000000000000000000100000000;
			// PEs: 8, 9 -> 9
			// srcs: (270, 59)(828) 1271, (858) 1184 --> (1683) 2455:PENB, NI1, +, NI0
			9'd79 : rdata = 43'b0000111011110101000011000000000000000000000;
			// PEs: 8, 9 -> 9
			// srcs: (272, 64)(830) 806, (860) 1536 --> (1721) 2342:PENB, NI2, +, NI1
			9'd80 : rdata = 43'b0000111011110101000101000010000000000000000;
			// PEs: 8, 9 -> 8
			// srcs: (273, 65)(831) 744, (861) 1376 --> (1740) 2120:PENB, NI3, +, PEGB0
			9'd81 : rdata = 43'b0000111011110101000110000000000000010000000;
			// PEs: 8, 9 -> 8
			// srcs: (275, 70)(833) 465, (863) 1120 --> (1778) 1585:PENB, NI4, +, PEGB0
			9'd82 : rdata = 43'b0000111011110101001000000000000000010000000;
			// PEs: 8 -> 
			// srcs: (277, 71)(1345) 1815 --> (1345) 1815:PENB, pass, 
			9'd83 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 8, 9 -> 8
			// srcs: (283, 72)(1344) 60, (1345) 1815 --> (1351) 1875:PENB, ALU, +, PEGB0
			9'd84 : rdata = 43'b0000111011110001111110000000000000010000000;
			// PEs: 9 -> 10
			// srcs: (284, 80)(1663) 1071 --> (1663) 1071:NI8, pass, PENB
			9'd85 : rdata = 43'b1100010101000000000000000000000000100000000;
			// PEs: 9 -> 10
			// srcs: (285, 85)(1760) 1062 --> (1760) 1062:NI5, pass, PENB
			9'd86 : rdata = 43'b1100010100101000000000000000000000100000000;
			// PEs: 9 -> 10
			// srcs: (286, 86)(1594) 847 --> (1594) 847:NI7, pass, PENB
			9'd87 : rdata = 43'b1100010100111000000000000000000000100000000;
			// PEs: 9 -> 10
			// srcs: (287, 91)(1633) 1981 --> (1633) 1981:NI12, pass, PENB
			9'd88 : rdata = 43'b1100010101100000000000000000000000100000000;
			// PEs: 9 -> 10
			// srcs: (288, 92)(1652) 2643 --> (1652) 2643:NI13, pass, PENB
			9'd89 : rdata = 43'b1100010101101000000000000000000000100000000;
			// PEs: 9 -> 10
			// srcs: (403, 87)(1593) 1228 --> (1593) 1228:NI6, pass, PENB
			9'd90 : rdata = 43'b1100010100110000000000000000000000100000000;
			// PEs: 8 -> 
			// srcs: (496, 76)(1630) 1473 --> (1630) 1473:PENB, pass, 
			9'd91 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 8, 9 -> 8
			// srcs: (503, 77)(1629) 374, (1630) 1473 --> (1636) 1847:PENB, ALU, +, PEGB0
			9'd92 : rdata = 43'b0000111011110001111110000000000000010000000;
			// PEs: 8, 9 -> 8
			// srcs: (504, 81)(1682) 1636, (1683) 2455 --> (1691) 4091:PENB, NI0, +, PEGB0
			9'd93 : rdata = 43'b0000111011110101000000000000000000010000000;
			// PEs: 8, 9 -> 9
			// srcs: (505, 82)(1720) 613, (1721) 2342 --> (1729) 2955:PENB, NI1, +, NI0
			9'd94 : rdata = 43'b0000111011110101000011000000000000000000000;
			// PEs: 8, 10 -> 9
			// srcs: (506, 84)(1758) 1534, (1759) 1493 --> (1767) 3027:PENB, PEGB2, +, NI1
			9'd95 : rdata = 43'b0000111011110111001001000010000000000000000;
			// PEs: 9, 10 -> 9
			// srcs: (507, 93)(1671) 1615, (1672) 1832 --> (1676) 3447:NI14, PEGB2, +, NI2
			9'd96 : rdata = 43'b0000110101110111001001000100000000000000000;
			// PEs: 8 -> 
			// srcs: (508, 88)(1292) 3317 --> (1292) 3317:PENB, pass, 
			9'd97 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 8, 9 -> 9
			// srcs: (514, 89)(1291) 1070, (1292) 3317 --> (1296) 4387:PENB, ALU, +, NI3
			9'd98 : rdata = 43'b0000111011110001111111000110000000000000000;
			// PEs: 8, 9 -> 9
			// srcs: (515, 94)(1728) 2715, (1729) 2955 --> (1733) 5670:PENB, NI0, +, NI4
			9'd99 : rdata = 43'b0000111011110101000001001000000000000000000;
			// PEs: 8, 9 -> 9
			// srcs: (516, 95)(1766) 3199, (1767) 3027 --> (1771) 6226:PENB, NI1, +, NI0
			9'd100 : rdata = 43'b0000111011110101000011000000000000000000000;
			// PEs: 9 -> 8
			// srcs: (517, 103)(1619) 3843 --> (1619) 3843:NI9, pass, PEGB0
			9'd101 : rdata = 43'b1100010101001000000000000000000000010000000;
			// PEs: 9 -> 8
			// srcs: (529, 105)(1733) 5670 --> (1733) 5670:NI4, pass, PEGB0
			9'd102 : rdata = 43'b1100010100100000000000000000000000010000000;
			// PEs: 9 -> 8
			// srcs: (538, 106)(1771) 6226 --> (1771) 6226:NI0, pass, PEGB0
			9'd103 : rdata = 43'b1100010100000000000000000000000000010000000;
			// PEs: 9 -> 8
			// srcs: (545, 104)(1676) 3447 --> (1676) 3447:NI2, pass, PEGB0
			9'd104 : rdata = 43'b1100010100010000000000000000000000010000000;
			// PEs: 8, 9 -> 8
			// srcs: (609, 96)(1295) 2557, (1296) 4387 --> (1298) 6944:PENB, NI3, +, PEGB0
			9'd105 : rdata = 43'b0000111011110101000110000000000000010000000;
			// PEs: 8 -> 
			// srcs: (851, 97)(1315) 4919 --> (1315) 4919:PENB, pass, 
			9'd106 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 8, 9 -> 8
			// srcs: (857, 98)(1314) 3020, (1315) 4919 --> (1317) 7939:PENB, ALU, +, PEGB0
			9'd107 : rdata = 43'b0000111011110001111110000000000000010000000;
			// PEs: 8 -> 
			// srcs: (859, 99)(1391) 5170 --> (1391) 5170:PENB, pass, 
			9'd108 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 8, 9 -> 9
			// srcs: (865, 100)(1390) 1954, (1391) 5170 --> (1393) 7124:PENB, ALU, +, NI0
			9'd109 : rdata = 43'b0000111011110001111111000000000000000000000;
			// PEs: 8 -> 
			// srcs: (867, 101)(1429) 4852 --> (1429) 4852:PENB, pass, 
			9'd110 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 8, 9 -> 8
			// srcs: (873, 102)(1428) 1960, (1429) 4852 --> (1431) 6812:PENB, ALU, +, PEGB0
			9'd111 : rdata = 43'b0000111011110001111110000000000000010000000;
			// PEs: 8, 9 -> 9
			// srcs: (875, 107)(1392) 2905, (1393) 7124 --> (1394) 10029:PENB, NI0, +, NW30
			9'd112 : rdata = 43'b0000111011110101000000000001111100000000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 10) begin
	always @(*) begin
		case(address)
			// PEs: 10, 10 -> 8
			// srcs: (1, 0)(264) 38, (12) 32 --> (864) 1216:NW0, ND0, *, PEGB0
			9'd0 : rdata = 43'b0001101000000011000000000000000000010000000;
			// PEs: 10, 10 -> 8
			// srcs: (2, 1)(265) 41, (12) 32 --> (865) 1312:NW1, ND0, *, PEGB0
			9'd1 : rdata = 43'b0001101000001011000000000000000000010000000;
			// PEs: 10, 10 -> 8
			// srcs: (3, 2)(266) 13, (12) 32 --> (866) 416:NW2, ND0, *, PEGB0
			9'd2 : rdata = 43'b0001101000010011000000000000000000010000000;
			// PEs: 10, 10 -> 8
			// srcs: (4, 3)(267) 28, (12) 32 --> (867) 896:NW3, ND0, *, PEGB0
			9'd3 : rdata = 43'b0001101000011011000000000000000000010000000;
			// PEs: 10, 10 -> 8
			// srcs: (5, 4)(268) 1, (12) 32 --> (868) 32:NW4, ND0, *, PEGB0
			9'd4 : rdata = 43'b0001101000100011000000000000000000010000000;
			// PEs: 10, 10 -> 8
			// srcs: (6, 5)(269) 22, (12) 32 --> (869) 704:NW5, ND0, *, PEGB0
			9'd5 : rdata = 43'b0001101000101011000000000000000000010000000;
			// PEs: 10, 10 -> 8
			// srcs: (7, 6)(270) 32, (12) 32 --> (870) 1024:NW6, ND0, *, PEGB0
			9'd6 : rdata = 43'b0001101000110011000000000000000000010000000;
			// PEs: 10, 10 -> 8
			// srcs: (8, 7)(271) 29, (12) 32 --> (871) 928:NW7, ND0, *, PEGB0
			9'd7 : rdata = 43'b0001101000111011000000000000000000010000000;
			// PEs: 10, 10 -> 8
			// srcs: (9, 8)(272) 32, (12) 32 --> (872) 1024:NW8, ND0, *, PEGB0
			9'd8 : rdata = 43'b0001101001000011000000000000000000010000000;
			// PEs: 10, 10 -> 8
			// srcs: (10, 9)(273) 11, (12) 32 --> (873) 352:NW9, ND0, *, PEGB0
			9'd9 : rdata = 43'b0001101001001011000000000000000000010000000;
			// PEs: 10, 10 -> 8
			// srcs: (11, 10)(274) 49, (12) 32 --> (874) 1568:NW10, ND0, *, PEGB0
			9'd10 : rdata = 43'b0001101001010011000000000000000000010000000;
			// PEs: 10, 10 -> 8
			// srcs: (12, 11)(275) 48, (12) 32 --> (875) 1536:NW11, ND0, *, PEGB0
			9'd11 : rdata = 43'b0001101001011011000000000000000000010000000;
			// PEs: 10, 10 -> 8
			// srcs: (13, 12)(276) 22, (12) 32 --> (876) 704:NW12, ND0, *, PEGB0
			9'd12 : rdata = 43'b0001101001100011000000000000000000010000000;
			// PEs: 10, 10 -> 8
			// srcs: (14, 13)(277) 32, (12) 32 --> (877) 1024:NW13, ND0, *, PEGB0
			9'd13 : rdata = 43'b0001101001101011000000000000000000010000000;
			// PEs: 10, 10 -> 8
			// srcs: (15, 14)(278) 19, (12) 32 --> (878) 608:NW14, ND0, *, PEGB0
			9'd14 : rdata = 43'b0001101001110011000000000000000000010000000;
			// PEs: 10, 10 -> 8
			// srcs: (16, 15)(279) 4, (12) 32 --> (879) 128:NW15, ND0, *, PEGB0
			9'd15 : rdata = 43'b0001101001111011000000000000000000010000000;
			// PEs: 10, 10 -> 8
			// srcs: (17, 16)(280) 22, (12) 32 --> (880) 704:NW16, ND0, *, PEGB0
			9'd16 : rdata = 43'b0001101010000011000000000000000000010000000;
			// PEs: 10, 10 -> 8
			// srcs: (18, 17)(281) 7, (12) 32 --> (881) 224:NW17, ND0, *, PEGB0
			9'd17 : rdata = 43'b0001101010001011000000000000000000010000000;
			// PEs: 10, 10 -> 8
			// srcs: (19, 18)(282) 18, (12) 32 --> (882) 576:NW18, ND0, *, PEGB0
			9'd18 : rdata = 43'b0001101010010011000000000000000000010000000;
			// PEs: 10, 10 -> 8
			// srcs: (20, 19)(283) -3, (12) 32 --> (883) -96:NW19, ND0, *, PEGB0
			9'd19 : rdata = 43'b0001101010011011000000000000000000010000000;
			// PEs: 10, 10 -> 8
			// srcs: (21, 20)(284) 20, (12) 32 --> (884) 640:NW20, ND0, *, PEGB0
			9'd20 : rdata = 43'b0001101010100011000000000000000000010000000;
			// PEs: 10, 10 -> 8
			// srcs: (22, 21)(285) 4, (12) 32 --> (885) 128:NW21, ND0, *, PEGB0
			9'd21 : rdata = 43'b0001101010101011000000000000000000010000000;
			// PEs: 10, 10 -> 8
			// srcs: (23, 22)(286) 32, (12) 32 --> (886) 1024:NW22, ND0, *, PEGB0
			9'd22 : rdata = 43'b0001101010110011000000000000000000010000000;
			// PEs: 10, 10 -> 8
			// srcs: (24, 23)(287) 4, (12) 32 --> (887) 128:NW23, ND0, *, PEGB0
			9'd23 : rdata = 43'b0001101010111011000000000000000000010000000;
			// PEs: 10, 10 -> 9
			// srcs: (25, 24)(288) -1, (12) 32 --> (888) -32:NW24, ND0, *, PEGB1
			9'd24 : rdata = 43'b0001101011000011000000000000000000010010000;
			// PEs: 10, 10 -> 9
			// srcs: (26, 25)(289) 18, (12) 32 --> (889) 576:NW25, ND0, *, PEGB1
			9'd25 : rdata = 43'b0001101011001011000000000000000000010010000;
			// PEs: 10, 10 -> 12
			// srcs: (27, 26)(290) 40, (12) 32 --> (890) 1280:NW26, ND0, *, PEGB4
			9'd26 : rdata = 43'b0001101011010011000000000000000000011000000;
			// PEs: 10, 10 -> 9
			// srcs: (28, 27)(291) 17, (12) 32 --> (891) 544:NW27, ND0, *, PEGB1
			9'd27 : rdata = 43'b0001101011011011000000000000000000010010000;
			// PEs: 10, 10 -> 9
			// srcs: (29, 28)(292) 34, (12) 32 --> (892) 1088:NW28, ND0, *, PEGB1
			9'd28 : rdata = 43'b0001101011100011000000000000000000010010000;
			// PEs: 10, 10 -> 12
			// srcs: (30, 29)(293) 43, (12) 32 --> (893) 1376:NW29, ND0, *, PEGB4
			9'd29 : rdata = 43'b0001101011101011000000000000000000011000000;
			// PEs: 13 -> 10
			// srcs: (31, 38)(978) 1386 --> (978) 1386:PEGB5, pass, NI0
			9'd30 : rdata = 43'b1100011101010000000001000000000000000000000;
			// PEs: 13 -> 10
			// srcs: (32, 41)(979) 363 --> (979) 363:PEGB5, pass, NI1
			9'd31 : rdata = 43'b1100011101010000000001000010000000000000000;
			// PEs: 12, 10 -> 15
			// srcs: (33, 39)(948) 58, (978) 1386 --> (1685) 1444:PEGB4, NI0, +, PEGB7
			9'd32 : rdata = 43'b0000111101000101000000000000000000011110000;
			// PEs: 13 -> 10
			// srcs: (34, 44)(982) 726 --> (982) 726:PEGB5, pass, NI0
			9'd33 : rdata = 43'b1100011101010000000001000000000000000000000;
			// PEs: 12, 10 -> 11
			// srcs: (36, 42)(949) 696, (979) 363 --> (1704) 1059:PEGB4, NI1, +, PENB
			9'd34 : rdata = 43'b0000111101000101000010000000000000100000000;
			// PEs: 12, 10 -> 10
			// srcs: (39, 45)(952) 1363, (982) 726 --> (1761) 2089:PEGB4, NI0, +, NI1
			9'd35 : rdata = 43'b0000111101000101000001000010000000000000000;
			// PEs: 8 -> 
			// srcs: (145, 30)(673) 143 --> (673) 143:PEGB0, pass, 
			9'd36 : rdata = 43'b1100011100000000000000000000000000000000000;
			// PEs: 8, 10 -> 10
			// srcs: (154, 31)(643) 266, (673) 143 --> (1585) 409:PEGB0, ALU, +, NI0
			9'd37 : rdata = 43'b0000111100000001111111000000000000000000000;
			// PEs: 8 -> 
			// srcs: (156, 32)(733) 460 --> (733) 460:PEGB0, pass, 
			9'd38 : rdata = 43'b1100011100000000000000000000000000000000000;
			// PEs: 8, 10 -> 10
			// srcs: (165, 33)(703) 72, (733) 460 --> (1586) 532:PEGB0, ALU, +, NI2
			9'd39 : rdata = 43'b0000111100000001111111000100000000000000000;
			// PEs: 8 -> 10
			// srcs: (167, 34)(793) 95 --> (793) 95:PEGB0, pass, NI3
			9'd40 : rdata = 43'b1100011100000000000001000110000000000000000;
			// PEs: 10 -> 10
			// srcs: (168, 59)(1585) 409 --> (1585) 409:NI0, pass, NI0
			9'd41 : rdata = 43'b1100010100000000000001000000000000000000000;
			// PEs: 10, 10 -> 10
			// srcs: (168, 46)(1585) 409, (1586) 532 --> (1595) 941:ALU, NI2, +, NI4
			9'd42 : rdata = 43'b0000100111111101000101001000000000000000000;
			// PEs: 8, 10 -> 8
			// srcs: (176, 35)(763) -72, (793) 95 --> (1587) 23:PEGB0, NI3, +, PEGB0
			9'd43 : rdata = 43'b0000111100000101000110000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (209, 54)(1595) 941 --> (1595) 941:NI4, pass, PEGB0
			9'd44 : rdata = 43'b1100010100100000000000000000000000010000000;
			// PEs: 8, 9 -> 10
			// srcs: (218, 36)(825) 403, (855) -64 --> (1626) 339:PEGB0, PENB, +, NI0
			9'd45 : rdata = 43'b0000111100000110111101000000000000000000000;
			// PEs: 8, 9 -> 10
			// srcs: (242, 37)(826) 248, (856) 192 --> (1645) 440:PEGB0, PENB, +, NI2
			9'd46 : rdata = 43'b0000111100000110111101000100000000000000000;
			// PEs: 8, 9 -> 8
			// srcs: (274, 40)(829) 992, (859) 320 --> (1702) 1312:PEGB0, PENB, +, PEGB0
			9'd47 : rdata = 43'b0000111100000110111100000000000000010000000;
			// PEs: 8, 9 -> 9
			// srcs: (277, 43)(832) 341, (862) 1152 --> (1759) 1493:PEGB0, PENB, +, PEGB1
			9'd48 : rdata = 43'b0000111100000110111100000000000000010010000;
			// PEs: 9, 10 -> 10
			// srcs: (278, 47)(1625) 761, (1626) 339 --> (1634) 1100:PENB, NI0, +, NI3
			9'd49 : rdata = 43'b0000111011110101000001000110000000000000000;
			// PEs: 9, 10 -> 10
			// srcs: (279, 48)(1644) 960, (1645) 440 --> (1653) 1400:PENB, NI2, +, NI0
			9'd50 : rdata = 43'b0000111011110101000101000000000000000000000;
			// PEs: 9 -> 
			// srcs: (280, 49)(1664) 761 --> (1664) 761:PENB, pass, 
			9'd51 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 9, 10 -> 9
			// srcs: (286, 50)(1663) 1071, (1664) 761 --> (1672) 1832:PENB, ALU, +, PEGB1
			9'd52 : rdata = 43'b0000111011110001111110000000000000010010000;
			// PEs: 9, 10 -> 8
			// srcs: (287, 51)(1760) 1062, (1761) 2089 --> (1768) 3151:PENB, NI1, +, PEGB0
			9'd53 : rdata = 43'b0000111011110101000010000000000000010000000;
			// PEs: 9 -> 10
			// srcs: (288, 52)(1594) 847 --> (1594) 847:PENB, pass, NI1
			9'd54 : rdata = 43'b1100011011110000000001000010000000000000000;
			// PEs: 9, 10 -> 10
			// srcs: (289, 55)(1633) 1981, (1634) 1100 --> (1638) 3081:PENB, NI3, +, NI2
			9'd55 : rdata = 43'b0000111011110101000111000100000000000000000;
			// PEs: 9, 10 -> 10
			// srcs: (290, 56)(1652) 2643, (1653) 1400 --> (1657) 4043:PENB, NI0, +, NI3
			9'd56 : rdata = 43'b0000111011110101000001000110000000000000000;
			// PEs: 9, 10 -> 8
			// srcs: (405, 53)(1593) 1228, (1594) 847 --> (1599) 2075:PENB, NI1, +, PEGB0
			9'd57 : rdata = 43'b0000111011110101000010000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (529, 57)(1638) 3081 --> (1638) 3081:NI2, pass, PEGB0
			9'd58 : rdata = 43'b1100010100010000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (537, 58)(1657) 4043 --> (1657) 4043:NI3, pass, PEGB0
			9'd59 : rdata = 43'b1100010100011000000000000000000000010000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 11) begin
	always @(*) begin
		case(address)
			// PEs: 11, 11 -> 8
			// srcs: (1, 0)(294) 22, (13) -1 --> (894) -22:NW0, ND0, *, PEGB0
			9'd0 : rdata = 43'b0001101000000011000000000000000000010000000;
			// PEs: 11, 11 -> 8
			// srcs: (2, 1)(295) 23, (13) -1 --> (895) -23:NW1, ND0, *, PEGB0
			9'd1 : rdata = 43'b0001101000001011000000000000000000010000000;
			// PEs: 11, 11 -> 8
			// srcs: (3, 2)(296) 5, (13) -1 --> (896) -5:NW2, ND0, *, PEGB0
			9'd2 : rdata = 43'b0001101000010011000000000000000000010000000;
			// PEs: 11, 11 -> 8
			// srcs: (4, 3)(297) 9, (13) -1 --> (897) -9:NW3, ND0, *, PEGB0
			9'd3 : rdata = 43'b0001101000011011000000000000000000010000000;
			// PEs: 11, 11 -> 8
			// srcs: (5, 4)(298) 9, (13) -1 --> (898) -9:NW4, ND0, *, PEGB0
			9'd4 : rdata = 43'b0001101000100011000000000000000000010000000;
			// PEs: 11, 11 -> 8
			// srcs: (6, 5)(299) 4, (13) -1 --> (899) -4:NW5, ND0, *, PEGB0
			9'd5 : rdata = 43'b0001101000101011000000000000000000010000000;
			// PEs: 11, 11 -> 8
			// srcs: (7, 6)(300) -2, (13) -1 --> (900) 2:NW6, ND0, *, PEGB0
			9'd6 : rdata = 43'b0001101000110011000000000000000000010000000;
			// PEs: 11, 11 -> 8
			// srcs: (8, 7)(301) 47, (13) -1 --> (901) -47:NW7, ND0, *, PEGB0
			9'd7 : rdata = 43'b0001101000111011000000000000000000010000000;
			// PEs: 11, 11 -> 8
			// srcs: (9, 8)(302) 45, (13) -1 --> (902) -45:NW8, ND0, *, PEGB0
			9'd8 : rdata = 43'b0001101001000011000000000000000000010000000;
			// PEs: 11, 11 -> 8
			// srcs: (10, 9)(303) 37, (13) -1 --> (903) -37:NW9, ND0, *, PEGB0
			9'd9 : rdata = 43'b0001101001001011000000000000000000010000000;
			// PEs: 11, 11 -> 8
			// srcs: (11, 10)(304) 4, (13) -1 --> (904) -4:NW10, ND0, *, PEGB0
			9'd10 : rdata = 43'b0001101001010011000000000000000000010000000;
			// PEs: 11, 11 -> 8
			// srcs: (12, 11)(305) 35, (13) -1 --> (905) -35:NW11, ND0, *, PEGB0
			9'd11 : rdata = 43'b0001101001011011000000000000000000010000000;
			// PEs: 11, 11 -> 8
			// srcs: (13, 12)(306) 28, (13) -1 --> (906) -28:NW12, ND0, *, PEGB0
			9'd12 : rdata = 43'b0001101001100011000000000000000000010000000;
			// PEs: 11, 11 -> 8
			// srcs: (14, 13)(307) 13, (13) -1 --> (907) -13:NW13, ND0, *, PEGB0
			9'd13 : rdata = 43'b0001101001101011000000000000000000010000000;
			// PEs: 11, 11 -> 8
			// srcs: (15, 14)(308) 20, (13) -1 --> (908) -20:NW14, ND0, *, PEGB0
			9'd14 : rdata = 43'b0001101001110011000000000000000000010000000;
			// PEs: 11, 11 -> 8
			// srcs: (16, 15)(309) 37, (13) -1 --> (909) -37:NW15, ND0, *, PEGB0
			9'd15 : rdata = 43'b0001101001111011000000000000000000010000000;
			// PEs: 11, 11 -> 8
			// srcs: (17, 16)(310) 2, (13) -1 --> (910) -2:NW16, ND0, *, PEGB0
			9'd16 : rdata = 43'b0001101010000011000000000000000000010000000;
			// PEs: 11, 11 -> 8
			// srcs: (18, 17)(311) 14, (13) -1 --> (911) -14:NW17, ND0, *, PEGB0
			9'd17 : rdata = 43'b0001101010001011000000000000000000010000000;
			// PEs: 11, 11 -> 8
			// srcs: (19, 18)(312) 20, (13) -1 --> (912) -20:NW18, ND0, *, PEGB0
			9'd18 : rdata = 43'b0001101010010011000000000000000000010000000;
			// PEs: 11, 11 -> 8
			// srcs: (20, 19)(313) 30, (13) -1 --> (913) -30:NW19, ND0, *, PEGB0
			9'd19 : rdata = 43'b0001101010011011000000000000000000010000000;
			// PEs: 11, 11 -> 8
			// srcs: (21, 20)(314) 19, (13) -1 --> (914) -19:NW20, ND0, *, PEGB0
			9'd20 : rdata = 43'b0001101010100011000000000000000000010000000;
			// PEs: 11, 11 -> 8
			// srcs: (22, 21)(315) 2, (13) -1 --> (915) -2:NW21, ND0, *, PEGB0
			9'd21 : rdata = 43'b0001101010101011000000000000000000010000000;
			// PEs: 11, 11 -> 8
			// srcs: (23, 22)(316) 23, (13) -1 --> (916) -23:NW22, ND0, *, PEGB0
			9'd22 : rdata = 43'b0001101010110011000000000000000000010000000;
			// PEs: 11, 11 -> 8
			// srcs: (24, 23)(317) 39, (13) -1 --> (917) -39:NW23, ND0, *, PEGB0
			9'd23 : rdata = 43'b0001101010111011000000000000000000010000000;
			// PEs: 11, 11 -> 9
			// srcs: (25, 24)(318) 2, (13) -1 --> (918) -2:NW24, ND0, *, PEGB1
			9'd24 : rdata = 43'b0001101011000011000000000000000000010010000;
			// PEs: 11, 11 -> 9
			// srcs: (26, 25)(319) 21, (13) -1 --> (919) -21:NW25, ND0, *, PEGB1
			9'd25 : rdata = 43'b0001101011001011000000000000000000010010000;
			// PEs: 11, 11 -> 12
			// srcs: (27, 26)(320) 27, (13) -1 --> (920) -27:NW26, ND0, *, PENB
			9'd26 : rdata = 43'b0001101011010011000000000000000000100000000;
			// PEs: 11, 11 -> 9
			// srcs: (28, 27)(321) 10, (13) -1 --> (921) -10:NW27, ND0, *, PEGB1
			9'd27 : rdata = 43'b0001101011011011000000000000000000010010000;
			// PEs: 11, 11 -> 9
			// srcs: (29, 28)(322) 26, (13) -1 --> (922) -26:NW28, ND0, *, PEGB1
			9'd28 : rdata = 43'b0001101011100011000000000000000000010010000;
			// PEs: 11, 11 -> 12
			// srcs: (30, 29)(323) 6, (13) -1 --> (923) -6:NW29, ND0, *, PENB
			9'd29 : rdata = 43'b0001101011101011000000000000000000100000000;
			// PEs: 15 -> 11
			// srcs: (31, 30)(1038) 682 --> (1038) 682:PEGB7, pass, NI0
			9'd30 : rdata = 43'b1100011101110000000001000000000000000000000;
			// PEs: 15 -> 11
			// srcs: (32, 32)(1039) 330 --> (1039) 330:PEGB7, pass, NI1
			9'd31 : rdata = 43'b1100011101110000000001000010000000000000000;
			// PEs: 14, 11 -> 8
			// srcs: (33, 31)(1008) 42, (1038) 682 --> (1686) 724:PEGB6, NI0, +, PEGB0
			9'd32 : rdata = 43'b0000111101100101000000000000000000010000000;
			// PEs: 14, 11 -> 8
			// srcs: (36, 33)(1009) 28, (1039) 330 --> (1705) 358:PEGB6, NI1, +, PEGB0
			9'd33 : rdata = 43'b0000111101100101000010000000000000010000000;
			// PEs: 14 -> 
			// srcs: (38, 35)(1723) 1296 --> (1723) 1296:PEGB6, pass, 
			9'd34 : rdata = 43'b1100011101100000000000000000000000000000000;
			// PEs: 12, 11 -> 11
			// srcs: (41, 36)(1722) 1253, (1723) 1296 --> (1730) 2549:PEGB4, ALU, +, NI0
			9'd35 : rdata = 43'b0000111101000001111111000000000000000000000;
			// PEs: 9, 10 -> 8
			// srcs: (42, 34)(1703) 555, (1704) 1059 --> (1711) 1614:PEGB1, PENB, +, PEGB0
			9'd36 : rdata = 43'b0000111100010110111100000000000000010000000;
			// PEs: 11 -> 8
			// srcs: (517, 37)(1730) 2549 --> (1730) 2549:NI0, pass, PEGB0
			9'd37 : rdata = 43'b1100010100000000000000000000000000010000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 12) begin
	always @(*) begin
		case(address)
			// PEs: 12, 12 -> 8
			// srcs: (1, 0)(324) 23, (14) 29 --> (924) 667:NW0, ND0, *, PEGB0
			9'd0 : rdata = 43'b0001101000000011000000000000000000010000000;
			// PEs: 12, 12 -> 8
			// srcs: (2, 1)(325) 22, (14) 29 --> (925) 638:NW1, ND0, *, PEGB0
			9'd1 : rdata = 43'b0001101000001011000000000000000000010000000;
			// PEs: 12, 12 -> 8
			// srcs: (3, 2)(326) 4, (14) 29 --> (926) 116:NW2, ND0, *, PEGB0
			9'd2 : rdata = 43'b0001101000010011000000000000000000010000000;
			// PEs: 12, 12 -> 8
			// srcs: (4, 3)(327) 1, (14) 29 --> (927) 29:NW3, ND0, *, PEGB0
			9'd3 : rdata = 43'b0001101000011011000000000000000000010000000;
			// PEs: 12, 12 -> 8
			// srcs: (5, 4)(328) 1, (14) 29 --> (928) 29:NW4, ND0, *, PEGB0
			9'd4 : rdata = 43'b0001101000100011000000000000000000010000000;
			// PEs: 12, 12 -> 8
			// srcs: (6, 5)(329) 35, (14) 29 --> (929) 1015:NW5, ND0, *, PEGB0
			9'd5 : rdata = 43'b0001101000101011000000000000000000010000000;
			// PEs: 12, 12 -> 8
			// srcs: (7, 6)(330) 45, (14) 29 --> (930) 1305:NW6, ND0, *, PEGB0
			9'd6 : rdata = 43'b0001101000110011000000000000000000010000000;
			// PEs: 12, 12 -> 8
			// srcs: (8, 7)(331) 16, (14) 29 --> (931) 464:NW7, ND0, *, PEGB0
			9'd7 : rdata = 43'b0001101000111011000000000000000000010000000;
			// PEs: 12, 12 -> 8
			// srcs: (9, 8)(332) 20, (14) 29 --> (932) 580:NW8, ND0, *, PEGB0
			9'd8 : rdata = 43'b0001101001000011000000000000000000010000000;
			// PEs: 12, 12 -> 8
			// srcs: (10, 9)(333) 14, (14) 29 --> (933) 406:NW9, ND0, *, PEGB0
			9'd9 : rdata = 43'b0001101001001011000000000000000000010000000;
			// PEs: 12, 12 -> 8
			// srcs: (11, 10)(334) 39, (14) 29 --> (934) 1131:NW10, ND0, *, PEGB0
			9'd10 : rdata = 43'b0001101001010011000000000000000000010000000;
			// PEs: 12, 12 -> 8
			// srcs: (12, 11)(335) 36, (14) 29 --> (935) 1044:NW11, ND0, *, PEGB0
			9'd11 : rdata = 43'b0001101001011011000000000000000000010000000;
			// PEs: 12, 12 -> 8
			// srcs: (13, 12)(336) 10, (14) 29 --> (936) 290:NW12, ND0, *, PEGB0
			9'd12 : rdata = 43'b0001101001100011000000000000000000010000000;
			// PEs: 12, 12 -> 8
			// srcs: (14, 13)(337) 19, (14) 29 --> (937) 551:NW13, ND0, *, PEGB0
			9'd13 : rdata = 43'b0001101001101011000000000000000000010000000;
			// PEs: 12, 12 -> 8
			// srcs: (15, 14)(338) -3, (14) 29 --> (938) -87:NW14, ND0, *, PEGB0
			9'd14 : rdata = 43'b0001101001110011000000000000000000010000000;
			// PEs: 12, 12 -> 8
			// srcs: (16, 15)(339) 27, (14) 29 --> (939) 783:NW15, ND0, *, PEGB0
			9'd15 : rdata = 43'b0001101001111011000000000000000000010000000;
			// PEs: 12, 12 -> 8
			// srcs: (17, 16)(340) 12, (14) 29 --> (940) 348:NW16, ND0, *, PEGB0
			9'd16 : rdata = 43'b0001101010000011000000000000000000010000000;
			// PEs: 12, 12 -> 8
			// srcs: (18, 17)(341) 46, (14) 29 --> (941) 1334:NW17, ND0, *, PEGB0
			9'd17 : rdata = 43'b0001101010001011000000000000000000010000000;
			// PEs: 12, 12 -> 8
			// srcs: (19, 18)(342) 44, (14) 29 --> (942) 1276:NW18, ND0, *, PEGB0
			9'd18 : rdata = 43'b0001101010010011000000000000000000010000000;
			// PEs: 12, 12 -> 8
			// srcs: (20, 19)(343) 7, (14) 29 --> (943) 203:NW19, ND0, *, PEGB0
			9'd19 : rdata = 43'b0001101010011011000000000000000000010000000;
			// PEs: 12, 12 -> 8
			// srcs: (21, 20)(344) 20, (14) 29 --> (944) 580:NW20, ND0, *, PEGB0
			9'd20 : rdata = 43'b0001101010100011000000000000000000010000000;
			// PEs: 12, 12 -> 8
			// srcs: (22, 21)(345) 3, (14) 29 --> (945) 87:NW21, ND0, *, PEGB0
			9'd21 : rdata = 43'b0001101010101011000000000000000000010000000;
			// PEs: 12, 12 -> 8
			// srcs: (23, 22)(346) 49, (14) 29 --> (946) 1421:NW22, ND0, *, PEGB0
			9'd22 : rdata = 43'b0001101010110011000000000000000000010000000;
			// PEs: 12, 12 -> 8
			// srcs: (24, 23)(347) 35, (14) 29 --> (947) 1015:NW23, ND0, *, PEGB0
			9'd23 : rdata = 43'b0001101010111011000000000000000000010000000;
			// PEs: 12, 12 -> 10
			// srcs: (25, 24)(348) 2, (14) 29 --> (948) 58:NW24, ND0, *, PEGB2
			9'd24 : rdata = 43'b0001101011000011000000000000000000010100000;
			// PEs: 12, 12 -> 10
			// srcs: (26, 25)(349) 24, (14) 29 --> (949) 696:NW25, ND0, *, PEGB2
			9'd25 : rdata = 43'b0001101011001011000000000000000000010100000;
			// PEs: 12, 12 -> 14
			// srcs: (27, 26)(350) 6, (14) 29 --> (950) 174:NW26, ND0, *, PEGB6
			9'd26 : rdata = 43'b0001101011010011000000000000000000011100000;
			// PEs: 12, 12 -> 13
			// srcs: (28, 27)(351) 49, (14) 29 --> (951) 1421:NW27, ND0, *, PENB
			9'd27 : rdata = 43'b0001101011011011000000000000000000100000000;
			// PEs: 12, 12 -> 10
			// srcs: (29, 28)(352) 47, (14) 29 --> (952) 1363:NW28, ND0, *, PEGB2
			9'd28 : rdata = 43'b0001101011100011000000000000000000010100000;
			// PEs: 12, 12 -> 13
			// srcs: (30, 29)(353) 6, (14) 29 --> (953) 174:NW29, ND0, *, PENB
			9'd29 : rdata = 43'b0001101011101011000000000000000000100000000;
			// PEs: 10, 11 -> 11
			// srcs: (33, 32)(890) 1280, (920) -27 --> (1722) 1253:PEGB2, PENB, +, PEGB3
			9'd30 : rdata = 43'b0000111100100110111100000000000000010110000;
			// PEs: 10, 11 -> 13
			// srcs: (36, 33)(893) 1376, (923) -6 --> (1779) 1370:PEGB2, PENB, +, PENB
			9'd31 : rdata = 43'b0000111100100110111100000000000000100000000;
			// PEs: 8 -> 
			// srcs: (194, 30)(824) 713 --> (824) 713:PEGB0, pass, 
			9'd32 : rdata = 43'b1100011100000000000000000000000000000000000;
			// PEs: 12, 9 -> 9
			// srcs: (196, 31)(824) 713, (854) 1344 --> (1607) 2057:ALU, PEGB1, +, PEGB1
			9'd33 : rdata = 43'b0000100111111111000100000000000000010010000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 13) begin
	always @(*) begin
		case(address)
			// PEs: 13, 13 -> 8
			// srcs: (1, 0)(354) 47, (15) 33 --> (954) 1551:NW0, ND0, *, PEGB0
			9'd0 : rdata = 43'b0001101000000011000000000000000000010000000;
			// PEs: 13, 13 -> 8
			// srcs: (2, 1)(355) 14, (15) 33 --> (955) 462:NW1, ND0, *, PEGB0
			9'd1 : rdata = 43'b0001101000001011000000000000000000010000000;
			// PEs: 13, 13 -> 8
			// srcs: (3, 2)(356) 5, (15) 33 --> (956) 165:NW2, ND0, *, PEGB0
			9'd2 : rdata = 43'b0001101000010011000000000000000000010000000;
			// PEs: 13, 13 -> 8
			// srcs: (4, 3)(357) 40, (15) 33 --> (957) 1320:NW3, ND0, *, PEGB0
			9'd3 : rdata = 43'b0001101000011011000000000000000000010000000;
			// PEs: 13, 13 -> 8
			// srcs: (5, 4)(358) 23, (15) 33 --> (958) 759:NW4, ND0, *, PEGB0
			9'd4 : rdata = 43'b0001101000100011000000000000000000010000000;
			// PEs: 13, 13 -> 8
			// srcs: (6, 5)(359) 30, (15) 33 --> (959) 990:NW5, ND0, *, PEGB0
			9'd5 : rdata = 43'b0001101000101011000000000000000000010000000;
			// PEs: 13, 13 -> 8
			// srcs: (7, 6)(360) -1, (15) 33 --> (960) -33:NW6, ND0, *, PEGB0
			9'd6 : rdata = 43'b0001101000110011000000000000000000010000000;
			// PEs: 13, 13 -> 8
			// srcs: (8, 7)(361) 11, (15) 33 --> (961) 363:NW7, ND0, *, PEGB0
			9'd7 : rdata = 43'b0001101000111011000000000000000000010000000;
			// PEs: 13, 13 -> 8
			// srcs: (9, 8)(362) 3, (15) 33 --> (962) 99:NW8, ND0, *, PEGB0
			9'd8 : rdata = 43'b0001101001000011000000000000000000010000000;
			// PEs: 13, 13 -> 8
			// srcs: (10, 9)(363) 1, (15) 33 --> (963) 33:NW9, ND0, *, PEGB0
			9'd9 : rdata = 43'b0001101001001011000000000000000000010000000;
			// PEs: 13, 13 -> 8
			// srcs: (11, 10)(364) 22, (15) 33 --> (964) 726:NW10, ND0, *, PEGB0
			9'd10 : rdata = 43'b0001101001010011000000000000000000010000000;
			// PEs: 13, 13 -> 8
			// srcs: (12, 11)(365) -3, (15) 33 --> (965) -99:NW11, ND0, *, PEGB0
			9'd11 : rdata = 43'b0001101001011011000000000000000000010000000;
			// PEs: 13, 13 -> 8
			// srcs: (13, 12)(366) 46, (15) 33 --> (966) 1518:NW12, ND0, *, PEGB0
			9'd12 : rdata = 43'b0001101001100011000000000000000000010000000;
			// PEs: 13, 13 -> 8
			// srcs: (14, 13)(367) 45, (15) 33 --> (967) 1485:NW13, ND0, *, PEGB0
			9'd13 : rdata = 43'b0001101001101011000000000000000000010000000;
			// PEs: 13, 13 -> 8
			// srcs: (15, 14)(368) 7, (15) 33 --> (968) 231:NW14, ND0, *, PEGB0
			9'd14 : rdata = 43'b0001101001110011000000000000000000010000000;
			// PEs: 13, 13 -> 8
			// srcs: (16, 15)(369) 26, (15) 33 --> (969) 858:NW15, ND0, *, PEGB0
			9'd15 : rdata = 43'b0001101001111011000000000000000000010000000;
			// PEs: 13, 13 -> 8
			// srcs: (17, 16)(370) 27, (15) 33 --> (970) 891:NW16, ND0, *, PEGB0
			9'd16 : rdata = 43'b0001101010000011000000000000000000010000000;
			// PEs: 13, 13 -> 8
			// srcs: (18, 17)(371) 48, (15) 33 --> (971) 1584:NW17, ND0, *, PEGB0
			9'd17 : rdata = 43'b0001101010001011000000000000000000010000000;
			// PEs: 13, 13 -> 8
			// srcs: (19, 18)(372) 17, (15) 33 --> (972) 561:NW18, ND0, *, PEGB0
			9'd18 : rdata = 43'b0001101010010011000000000000000000010000000;
			// PEs: 13, 13 -> 8
			// srcs: (20, 19)(373) 11, (15) 33 --> (973) 363:NW19, ND0, *, PEGB0
			9'd19 : rdata = 43'b0001101010011011000000000000000000010000000;
			// PEs: 13, 13 -> 8
			// srcs: (21, 20)(374) 23, (15) 33 --> (974) 759:NW20, ND0, *, PEGB0
			9'd20 : rdata = 43'b0001101010100011000000000000000000010000000;
			// PEs: 13, 13 -> 8
			// srcs: (22, 21)(375) 33, (15) 33 --> (975) 1089:NW21, ND0, *, PEGB0
			9'd21 : rdata = 43'b0001101010101011000000000000000000010000000;
			// PEs: 13, 13 -> 8
			// srcs: (23, 22)(376) 27, (15) 33 --> (976) 891:NW22, ND0, *, PEGB0
			9'd22 : rdata = 43'b0001101010110011000000000000000000010000000;
			// PEs: 13, 13 -> 8
			// srcs: (24, 23)(377) 4, (15) 33 --> (977) 132:NW23, ND0, *, PEGB0
			9'd23 : rdata = 43'b0001101010111011000000000000000000010000000;
			// PEs: 13, 13 -> 10
			// srcs: (25, 24)(378) 42, (15) 33 --> (978) 1386:NW24, ND0, *, PEGB2
			9'd24 : rdata = 43'b0001101011000011000000000000000000010100000;
			// PEs: 13, 13 -> 10
			// srcs: (26, 25)(379) 11, (15) 33 --> (979) 363:NW25, ND0, *, PEGB2
			9'd25 : rdata = 43'b0001101011001011000000000000000000010100000;
			// PEs: 13, 13 -> 14
			// srcs: (27, 26)(380) 34, (15) 33 --> (980) 1122:NW26, ND0, *, PENB
			9'd26 : rdata = 43'b0001101011010011000000000000000000100000000;
			// PEs: 13, 13 -> 13
			// srcs: (28, 27)(381) 1, (15) 33 --> (981) 33:NW27, ND0, *, NI0
			9'd27 : rdata = 43'b0001101011011011000001000000000000000000000;
			// PEs: 13, 13 -> 10
			// srcs: (29, 28)(382) 22, (15) 33 --> (982) 726:NW28, ND0, *, PEGB2
			9'd28 : rdata = 43'b0001101011100011000000000000000000010100000;
			// PEs: 13, 13 -> 13
			// srcs: (30, 29)(383) 23, (15) 33 --> (983) 759:NW29, ND0, *, NI1
			9'd29 : rdata = 43'b0001101011101011000001000010000000000000000;
			// PEs: 12, 13 -> 9
			// srcs: (31, 32)(951) 1421, (981) 33 --> (1742) 1454:PENB, NI0, +, PEGB1
			9'd30 : rdata = 43'b0000111011110101000000000000000000010010000;
			// PEs: 15 -> 13
			// srcs: (32, 30)(1040) 440 --> (1040) 440:PEGB7, pass, NI0
			9'd31 : rdata = 43'b1100011101110000000001000000000000000000000;
			// PEs: 12, 13 -> 13
			// srcs: (33, 33)(953) 174, (983) 759 --> (1780) 933:PENB, NI1, +, NI2
			9'd32 : rdata = 43'b0000111011110101000011000100000000000000000;
			// PEs: 14, 13 -> 8
			// srcs: (35, 31)(1010) 42, (1040) 440 --> (1724) 482:PEGB6, NI0, +, PEGB0
			9'd33 : rdata = 43'b0000111101100101000000000000000000010000000;
			// PEs: 12, 13 -> 8
			// srcs: (39, 34)(1779) 1370, (1780) 933 --> (1787) 2303:PENB, NI2, +, PEGB0
			9'd34 : rdata = 43'b0000111011110101000100000000000000010000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 14) begin
	always @(*) begin
		case(address)
			// PEs: 14, 14 -> 8
			// srcs: (1, 0)(384) 46, (16) 2 --> (984) 92:NW0, ND0, *, PEGB0
			9'd0 : rdata = 43'b0001101000000011000000000000000000010000000;
			// PEs: 14, 14 -> 8
			// srcs: (2, 1)(385) 26, (16) 2 --> (985) 52:NW1, ND0, *, PEGB0
			9'd1 : rdata = 43'b0001101000001011000000000000000000010000000;
			// PEs: 14, 14 -> 8
			// srcs: (3, 2)(386) 28, (16) 2 --> (986) 56:NW2, ND0, *, PEGB0
			9'd2 : rdata = 43'b0001101000010011000000000000000000010000000;
			// PEs: 14, 14 -> 8
			// srcs: (4, 3)(387) 47, (16) 2 --> (987) 94:NW3, ND0, *, PEGB0
			9'd3 : rdata = 43'b0001101000011011000000000000000000010000000;
			// PEs: 14, 14 -> 8
			// srcs: (5, 4)(388) 9, (16) 2 --> (988) 18:NW4, ND0, *, PEGB0
			9'd4 : rdata = 43'b0001101000100011000000000000000000010000000;
			// PEs: 14, 14 -> 8
			// srcs: (6, 5)(389) 45, (16) 2 --> (989) 90:NW5, ND0, *, PEGB0
			9'd5 : rdata = 43'b0001101000101011000000000000000000010000000;
			// PEs: 14, 14 -> 8
			// srcs: (7, 6)(390) 41, (16) 2 --> (990) 82:NW6, ND0, *, PEGB0
			9'd6 : rdata = 43'b0001101000110011000000000000000000010000000;
			// PEs: 14, 14 -> 8
			// srcs: (8, 7)(391) 25, (16) 2 --> (991) 50:NW7, ND0, *, PEGB0
			9'd7 : rdata = 43'b0001101000111011000000000000000000010000000;
			// PEs: 14, 14 -> 8
			// srcs: (9, 8)(392) 25, (16) 2 --> (992) 50:NW8, ND0, *, PEGB0
			9'd8 : rdata = 43'b0001101001000011000000000000000000010000000;
			// PEs: 14, 14 -> 8
			// srcs: (10, 9)(393) 37, (16) 2 --> (993) 74:NW9, ND0, *, PEGB0
			9'd9 : rdata = 43'b0001101001001011000000000000000000010000000;
			// PEs: 14, 14 -> 8
			// srcs: (11, 10)(394) 11, (16) 2 --> (994) 22:NW10, ND0, *, PEGB0
			9'd10 : rdata = 43'b0001101001010011000000000000000000010000000;
			// PEs: 14, 14 -> 8
			// srcs: (12, 11)(395) 30, (16) 2 --> (995) 60:NW11, ND0, *, PEGB0
			9'd11 : rdata = 43'b0001101001011011000000000000000000010000000;
			// PEs: 14, 14 -> 8
			// srcs: (13, 12)(396) 32, (16) 2 --> (996) 64:NW12, ND0, *, PEGB0
			9'd12 : rdata = 43'b0001101001100011000000000000000000010000000;
			// PEs: 14, 14 -> 8
			// srcs: (14, 13)(397) 39, (16) 2 --> (997) 78:NW13, ND0, *, PEGB0
			9'd13 : rdata = 43'b0001101001101011000000000000000000010000000;
			// PEs: 14, 14 -> 8
			// srcs: (15, 14)(398) 0, (16) 2 --> (998) 0:NW14, ND0, *, PEGB0
			9'd14 : rdata = 43'b0001101001110011000000000000000000010000000;
			// PEs: 14, 14 -> 8
			// srcs: (16, 15)(399) 22, (16) 2 --> (999) 44:NW15, ND0, *, PEGB0
			9'd15 : rdata = 43'b0001101001111011000000000000000000010000000;
			// PEs: 14, 14 -> 8
			// srcs: (17, 16)(400) 26, (16) 2 --> (1000) 52:NW16, ND0, *, PEGB0
			9'd16 : rdata = 43'b0001101010000011000000000000000000010000000;
			// PEs: 14, 14 -> 8
			// srcs: (18, 17)(401) 15, (16) 2 --> (1001) 30:NW17, ND0, *, PEGB0
			9'd17 : rdata = 43'b0001101010001011000000000000000000010000000;
			// PEs: 14, 14 -> 8
			// srcs: (19, 18)(402) 21, (16) 2 --> (1002) 42:NW18, ND0, *, PEGB0
			9'd18 : rdata = 43'b0001101010010011000000000000000000010000000;
			// PEs: 14, 14 -> 8
			// srcs: (20, 19)(403) 47, (16) 2 --> (1003) 94:NW19, ND0, *, PEGB0
			9'd19 : rdata = 43'b0001101010011011000000000000000000010000000;
			// PEs: 14, 14 -> 8
			// srcs: (21, 20)(404) 16, (16) 2 --> (1004) 32:NW20, ND0, *, PEGB0
			9'd20 : rdata = 43'b0001101010100011000000000000000000010000000;
			// PEs: 14, 14 -> 8
			// srcs: (22, 21)(405) 22, (16) 2 --> (1005) 44:NW21, ND0, *, PEGB0
			9'd21 : rdata = 43'b0001101010101011000000000000000000010000000;
			// PEs: 14, 14 -> 8
			// srcs: (23, 22)(406) 35, (16) 2 --> (1006) 70:NW22, ND0, *, PEGB0
			9'd22 : rdata = 43'b0001101010110011000000000000000000010000000;
			// PEs: 14, 14 -> 8
			// srcs: (24, 23)(407) 36, (16) 2 --> (1007) 72:NW23, ND0, *, PEGB0
			9'd23 : rdata = 43'b0001101010111011000000000000000000010000000;
			// PEs: 14, 14 -> 11
			// srcs: (25, 24)(408) 21, (16) 2 --> (1008) 42:NW24, ND0, *, PEGB3
			9'd24 : rdata = 43'b0001101011000011000000000000000000010110000;
			// PEs: 14, 14 -> 11
			// srcs: (26, 25)(409) 14, (16) 2 --> (1009) 28:NW25, ND0, *, PEGB3
			9'd25 : rdata = 43'b0001101011001011000000000000000000010110000;
			// PEs: 14, 14 -> 13
			// srcs: (27, 26)(410) 21, (16) 2 --> (1010) 42:NW26, ND0, *, PEGB5
			9'd26 : rdata = 43'b0001101011010011000000000000000000011010000;
			// PEs: 14, 14 -> 15
			// srcs: (28, 27)(411) 49, (16) 2 --> (1011) 98:NW27, ND0, *, PENB
			9'd27 : rdata = 43'b0001101011011011000000000000000000100000000;
			// PEs: 14, 14 -> 15
			// srcs: (29, 28)(412) 7, (16) 2 --> (1012) 14:NW28, ND0, *, PENB
			9'd28 : rdata = 43'b0001101011100011000000000000000000100000000;
			// PEs: 14, 14 -> 15
			// srcs: (30, 29)(413) 37, (16) 2 --> (1013) 74:NW29, ND0, *, PENB
			9'd29 : rdata = 43'b0001101011101011000000000000000000100000000;
			// PEs: 12, 13 -> 11
			// srcs: (33, 30)(950) 174, (980) 1122 --> (1723) 1296:PEGB4, PENB, +, PEGB3
			9'd30 : rdata = 43'b0000111101000110111100000000000000010110000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 15) begin
	always @(*) begin
		case(address)
			// PEs: 15, 15 -> 8
			// srcs: (1, 0)(414) 21, (17) 22 --> (1014) 462:NW0, ND0, *, PENB
			9'd0 : rdata = 43'b0001101000000011000000000000000000100000000;
			// PEs: 15, 15 -> 8
			// srcs: (2, 1)(415) 2, (17) 22 --> (1015) 44:NW1, ND0, *, PENB
			9'd1 : rdata = 43'b0001101000001011000000000000000000100000000;
			// PEs: 15, 15 -> 8
			// srcs: (3, 2)(416) -1, (17) 22 --> (1016) -22:NW2, ND0, *, PENB
			9'd2 : rdata = 43'b0001101000010011000000000000000000100000000;
			// PEs: 15, 15 -> 8
			// srcs: (4, 3)(417) 44, (17) 22 --> (1017) 968:NW3, ND0, *, PENB
			9'd3 : rdata = 43'b0001101000011011000000000000000000100000000;
			// PEs: 15, 15 -> 8
			// srcs: (5, 4)(418) 20, (17) 22 --> (1018) 440:NW4, ND0, *, PENB
			9'd4 : rdata = 43'b0001101000100011000000000000000000100000000;
			// PEs: 15, 15 -> 8
			// srcs: (6, 5)(419) 23, (17) 22 --> (1019) 506:NW5, ND0, *, PENB
			9'd5 : rdata = 43'b0001101000101011000000000000000000100000000;
			// PEs: 15, 15 -> 8
			// srcs: (7, 6)(420) -1, (17) 22 --> (1020) -22:NW6, ND0, *, PENB
			9'd6 : rdata = 43'b0001101000110011000000000000000000100000000;
			// PEs: 15, 15 -> 8
			// srcs: (8, 7)(421) 40, (17) 22 --> (1021) 880:NW7, ND0, *, PENB
			9'd7 : rdata = 43'b0001101000111011000000000000000000100000000;
			// PEs: 15, 15 -> 8
			// srcs: (9, 8)(422) 3, (17) 22 --> (1022) 66:NW8, ND0, *, PENB
			9'd8 : rdata = 43'b0001101001000011000000000000000000100000000;
			// PEs: 15, 15 -> 8
			// srcs: (10, 9)(423) 28, (17) 22 --> (1023) 616:NW9, ND0, *, PENB
			9'd9 : rdata = 43'b0001101001001011000000000000000000100000000;
			// PEs: 15, 15 -> 8
			// srcs: (11, 10)(424) 38, (17) 22 --> (1024) 836:NW10, ND0, *, PENB
			9'd10 : rdata = 43'b0001101001010011000000000000000000100000000;
			// PEs: 15, 15 -> 8
			// srcs: (12, 11)(425) 14, (17) 22 --> (1025) 308:NW11, ND0, *, PENB
			9'd11 : rdata = 43'b0001101001011011000000000000000000100000000;
			// PEs: 15, 15 -> 8
			// srcs: (13, 12)(426) -1, (17) 22 --> (1026) -22:NW12, ND0, *, PENB
			9'd12 : rdata = 43'b0001101001100011000000000000000000100000000;
			// PEs: 15, 15 -> 8
			// srcs: (14, 13)(427) 36, (17) 22 --> (1027) 792:NW13, ND0, *, PENB
			9'd13 : rdata = 43'b0001101001101011000000000000000000100000000;
			// PEs: 15, 15 -> 8
			// srcs: (15, 14)(428) 45, (17) 22 --> (1028) 990:NW14, ND0, *, PENB
			9'd14 : rdata = 43'b0001101001110011000000000000000000100000000;
			// PEs: 15, 15 -> 8
			// srcs: (16, 15)(429) -1, (17) 22 --> (1029) -22:NW15, ND0, *, PENB
			9'd15 : rdata = 43'b0001101001111011000000000000000000100000000;
			// PEs: 15, 15 -> 8
			// srcs: (17, 16)(430) 21, (17) 22 --> (1030) 462:NW16, ND0, *, PENB
			9'd16 : rdata = 43'b0001101010000011000000000000000000100000000;
			// PEs: 15, 15 -> 8
			// srcs: (18, 17)(431) -2, (17) 22 --> (1031) -44:NW17, ND0, *, PENB
			9'd17 : rdata = 43'b0001101010001011000000000000000000100000000;
			// PEs: 15, 15 -> 8
			// srcs: (19, 18)(432) 27, (17) 22 --> (1032) 594:NW18, ND0, *, PENB
			9'd18 : rdata = 43'b0001101010010011000000000000000000100000000;
			// PEs: 15, 15 -> 8
			// srcs: (20, 19)(433) 29, (17) 22 --> (1033) 638:NW19, ND0, *, PENB
			9'd19 : rdata = 43'b0001101010011011000000000000000000100000000;
			// PEs: 15, 15 -> 8
			// srcs: (21, 20)(434) 10, (17) 22 --> (1034) 220:NW20, ND0, *, PENB
			9'd20 : rdata = 43'b0001101010100011000000000000000000100000000;
			// PEs: 15, 15 -> 8
			// srcs: (22, 21)(435) 15, (17) 22 --> (1035) 330:NW21, ND0, *, PENB
			9'd21 : rdata = 43'b0001101010101011000000000000000000100000000;
			// PEs: 15, 15 -> 8
			// srcs: (23, 22)(436) 0, (17) 22 --> (1036) 0:NW22, ND0, *, PENB
			9'd22 : rdata = 43'b0001101010110011000000000000000000100000000;
			// PEs: 15, 15 -> 8
			// srcs: (24, 23)(437) 10, (17) 22 --> (1037) 220:NW23, ND0, *, PENB
			9'd23 : rdata = 43'b0001101010111011000000000000000000100000000;
			// PEs: 15, 15 -> 11
			// srcs: (25, 24)(438) 31, (17) 22 --> (1038) 682:NW24, ND0, *, PEGB3
			9'd24 : rdata = 43'b0001101011000011000000000000000000010110000;
			// PEs: 15, 15 -> 11
			// srcs: (26, 25)(439) 15, (17) 22 --> (1039) 330:NW25, ND0, *, PEGB3
			9'd25 : rdata = 43'b0001101011001011000000000000000000010110000;
			// PEs: 15, 15 -> 13
			// srcs: (27, 26)(440) 20, (17) 22 --> (1040) 440:NW26, ND0, *, PEGB5
			9'd26 : rdata = 43'b0001101011010011000000000000000000011010000;
			// PEs: 15, 15 -> 15
			// srcs: (28, 27)(441) 21, (17) 22 --> (1041) 462:NW27, ND0, *, NI0
			9'd27 : rdata = 43'b0001101011011011000001000000000000000000000;
			// PEs: 15, 15 -> 15
			// srcs: (29, 28)(442) 4, (17) 22 --> (1042) 88:NW28, ND0, *, NI1
			9'd28 : rdata = 43'b0001101011100011000001000010000000000000000;
			// PEs: 15, 15 -> 15
			// srcs: (30, 29)(443) 21, (17) 22 --> (1043) 462:NW29, ND0, *, NI2
			9'd29 : rdata = 43'b0001101011101011000001000100000000000000000;
			// PEs: 14, 15 -> 8
			// srcs: (31, 30)(1011) 98, (1041) 462 --> (1743) 560:PENB, NI0, +, PENB
			9'd30 : rdata = 43'b0000111011110101000000000000000000100000000;
			// PEs: 14, 15 -> 8
			// srcs: (32, 31)(1012) 14, (1042) 88 --> (1762) 102:PENB, NI1, +, PENB
			9'd31 : rdata = 43'b0000111011110101000010000000000000100000000;
			// PEs: 14, 15 -> 8
			// srcs: (33, 32)(1013) 74, (1043) 462 --> (1781) 536:PENB, NI2, +, PENB
			9'd32 : rdata = 43'b0000111011110101000100000000000000100000000;
			// PEs: 10 -> 
			// srcs: (38, 33)(1685) 1444 --> (1685) 1444:PEGB2, pass, 
			9'd33 : rdata = 43'b1100011100100000000000000000000000000000000;
			// PEs: 9, 15 -> 8
			// srcs: (41, 34)(1684) -34, (1685) 1444 --> (1692) 1410:PEGB1, ALU, +, PENB
			9'd34 : rdata = 43'b0000111100010001111110000000000000100000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 16) begin
	always @(*) begin
		case(address)
			// PEs: 21 -> 24
			// srcs: (6, 3)(1164) -9 --> (1164) -9:PEGB5, pass, PUNB
			9'd0 : rdata = 43'b1100011101010000000000000000000001000000000;
			// PEs: 22 -> 24
			// srcs: (7, 4)(1194) 341 --> (1194) 341:PEGB6, pass, PUNB
			9'd1 : rdata = 43'b1100011101100000000000000000000001000000000;
			// PEs: 0 -> 16
			// srcs: (8, 0)(804) 1395 --> (804) 1395:PUGB0, pass, NI0
			9'd2 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 8 -> 23
			// srcs: (9, 1)(834) 992 --> (834) 992:PUNB, pass, PEGB7
			9'd3 : rdata = 43'b1100011011111000000000000000000000011110000;
			// PEs: 19 -> 24
			// srcs: (10, 17)(1105) 897 --> (1105) 897:PEGB3, pass, PUNB
			9'd4 : rdata = 43'b1100011100110000000000000000000001000000000;
			// PEs: 20 -> 24
			// srcs: (11, 18)(1135) -39 --> (1135) -39:PEGB4, pass, PUNB
			9'd5 : rdata = 43'b1100011101000000000000000000000001000000000;
			// PEs: 21 -> 24
			// srcs: (12, 19)(1165) 117 --> (1165) 117:PEGB5, pass, PUNB
			9'd6 : rdata = 43'b1100011101010000000000000000000001000000000;
			// PEs: 22 -> 24
			// srcs: (13, 20)(1195) 93 --> (1195) 93:PEGB6, pass, PUNB
			9'd7 : rdata = 43'b1100011101100000000000000000000001000000000;
			// PEs: 17 -> 24
			// srcs: (14, 21)(1046) 1152 --> (1046) 1152:PEGB1, pass, PUNB
			9'd8 : rdata = 43'b1100011100010000000000000000000001000000000;
			// PEs: 18 -> 24
			// srcs: (15, 22)(1076) 273 --> (1076) 273:PEGB2, pass, PUNB
			9'd9 : rdata = 43'b1100011100100000000000000000000001000000000;
			// PEs: 19 -> 24
			// srcs: (16, 23)(1106) 437 --> (1106) 437:PEGB3, pass, PUNB
			9'd10 : rdata = 43'b1100011100110000000000000000000001000000000;
			// PEs: 20 -> 24
			// srcs: (17, 24)(1136) 468 --> (1136) 468:PEGB4, pass, PUNB
			9'd11 : rdata = 43'b1100011101000000000000000000000001000000000;
			// PEs: 16 -> 23
			// srcs: (18, 2)(804) 1395 --> (804) 1395:NI0, pass, PEGB7
			9'd12 : rdata = 43'b1100010100000000000000000000000000011110000;
			// PEs: 0 -> 16
			// srcs: (19, 5)(805) 930 --> (805) 930:PUGB0, pass, NI0
			9'd13 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 8 -> 23
			// srcs: (20, 6)(835) 32 --> (835) 32:PUNB, pass, PEGB7
			9'd14 : rdata = 43'b1100011011111000000000000000000000011110000;
			// PEs: 21 -> 24
			// srcs: (21, 25)(1166) 162 --> (1166) 162:PEGB5, pass, PUNB
			9'd15 : rdata = 43'b1100011101010000000000000000000001000000000;
			// PEs: 22 -> 24
			// srcs: (22, 26)(1196) 1240 --> (1196) 1240:PEGB6, pass, PUNB
			9'd16 : rdata = 43'b1100011101100000000000000000000001000000000;
			// PEs: 17 -> 40
			// srcs: (23, 27)(1047) 1044 --> (1047) 1044:PEGB1, pass, PUGB5
			9'd17 : rdata = 43'b1100011100010000000000000000000000000001101;
			// PEs: 18 -> 40
			// srcs: (24, 28)(1077) 882 --> (1077) 882:PEGB2, pass, PUGB5
			9'd18 : rdata = 43'b1100011100100000000000000000000000000001101;
			// PEs: 19 -> 40
			// srcs: (25, 29)(1107) 805 --> (1107) 805:PEGB3, pass, PUGB5
			9'd19 : rdata = 43'b1100011100110000000000000000000000000001101;
			// PEs: 20 -> 40
			// srcs: (26, 30)(1137) 598 --> (1137) 598:PEGB4, pass, PUGB5
			9'd20 : rdata = 43'b1100011101000000000000000000000000000001101;
			// PEs: 21 -> 40
			// srcs: (27, 31)(1167) 162 --> (1167) 162:PEGB5, pass, PUGB5
			9'd21 : rdata = 43'b1100011101010000000000000000000000000001101;
			// PEs: 22 -> 40
			// srcs: (28, 32)(1197) 992 --> (1197) 992:PEGB6, pass, PUGB5
			9'd22 : rdata = 43'b1100011101100000000000000000000000000001101;
			// PEs: 16 -> 23
			// srcs: (29, 7)(805) 930 --> (805) 930:NI0, pass, PEGB7
			9'd23 : rdata = 43'b1100010100000000000000000000000000011110000;
			// PEs: 8 -> 16
			// srcs: (30, 8)(865) 1312 --> (865) 1312:PUNB, pass, NI0
			9'd24 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 8 -> 23
			// srcs: (31, 9)(895) -23 --> (895) -23:PUNB, pass, PEGB7
			9'd25 : rdata = 43'b1100011011111000000000000000000000011110000;
			// PEs: 19 -> 24
			// srcs: (32, 33)(1108) 1058 --> (1108) 1058:PEGB3, pass, PUNB
			9'd26 : rdata = 43'b1100011100110000000000000000000001000000000;
			// PEs: 20 -> 24
			// srcs: (33, 34)(1138) 429 --> (1138) 429:PEGB4, pass, PUNB
			9'd27 : rdata = 43'b1100011101000000000000000000000001000000000;
			// PEs: 21 -> 24
			// srcs: (34, 35)(1168) 45 --> (1168) 45:PEGB5, pass, PUNB
			9'd28 : rdata = 43'b1100011101010000000000000000000001000000000;
			// PEs: 22 -> 24
			// srcs: (35, 36)(1198) 1488 --> (1198) 1488:PEGB6, pass, PUNB
			9'd29 : rdata = 43'b1100011101100000000000000000000001000000000;
			// PEs: 19 -> 24
			// srcs: (36, 37)(1109) 46 --> (1109) 46:PEGB3, pass, PUNB
			9'd30 : rdata = 43'b1100011100110000000000000000000001000000000;
			// PEs: 20 -> 24
			// srcs: (37, 38)(1139) 143 --> (1139) 143:PEGB4, pass, PUNB
			9'd31 : rdata = 43'b1100011101000000000000000000000001000000000;
			// PEs: 21 -> 24
			// srcs: (38, 39)(1169) 405 --> (1169) 405:PEGB5, pass, PUNB
			9'd32 : rdata = 43'b1100011101010000000000000000000001000000000;
			// PEs: 22 -> 24
			// srcs: (39, 40)(1199) -62 --> (1199) -62:PEGB6, pass, PUNB
			9'd33 : rdata = 43'b1100011101100000000000000000000001000000000;
			// PEs: 16 -> 23
			// srcs: (40, 10)(865) 1312 --> (865) 1312:NI0, pass, PEGB7
			9'd34 : rdata = 43'b1100010100000000000000000000000000011110000;
			// PEs: 8 -> 16
			// srcs: (41, 11)(925) 638 --> (925) 638:PUNB, pass, NI0
			9'd35 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 8 -> 23
			// srcs: (42, 12)(955) 462 --> (955) 462:PUNB, pass, PEGB7
			9'd36 : rdata = 43'b1100011011111000000000000000000000011110000;
			// PEs: 17 -> 24
			// srcs: (43, 41)(1050) 1332 --> (1050) 1332:PEGB1, pass, PUNB
			9'd37 : rdata = 43'b1100011100010000000000000000000001000000000;
			// PEs: 18 -> 24
			// srcs: (44, 42)(1080) 483 --> (1080) 483:PEGB2, pass, PUNB
			9'd38 : rdata = 43'b1100011100100000000000000000000001000000000;
			// PEs: 19 -> 24
			// srcs: (45, 43)(1110) 391 --> (1110) 391:PEGB3, pass, PUNB
			9'd39 : rdata = 43'b1100011100110000000000000000000001000000000;
			// PEs: 20 -> 24
			// srcs: (46, 44)(1140) 39 --> (1140) 39:PEGB4, pass, PUNB
			9'd40 : rdata = 43'b1100011101000000000000000000000001000000000;
			// PEs: 21 -> 24
			// srcs: (47, 45)(1170) -9 --> (1170) -9:PEGB5, pass, PUNB
			9'd41 : rdata = 43'b1100011101010000000000000000000001000000000;
			// PEs: 22 -> 24
			// srcs: (48, 46)(1200) 434 --> (1200) 434:PEGB6, pass, PUNB
			9'd42 : rdata = 43'b1100011101100000000000000000000001000000000;
			// PEs: 17 -> 24
			// srcs: (49, 59)(1051) 108 --> (1051) 108:PEGB1, pass, PUNB
			9'd43 : rdata = 43'b1100011100010000000000000000000001000000000;
			// PEs: 18 -> 24
			// srcs: (50, 60)(1081) 231 --> (1081) 231:PEGB2, pass, PUNB
			9'd44 : rdata = 43'b1100011100100000000000000000000001000000000;
			// PEs: 16 -> 23
			// srcs: (51, 13)(925) 638 --> (925) 638:NI0, pass, PEGB7
			9'd45 : rdata = 43'b1100010100000000000000000000000000011110000;
			// PEs: 8 -> 16
			// srcs: (52, 14)(985) 52 --> (985) 52:PUNB, pass, NI0
			9'd46 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 8 -> 23
			// srcs: (53, 15)(1015) 44 --> (1015) 44:PUNB, pass, PEGB7
			9'd47 : rdata = 43'b1100011011111000000000000000000000011110000;
			// PEs: 19 -> 24
			// srcs: (54, 61)(1111) 437 --> (1111) 437:PEGB3, pass, PUNB
			9'd48 : rdata = 43'b1100011100110000000000000000000001000000000;
			// PEs: 20 -> 24
			// srcs: (55, 62)(1141) 91 --> (1141) 91:PEGB4, pass, PUNB
			9'd49 : rdata = 43'b1100011101000000000000000000000001000000000;
			// PEs: 21 -> 24
			// srcs: (56, 63)(1171) 369 --> (1171) 369:PEGB5, pass, PUNB
			9'd50 : rdata = 43'b1100011101010000000000000000000001000000000;
			// PEs: 22 -> 24
			// srcs: (57, 64)(1201) 186 --> (1201) 186:PEGB6, pass, PUNB
			9'd51 : rdata = 43'b1100011101100000000000000000000001000000000;
			// PEs: 19 -> 24
			// srcs: (58, 77)(1112) 161 --> (1112) 161:PEGB3, pass, PUNB
			9'd52 : rdata = 43'b1100011100110000000000000000000001000000000;
			// PEs: 20 -> 24
			// srcs: (59, 78)(1142) 91 --> (1142) 91:PEGB4, pass, PUNB
			9'd53 : rdata = 43'b1100011101000000000000000000000001000000000;
			// PEs: 21 -> 24
			// srcs: (60, 79)(1172) 369 --> (1172) 369:PEGB5, pass, PUNB
			9'd54 : rdata = 43'b1100011101010000000000000000000001000000000;
			// PEs: 22 -> 24
			// srcs: (61, 80)(1202) 1333 --> (1202) 1333:PEGB6, pass, PUNB
			9'd55 : rdata = 43'b1100011101100000000000000000000001000000000;
			// PEs: 16 -> 23
			// srcs: (62, 16)(985) 52 --> (985) 52:NI0, pass, PEGB7
			9'd56 : rdata = 43'b1100010100000000000000000000000000011110000;
			// PEs: 19 -> 40
			// srcs: (63, 81)(1113) 299 --> (1113) 299:PEGB3, pass, PUGB5
			9'd57 : rdata = 43'b1100011100110000000000000000000000000001101;
			// PEs: 0 -> 16
			// srcs: (64, 47)(811) 279 --> (811) 279:PUGB0, pass, NI0
			9'd58 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 8 -> 23
			// srcs: (65, 48)(841) -96 --> (841) -96:PUNB, pass, PEGB7
			9'd59 : rdata = 43'b1100011011111000000000000000000000011110000;
			// PEs: 20 -> 40
			// srcs: (66, 82)(1143) 390 --> (1143) 390:PEGB4, pass, PUGB5
			9'd60 : rdata = 43'b1100011101000000000000000000000000000001101;
			// PEs: 21 -> 40
			// srcs: (67, 83)(1173) 36 --> (1173) 36:PEGB5, pass, PUGB5
			9'd61 : rdata = 43'b1100011101010000000000000000000000000001101;
			// PEs: 22 -> 40
			// srcs: (68, 84)(1203) 527 --> (1203) 527:PEGB6, pass, PUGB5
			9'd62 : rdata = 43'b1100011101100000000000000000000000000001101;
			// PEs: 17 -> 24
			// srcs: (69, 85)(1054) 1188 --> (1054) 1188:PEGB1, pass, PUNB
			9'd63 : rdata = 43'b1100011100010000000000000000000001000000000;
			// PEs: 18 -> 24
			// srcs: (70, 86)(1084) 525 --> (1084) 525:PEGB2, pass, PUNB
			9'd64 : rdata = 43'b1100011100100000000000000000000001000000000;
			// PEs: 19 -> 24
			// srcs: (71, 87)(1114) 483 --> (1114) 483:PEGB3, pass, PUNB
			9'd65 : rdata = 43'b1100011100110000000000000000000001000000000;
			// PEs: 20 -> 24
			// srcs: (72, 88)(1144) 13 --> (1144) 13:PEGB4, pass, PUNB
			9'd66 : rdata = 43'b1100011101000000000000000000000001000000000;
			// PEs: 21 -> 24
			// srcs: (73, 89)(1174) 162 --> (1174) 162:PEGB5, pass, PUNB
			9'd67 : rdata = 43'b1100011101010000000000000000000001000000000;
			// PEs: 16 -> 23
			// srcs: (74, 49)(811) 279 --> (811) 279:NI0, pass, PEGB7
			9'd68 : rdata = 43'b1100010100000000000000000000000000011110000;
			// PEs: 8 -> 16
			// srcs: (75, 50)(871) 928 --> (871) 928:PUNB, pass, NI0
			9'd69 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 8 -> 23
			// srcs: (76, 51)(901) -47 --> (901) -47:PUNB, pass, PEGB7
			9'd70 : rdata = 43'b1100011011111000000000000000000000011110000;
			// PEs: 22 -> 24
			// srcs: (77, 90)(1204) 1302 --> (1204) 1302:PEGB6, pass, PUNB
			9'd71 : rdata = 43'b1100011101100000000000000000000001000000000;
			// PEs: 19 -> 56
			// srcs: (78, 91)(1115) 69 --> (1115) 69:PEGB3, pass, PUGB7
			9'd72 : rdata = 43'b1100011100110000000000000000000000000001111;
			// PEs: 20 -> 56
			// srcs: (79, 92)(1145) 312 --> (1145) 312:PEGB4, pass, PUGB7
			9'd73 : rdata = 43'b1100011101000000000000000000000000000001111;
			// PEs: 21 -> 56
			// srcs: (80, 93)(1175) 198 --> (1175) 198:PEGB5, pass, PUGB7
			9'd74 : rdata = 43'b1100011101010000000000000000000000000001111;
			// PEs: 22 -> 56
			// srcs: (81, 94)(1205) 31 --> (1205) 31:PEGB6, pass, PUGB7
			9'd75 : rdata = 43'b1100011101100000000000000000000000000001111;
			// PEs: 19 -> 24
			// srcs: (82, 107)(1116) 598 --> (1116) 598:PEGB3, pass, PUNB
			9'd76 : rdata = 43'b1100011100110000000000000000000001000000000;
			// PEs: 20 -> 24
			// srcs: (83, 108)(1146) 195 --> (1146) 195:PEGB4, pass, PUNB
			9'd77 : rdata = 43'b1100011101000000000000000000000001000000000;
			// PEs: 21 -> 24
			// srcs: (84, 109)(1176) 360 --> (1176) 360:PEGB5, pass, PUNB
			9'd78 : rdata = 43'b1100011101010000000000000000000001000000000;
			// PEs: 16 -> 23
			// srcs: (85, 52)(871) 928 --> (871) 928:NI0, pass, PEGB7
			9'd79 : rdata = 43'b1100010100000000000000000000000000011110000;
			// PEs: 8 -> 16
			// srcs: (86, 53)(931) 464 --> (931) 464:PUNB, pass, NI0
			9'd80 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 8 -> 23
			// srcs: (87, 54)(961) 363 --> (961) 363:PUNB, pass, PEGB7
			9'd81 : rdata = 43'b1100011011111000000000000000000000011110000;
			// PEs: 22 -> 24
			// srcs: (88, 110)(1206) 1178 --> (1206) 1178:PEGB6, pass, PUNB
			9'd82 : rdata = 43'b1100011101100000000000000000000001000000000;
			// PEs: 17 -> 24
			// srcs: (89, 123)(1057) 1080 --> (1057) 1080:PEGB1, pass, PUNB
			9'd83 : rdata = 43'b1100011100010000000000000000000001000000000;
			// PEs: 18 -> 24
			// srcs: (90, 124)(1087) 903 --> (1087) 903:PEGB2, pass, PUNB
			9'd84 : rdata = 43'b1100011100100000000000000000000001000000000;
			// PEs: 19 -> 24
			// srcs: (91, 125)(1117) 1035 --> (1117) 1035:PEGB3, pass, PUNB
			9'd85 : rdata = 43'b1100011100110000000000000000000001000000000;
			// PEs: 20 -> 24
			// srcs: (92, 126)(1147) 377 --> (1147) 377:PEGB4, pass, PUNB
			9'd86 : rdata = 43'b1100011101000000000000000000000001000000000;
			// PEs: 21 -> 24
			// srcs: (93, 127)(1177) 396 --> (1177) 396:PEGB5, pass, PUNB
			9'd87 : rdata = 43'b1100011101010000000000000000000001000000000;
			// PEs: 22 -> 24
			// srcs: (94, 128)(1207) 372 --> (1207) 372:PEGB6, pass, PUNB
			9'd88 : rdata = 43'b1100011101100000000000000000000001000000000;
			// PEs: 19 -> 24
			// srcs: (95, 129)(1118) 391 --> (1118) 391:PEGB3, pass, PUNB
			9'd89 : rdata = 43'b1100011100110000000000000000000001000000000;
			// PEs: 16 -> 23
			// srcs: (96, 55)(931) 464 --> (931) 464:NI0, pass, PEGB7
			9'd90 : rdata = 43'b1100010100000000000000000000000000011110000;
			// PEs: 8 -> 16
			// srcs: (97, 56)(991) 50 --> (991) 50:PUNB, pass, NI0
			9'd91 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 8 -> 23
			// srcs: (98, 57)(1021) 880 --> (1021) 880:PUNB, pass, PEGB7
			9'd92 : rdata = 43'b1100011011111000000000000000000000011110000;
			// PEs: 20 -> 24
			// srcs: (99, 130)(1148) 273 --> (1148) 273:PEGB4, pass, PUNB
			9'd93 : rdata = 43'b1100011101000000000000000000000001000000000;
			// PEs: 21 -> 24
			// srcs: (100, 131)(1178) 81 --> (1178) 81:PEGB5, pass, PUNB
			9'd94 : rdata = 43'b1100011101010000000000000000000001000000000;
			// PEs: 22 -> 24
			// srcs: (101, 132)(1208) -62 --> (1208) -62:PEGB6, pass, PUNB
			9'd95 : rdata = 43'b1100011101100000000000000000000001000000000;
			// PEs: 19 -> 24
			// srcs: (102, 133)(1119) 322 --> (1119) 322:PEGB3, pass, PUNB
			9'd96 : rdata = 43'b1100011100110000000000000000000001000000000;
			// PEs: 20 -> 24
			// srcs: (103, 134)(1149) 429 --> (1149) 429:PEGB4, pass, PUNB
			9'd97 : rdata = 43'b1100011101000000000000000000000001000000000;
			// PEs: 21 -> 24
			// srcs: (104, 135)(1179) 333 --> (1179) 333:PEGB5, pass, PUNB
			9'd98 : rdata = 43'b1100011101010000000000000000000001000000000;
			// PEs: 22 -> 24
			// srcs: (105, 136)(1209) 806 --> (1209) 806:PEGB6, pass, PUNB
			9'd99 : rdata = 43'b1100011101100000000000000000000001000000000;
			// PEs: 17 -> 24
			// srcs: (106, 137)(1060) 720 --> (1060) 720:PEGB1, pass, PUNB
			9'd100 : rdata = 43'b1100011100010000000000000000000001000000000;
			// PEs: 16 -> 23
			// srcs: (107, 58)(991) 50 --> (991) 50:NI0, pass, PEGB7
			9'd101 : rdata = 43'b1100010100000000000000000000000000011110000;
			// PEs: 0 -> 16
			// srcs: (108, 65)(812) 1457 --> (812) 1457:PUGB0, pass, NI0
			9'd102 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 8 -> 23
			// srcs: (109, 66)(842) 416 --> (842) 416:PUNB, pass, PEGB7
			9'd103 : rdata = 43'b1100011011111000000000000000000000011110000;
			// PEs: 18 -> 24
			// srcs: (110, 138)(1090) 588 --> (1090) 588:PEGB2, pass, PUNB
			9'd104 : rdata = 43'b1100011100100000000000000000000001000000000;
			// PEs: 19 -> 24
			// srcs: (111, 139)(1120) 437 --> (1120) 437:PEGB3, pass, PUNB
			9'd105 : rdata = 43'b1100011100110000000000000000000001000000000;
			// PEs: 20 -> 24
			// srcs: (112, 140)(1150) 559 --> (1150) 559:PEGB4, pass, PUNB
			9'd106 : rdata = 43'b1100011101000000000000000000000001000000000;
			// PEs: 21 -> 24
			// srcs: (113, 141)(1180) 261 --> (1180) 261:PEGB5, pass, PUNB
			9'd107 : rdata = 43'b1100011101010000000000000000000001000000000;
			// PEs: 22 -> 24
			// srcs: (114, 142)(1210) 1209 --> (1210) 1209:PEGB6, pass, PUNB
			9'd108 : rdata = 43'b1100011101100000000000000000000001000000000;
			// PEs: 17 -> 56
			// srcs: (115, 143)(1061) 504 --> (1061) 504:PEGB1, pass, PUGB7
			9'd109 : rdata = 43'b1100011100010000000000000000000000000001111;
			// PEs: 18 -> 56
			// srcs: (116, 144)(1091) 126 --> (1091) 126:PEGB2, pass, PUGB7
			9'd110 : rdata = 43'b1100011100100000000000000000000000000001111;
			// PEs: 19 -> 56
			// srcs: (117, 145)(1121) 966 --> (1121) 966:PEGB3, pass, PUGB7
			9'd111 : rdata = 43'b1100011100110000000000000000000000000001111;
			// PEs: 16 -> 23
			// srcs: (118, 67)(812) 1457 --> (812) 1457:NI0, pass, PEGB7
			9'd112 : rdata = 43'b1100010100000000000000000000000000011110000;
			// PEs: 8 -> 16
			// srcs: (119, 68)(872) 1024 --> (872) 1024:PUNB, pass, NI0
			9'd113 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 8 -> 23
			// srcs: (120, 69)(902) -45 --> (902) -45:PUNB, pass, PEGB7
			9'd114 : rdata = 43'b1100011011111000000000000000000000011110000;
			// PEs: 20 -> 56
			// srcs: (121, 146)(1151) 533 --> (1151) 533:PEGB4, pass, PUGB7
			9'd115 : rdata = 43'b1100011101000000000000000000000000000001111;
			// PEs: 21 -> 56
			// srcs: (122, 147)(1181) 378 --> (1181) 378:PEGB5, pass, PUGB7
			9'd116 : rdata = 43'b1100011101010000000000000000000000000001111;
			// PEs: 22 -> 56
			// srcs: (123, 148)(1211) 1333 --> (1211) 1333:PEGB6, pass, PUGB7
			9'd117 : rdata = 43'b1100011101100000000000000000000000000001111;
			// PEs: 17 -> 24
			// srcs: (124, 149)(1062) 612 --> (1062) 612:PEGB1, pass, PUNB
			9'd118 : rdata = 43'b1100011100010000000000000000000001000000000;
			// PEs: 18 -> 24
			// srcs: (125, 150)(1092) 672 --> (1092) 672:PEGB2, pass, PUNB
			9'd119 : rdata = 43'b1100011100100000000000000000000001000000000;
			// PEs: 19 -> 24
			// srcs: (126, 151)(1122) 920 --> (1122) 920:PEGB3, pass, PUNB
			9'd120 : rdata = 43'b1100011100110000000000000000000001000000000;
			// PEs: 20 -> 24
			// srcs: (127, 152)(1152) 312 --> (1152) 312:PEGB4, pass, PUNB
			9'd121 : rdata = 43'b1100011101000000000000000000000001000000000;
			// PEs: 21 -> 24
			// srcs: (128, 153)(1182) 297 --> (1182) 297:PEGB5, pass, PUNB
			9'd122 : rdata = 43'b1100011101010000000000000000000001000000000;
			// PEs: 16 -> 23
			// srcs: (129, 70)(872) 1024 --> (872) 1024:NI0, pass, PEGB7
			9'd123 : rdata = 43'b1100010100000000000000000000000000011110000;
			// PEs: 8 -> 16
			// srcs: (130, 71)(932) 580 --> (932) 580:PUNB, pass, NI0
			9'd124 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 8 -> 23
			// srcs: (131, 72)(962) 99 --> (962) 99:PUNB, pass, PEGB7
			9'd125 : rdata = 43'b1100011011111000000000000000000000011110000;
			// PEs: 22 -> 24
			// srcs: (132, 154)(1212) 1085 --> (1212) 1085:PEGB6, pass, PUNB
			9'd126 : rdata = 43'b1100011101100000000000000000000001000000000;
			// PEs: 19 -> 8
			// srcs: (133, 167)(1123) 851 --> (1123) 851:PEGB3, pass, PUGB1
			9'd127 : rdata = 43'b1100011100110000000000000000000000000001001;
			// PEs: 20 -> 8
			// srcs: (134, 168)(1153) 377 --> (1153) 377:PEGB4, pass, PUGB1
			9'd128 : rdata = 43'b1100011101000000000000000000000000000001001;
			// PEs: 21 -> 8
			// srcs: (135, 169)(1183) 72 --> (1183) 72:PEGB5, pass, PUGB1
			9'd129 : rdata = 43'b1100011101010000000000000000000000000001001;
			// PEs: 22 -> 8
			// srcs: (136, 170)(1213) 775 --> (1213) 775:PEGB6, pass, PUGB1
			9'd130 : rdata = 43'b1100011101100000000000000000000000000001001;
			// PEs: 19 -> 24
			// srcs: (137, 180)(1124) 1127 --> (1124) 1127:PEGB3, pass, PUNB
			9'd131 : rdata = 43'b1100011100110000000000000000000001000000000;
			// PEs: 20 -> 24
			// srcs: (138, 181)(1154) 273 --> (1154) 273:PEGB4, pass, PUNB
			9'd132 : rdata = 43'b1100011101000000000000000000000001000000000;
			// PEs: 21 -> 24
			// srcs: (139, 182)(1184) 81 --> (1184) 81:PEGB5, pass, PUNB
			9'd133 : rdata = 43'b1100011101010000000000000000000001000000000;
			// PEs: 16 -> 23
			// srcs: (140, 73)(932) 580 --> (932) 580:NI0, pass, PEGB7
			9'd134 : rdata = 43'b1100010100000000000000000000000000011110000;
			// PEs: 8 -> 16
			// srcs: (141, 74)(992) 50 --> (992) 50:PUNB, pass, NI0
			9'd135 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 8 -> 23
			// srcs: (142, 75)(1022) 66 --> (1022) 66:PUNB, pass, PEGB7
			9'd136 : rdata = 43'b1100011011111000000000000000000000011110000;
			// PEs: 22 -> 24
			// srcs: (143, 183)(1214) -31 --> (1214) -31:PEGB6, pass, PUNB
			9'd137 : rdata = 43'b1100011101100000000000000000000001000000000;
			// PEs: 17 -> 24
			// srcs: (144, 193)(1065) 864 --> (1065) 864:PEGB1, pass, PUNB
			9'd138 : rdata = 43'b1100011100010000000000000000000001000000000;
			// PEs: 18 -> 24
			// srcs: (145, 194)(1095) 609 --> (1095) 609:PEGB2, pass, PUNB
			9'd139 : rdata = 43'b1100011100100000000000000000000001000000000;
			// PEs: 19 -> 24
			// srcs: (146, 195)(1125) 138 --> (1125) 138:PEGB3, pass, PUNB
			9'd140 : rdata = 43'b1100011100110000000000000000000001000000000;
			// PEs: 20 -> 24
			// srcs: (147, 196)(1155) 0 --> (1155) 0:PEGB4, pass, PUNB
			9'd141 : rdata = 43'b1100011101000000000000000000000001000000000;
			// PEs: 21 -> 24
			// srcs: (148, 197)(1185) 144 --> (1185) 144:PEGB5, pass, PUNB
			9'd142 : rdata = 43'b1100011101010000000000000000000001000000000;
			// PEs: 22 -> 24
			// srcs: (149, 198)(1215) -93 --> (1215) -93:PEGB6, pass, PUNB
			9'd143 : rdata = 43'b1100011101100000000000000000000001000000000;
			// PEs: 19 -> 24
			// srcs: (150, 208)(1126) 897 --> (1126) 897:PEGB3, pass, PUNB
			9'd144 : rdata = 43'b1100011100110000000000000000000001000000000;
			// PEs: 16 -> 23
			// srcs: (151, 76)(992) 50 --> (992) 50:NI0, pass, PEGB7
			9'd145 : rdata = 43'b1100010100000000000000000000000000011110000;
			// PEs: 0 -> 16
			// srcs: (152, 95)(816) 341 --> (816) 341:PUGB0, pass, NI0
			9'd146 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 8 -> 23
			// srcs: (153, 96)(846) 448 --> (846) 448:PUNB, pass, PEGB7
			9'd147 : rdata = 43'b1100011011111000000000000000000000011110000;
			// PEs: 20 -> 24
			// srcs: (154, 209)(1156) 39 --> (1156) 39:PEGB4, pass, PUNB
			9'd148 : rdata = 43'b1100011101000000000000000000000001000000000;
			// PEs: 21 -> 24
			// srcs: (155, 210)(1186) 198 --> (1186) 198:PEGB5, pass, PUNB
			9'd149 : rdata = 43'b1100011101010000000000000000000001000000000;
			// PEs: 22 -> 24
			// srcs: (156, 211)(1216) 341 --> (1216) 341:PEGB6, pass, PUNB
			9'd150 : rdata = 43'b1100011101100000000000000000000001000000000;
			// PEs: 19 -> 24
			// srcs: (157, 221)(1127) 989 --> (1127) 989:PEGB3, pass, PUNB
			9'd151 : rdata = 43'b1100011100110000000000000000000001000000000;
			// PEs: 20 -> 24
			// srcs: (158, 222)(1157) 195 --> (1157) 195:PEGB4, pass, PUNB
			9'd152 : rdata = 43'b1100011101000000000000000000000001000000000;
			// PEs: 21 -> 24
			// srcs: (159, 223)(1187) 441 --> (1187) 441:PEGB5, pass, PUNB
			9'd153 : rdata = 43'b1100011101010000000000000000000001000000000;
			// PEs: 22 -> 24
			// srcs: (160, 224)(1217) 310 --> (1217) 310:PEGB6, pass, PUNB
			9'd154 : rdata = 43'b1100011101100000000000000000000001000000000;
			// PEs: 23 -> 40
			// srcs: (161, 225)(1227) 2387 --> (1227) 2387:PENB, pass, PUGB5
			9'd155 : rdata = 43'b1100011011110000000000000000000000000001101;
			// PEs: 16 -> 23
			// srcs: (162, 97)(816) 341 --> (816) 341:NI0, pass, PEGB7
			9'd156 : rdata = 43'b1100010100000000000000000000000000011110000;
			// PEs: 8 -> 16
			// srcs: (163, 98)(876) 704 --> (876) 704:PUNB, pass, NI0
			9'd157 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 8 -> 23
			// srcs: (164, 99)(906) -28 --> (906) -28:PUNB, pass, PEGB7
			9'd158 : rdata = 43'b1100011011111000000000000000000000011110000;
			// PEs: 23 -> 24
			// srcs: (165, 227)(1246) 962 --> (1246) 962:PENB, pass, PUNB
			9'd159 : rdata = 43'b1100011011110000000000000000000001000000000;
			// PEs: 23 -> 24
			// srcs: (166, 230)(1360) 183 --> (1360) 183:PENB, pass, PUNB
			9'd160 : rdata = 43'b1100011011110000000000000000000001000000000;
			// PEs: 23 -> 24
			// srcs: (167, 231)(1363) 930 --> (1363) 930:PENB, pass, PUNB
			9'd161 : rdata = 43'b1100011011110000000000000000000001000000000;
			// PEs: 23 -> 48
			// srcs: (168, 232)(1379) 1873 --> (1379) 1873:PENB, pass, PUGB6
			9'd162 : rdata = 43'b1100011011110000000000000000000000000001110;
			// PEs: 23 -> 24
			// srcs: (169, 235)(1455) 789 --> (1455) 789:PENB, pass, PUNB
			9'd163 : rdata = 43'b1100011011110000000000000000000001000000000;
			// PEs: 23 -> 40
			// srcs: (170, 226)(1231) 756 --> (1231) 756:PENB, pass, PUGB5
			9'd164 : rdata = 43'b1100011011110000000000000000000000000001101;
			// PEs: 23 -> 56
			// srcs: (172, 228)(1307) 1302 --> (1307) 1302:PENB, pass, PUGB7
			9'd165 : rdata = 43'b1100011011110000000000000000000000000001111;
			// PEs: 16 -> 23
			// srcs: (173, 100)(876) 704 --> (876) 704:NI0, pass, PEGB7
			9'd166 : rdata = 43'b1100010100000000000000000000000000011110000;
			// PEs: 8 -> 16
			// srcs: (174, 101)(936) 290 --> (936) 290:PUNB, pass, NI0
			9'd167 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 8 -> 23
			// srcs: (175, 102)(966) 1518 --> (966) 1518:PUNB, pass, PEGB7
			9'd168 : rdata = 43'b1100011011111000000000000000000000011110000;
			// PEs: 23 -> 0
			// srcs: (176, 229)(1326) 1131 --> (1326) 1131:PENB, pass, PUGB0
			9'd169 : rdata = 43'b1100011011110000000000000000000000000001000;
			// PEs: 23 -> 40
			// srcs: (177, 233)(1402) 1053 --> (1402) 1053:PENB, pass, PUGB5
			9'd170 : rdata = 43'b1100011011110000000000000000000000000001101;
			// PEs: 23 -> 32
			// srcs: (178, 234)(1440) 1572 --> (1440) 1572:PENB, pass, PUGB4
			9'd171 : rdata = 43'b1100011011110000000000000000000000000001100;
			// PEs: 23 -> 40
			// srcs: (183, 238)(1497) 1764 --> (1497) 1764:PENB, pass, PUGB5
			9'd172 : rdata = 43'b1100011011110000000000000000000000000001101;
			// PEs: 16 -> 23
			// srcs: (184, 103)(936) 290 --> (936) 290:NI0, pass, PEGB7
			9'd173 : rdata = 43'b1100010100000000000000000000000000011110000;
			// PEs: 8 -> 16
			// srcs: (185, 104)(996) 64 --> (996) 64:PUNB, pass, NI0
			9'd174 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 8 -> 23
			// srcs: (186, 105)(1026) -22 --> (1026) -22:PUNB, pass, PEGB7
			9'd175 : rdata = 43'b1100011011111000000000000000000000011110000;
			// PEs: 23 -> 32
			// srcs: (187, 239)(1516) 474 --> (1516) 474:PENB, pass, PUGB4
			9'd176 : rdata = 43'b1100011011110000000000000000000000000001100;
			// PEs: 17 -> 32
			// srcs: (188, 275)(1751) 2005 --> (1751) 2005:PEGB1, pass, PUGB4
			9'd177 : rdata = 43'b1100011100010000000000000000000000000001100;
			// PEs: 20 -> 32
			// srcs: (189, 277)(1789) 2117 --> (1789) 2117:PEGB4, pass, PUGB4
			9'd178 : rdata = 43'b1100011101000000000000000000000000000001100;
			// PEs: 16 -> 23
			// srcs: (195, 106)(996) 64 --> (996) 64:NI0, pass, PEGB7
			9'd179 : rdata = 43'b1100010100000000000000000000000000011110000;
			// PEs: 0 -> 16
			// srcs: (196, 111)(817) 372 --> (817) 372:PUGB0, pass, NI0
			9'd180 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 8 -> 23
			// srcs: (197, 112)(847) 1568 --> (847) 1568:PUNB, pass, PEGB7
			9'd181 : rdata = 43'b1100011011111000000000000000000000011110000;
			// PEs: 0 -> 16
			// srcs: (198, 155)(823) 620 --> (823) 620:PUGB0, pass, NI1
			9'd182 : rdata = 43'b1100011100001000000001000010000000000000000;
			// PEs: 16 -> 23
			// srcs: (206, 113)(817) 372 --> (817) 372:NI0, pass, PEGB7
			9'd183 : rdata = 43'b1100010100000000000000000000000000011110000;
			// PEs: 8 -> 16
			// srcs: (207, 114)(877) 1024 --> (877) 1024:PUNB, pass, NI0
			9'd184 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 8 -> 23
			// srcs: (208, 115)(907) -13 --> (907) -13:PUNB, pass, PEGB7
			9'd185 : rdata = 43'b1100011011111000000000000000000000011110000;
			// PEs: 23 -> 24
			// srcs: (213, 236)(1474) 1940 --> (1474) 1940:PENB, pass, PUNB
			9'd186 : rdata = 43'b1100011011110000000000000000000001000000000;
			// PEs: 16 -> 23
			// srcs: (217, 116)(877) 1024 --> (877) 1024:NI0, pass, PEGB7
			9'd187 : rdata = 43'b1100010100000000000000000000000000011110000;
			// PEs: 8 -> 16
			// srcs: (218, 117)(937) 551 --> (937) 551:PUNB, pass, NI0
			9'd188 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 8 -> 23
			// srcs: (219, 118)(967) 1485 --> (967) 1485:PUNB, pass, PEGB7
			9'd189 : rdata = 43'b1100011011111000000000000000000000011110000;
			// PEs: 16 -> 23
			// srcs: (228, 119)(937) 551 --> (937) 551:NI0, pass, PEGB7
			9'd190 : rdata = 43'b1100010100000000000000000000000000011110000;
			// PEs: 8 -> 16
			// srcs: (229, 120)(997) 78 --> (997) 78:PUNB, pass, NI0
			9'd191 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 8 -> 23
			// srcs: (230, 121)(1027) 792 --> (1027) 792:PUNB, pass, PEGB7
			9'd192 : rdata = 43'b1100011011111000000000000000000000011110000;
			// PEs: 8 -> 18
			// srcs: (231, 156)(853) 160 --> (853) 160:PUNB, pass, PEGB2
			9'd193 : rdata = 43'b1100011011111000000000000000000000010100000;
			// PEs: 16 -> 23
			// srcs: (239, 122)(997) 78 --> (997) 78:NI0, pass, PEGB7
			9'd194 : rdata = 43'b1100010100000000000000000000000000011110000;
			// PEs: 16 -> 18
			// srcs: (240, 157)(823) 620 --> (823) 620:NI1, pass, PEGB2
			9'd195 : rdata = 43'b1100010100001000000000000000000000010100000;
			// PEs: 8 -> 16
			// srcs: (241, 158)(883) -96 --> (883) -96:PUNB, pass, NI0
			9'd196 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 8 -> 18
			// srcs: (242, 159)(913) -30 --> (913) -30:PUNB, pass, PEGB2
			9'd197 : rdata = 43'b1100011011111000000000000000000000010100000;
			// PEs: 23 -> 24
			// srcs: (246, 237)(1477) 870 --> (1477) 870:PENB, pass, PUNB
			9'd198 : rdata = 43'b1100011011110000000000000000000001000000000;
			// PEs: 16 -> 18
			// srcs: (251, 160)(883) -96 --> (883) -96:NI0, pass, PEGB2
			9'd199 : rdata = 43'b1100010100000000000000000000000000010100000;
			// PEs: 8 -> 16
			// srcs: (252, 161)(943) 203 --> (943) 203:PUNB, pass, NI0
			9'd200 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 8 -> 18
			// srcs: (253, 162)(973) 363 --> (973) 363:PUNB, pass, PEGB2
			9'd201 : rdata = 43'b1100011011111000000000000000000000010100000;
			// PEs: 23 -> 24
			// srcs: (254, 248)(1232) 613 --> (1232) 613:PENB, pass, PUNB
			9'd202 : rdata = 43'b1100011011110000000000000000000001000000000;
			// PEs: 23 -> 24
			// srcs: (259, 250)(1369) 1708 --> (1369) 1708:PENB, pass, PUNB
			9'd203 : rdata = 43'b1100011011110000000000000000000001000000000;
			// PEs: 16 -> 18
			// srcs: (262, 163)(943) 203 --> (943) 203:NI0, pass, PEGB2
			9'd204 : rdata = 43'b1100010100000000000000000000000000010100000;
			// PEs: 8 -> 16
			// srcs: (263, 164)(1003) 94 --> (1003) 94:PUNB, pass, NI0
			9'd205 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 8 -> 18
			// srcs: (264, 165)(1033) 638 --> (1033) 638:PUNB, pass, PEGB2
			9'd206 : rdata = 43'b1100011011111000000000000000000000010100000;
			// PEs: 8 -> 16
			// srcs: (265, 171)(884) 640 --> (884) 640:PUNB, pass, NI1
			9'd207 : rdata = 43'b1100011011111000000001000010000000000000000;
			// PEs: 8 -> 17
			// srcs: (266, 172)(914) -19 --> (914) -19:PUNB, pass, PENB
			9'd208 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 23 -> 24
			// srcs: (267, 251)(1483) 3047 --> (1483) 3047:PENB, pass, PUNB
			9'd209 : rdata = 43'b1100011011110000000000000000000001000000000;
			// PEs: 17 -> 24
			// srcs: (268, 272)(1694) 840 --> (1694) 840:PEGB1, pass, PUNB
			9'd210 : rdata = 43'b1100011100010000000000000000000001000000000;
			// PEs: 19 -> 24
			// srcs: (269, 273)(1713) 2173 --> (1713) 2173:PEGB3, pass, PUNB
			9'd211 : rdata = 43'b1100011100110000000000000000000001000000000;
			// PEs: 17 -> 24
			// srcs: (270, 278)(1259) 3298 --> (1259) 3298:PEGB1, pass, PUNB
			9'd212 : rdata = 43'b1100011100010000000000000000000001000000000;
			// PEs: 16 -> 17
			// srcs: (272, 173)(884) 640 --> (884) 640:NI1, pass, PENB
			9'd213 : rdata = 43'b1100010100001000000000000000000000100000000;
			// PEs: 16 -> 18
			// srcs: (273, 166)(1003) 94 --> (1003) 94:NI0, pass, PEGB2
			9'd214 : rdata = 43'b1100010100000000000000000000000000010100000;
			// PEs: 8 -> 16
			// srcs: (274, 174)(944) 580 --> (944) 580:PUNB, pass, NI0
			9'd215 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 8 -> 17
			// srcs: (275, 175)(974) 759 --> (974) 759:PUNB, pass, PENB
			9'd216 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 16 -> 17
			// srcs: (281, 176)(944) 580 --> (944) 580:NI0, pass, PENB
			9'd217 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 8 -> 16
			// srcs: (282, 177)(1004) 32 --> (1004) 32:PUNB, pass, NI0
			9'd218 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 8 -> 17
			// srcs: (283, 178)(1034) 220 --> (1034) 220:PUNB, pass, PENB
			9'd219 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 16 -> 17
			// srcs: (289, 179)(1004) 32 --> (1004) 32:NI0, pass, PENB
			9'd220 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 8 -> 16
			// srcs: (290, 184)(885) 128 --> (885) 128:PUNB, pass, NI0
			9'd221 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 8 -> 17
			// srcs: (291, 185)(915) -2 --> (915) -2:PUNB, pass, PENB
			9'd222 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 16 -> 17
			// srcs: (297, 186)(885) 128 --> (885) 128:NI0, pass, PENB
			9'd223 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 8 -> 16
			// srcs: (298, 187)(945) 87 --> (945) 87:PUNB, pass, NI0
			9'd224 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 8 -> 17
			// srcs: (299, 188)(975) 1089 --> (975) 1089:PUNB, pass, PENB
			9'd225 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 16 -> 17
			// srcs: (305, 189)(945) 87 --> (945) 87:NI0, pass, PENB
			9'd226 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 8 -> 16
			// srcs: (306, 190)(1005) 44 --> (1005) 44:PUNB, pass, NI0
			9'd227 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 8 -> 17
			// srcs: (307, 191)(1035) 330 --> (1035) 330:PUNB, pass, PENB
			9'd228 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 16 -> 17
			// srcs: (313, 192)(1005) 44 --> (1005) 44:NI0, pass, PENB
			9'd229 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 8 -> 16
			// srcs: (314, 199)(886) 1024 --> (886) 1024:PUNB, pass, NI0
			9'd230 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 8 -> 17
			// srcs: (315, 200)(916) -23 --> (916) -23:PUNB, pass, PENB
			9'd231 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 17 -> 8
			// srcs: (320, 241)(1629) 374 --> (1629) 374:PEGB1, pass, PUGB1
			9'd232 : rdata = 43'b1100011100010000000000000000000000000001001;
			// PEs: 16 -> 17
			// srcs: (321, 201)(886) 1024 --> (886) 1024:NI0, pass, PENB
			9'd233 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 8 -> 16
			// srcs: (322, 202)(946) 1421 --> (946) 1421:PUNB, pass, NI0
			9'd234 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 8 -> 17
			// srcs: (323, 203)(976) 891 --> (976) 891:PUNB, pass, PENB
			9'd235 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 23 -> 8
			// srcs: (328, 280)(1392) 2905 --> (1392) 2905:PENB, pass, PUGB1
			9'd236 : rdata = 43'b1100011011110000000000000000000000000001001;
			// PEs: 16 -> 17
			// srcs: (329, 204)(946) 1421 --> (946) 1421:NI0, pass, PENB
			9'd237 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 8 -> 16
			// srcs: (330, 205)(1006) 70 --> (1006) 70:PUNB, pass, NI0
			9'd238 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 8 -> 17
			// srcs: (331, 206)(1036) 0 --> (1036) 0:PUNB, pass, PENB
			9'd239 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 16 -> 17
			// srcs: (337, 207)(1006) 70 --> (1006) 70:NI0, pass, PENB
			9'd240 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 8 -> 16
			// srcs: (338, 212)(887) 128 --> (887) 128:PUNB, pass, NI0
			9'd241 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 8 -> 17
			// srcs: (339, 213)(917) -39 --> (917) -39:PUNB, pass, PENB
			9'd242 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 16 -> 17
			// srcs: (345, 214)(887) 128 --> (887) 128:NI0, pass, PENB
			9'd243 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 8 -> 16
			// srcs: (346, 215)(947) 1015 --> (947) 1015:PUNB, pass, NI0
			9'd244 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 8 -> 17
			// srcs: (347, 216)(977) 132 --> (977) 132:PUNB, pass, PENB
			9'd245 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 16 -> 17
			// srcs: (353, 217)(947) 1015 --> (947) 1015:NI0, pass, PENB
			9'd246 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 8 -> 16
			// srcs: (354, 218)(1007) 72 --> (1007) 72:PUNB, pass, NI0
			9'd247 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 8 -> 17
			// srcs: (355, 219)(1037) 220 --> (1037) 220:PUNB, pass, PENB
			9'd248 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 16 -> 17
			// srcs: (361, 220)(1007) 72 --> (1007) 72:NI0, pass, PENB
			9'd249 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 8 -> 17
			// srcs: (362, 240)(1587) 23 --> (1587) 23:PUNB, pass, PENB
			9'd250 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 8 -> 17
			// srcs: (363, 242)(1686) 724 --> (1686) 724:PUNB, pass, PENB
			9'd251 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 8 -> 17
			// srcs: (364, 243)(1705) 358 --> (1705) 358:PUNB, pass, PENB
			9'd252 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 8 -> 17
			// srcs: (365, 244)(1724) 482 --> (1724) 482:PUNB, pass, PENB
			9'd253 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 8 -> 17
			// srcs: (366, 245)(1743) 560 --> (1743) 560:PUNB, pass, PENB
			9'd254 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 8 -> 17
			// srcs: (367, 246)(1762) 102 --> (1762) 102:PUNB, pass, PENB
			9'd255 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 8 -> 17
			// srcs: (368, 247)(1781) 536 --> (1781) 536:PUNB, pass, PENB
			9'd256 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 8 -> 22
			// srcs: (369, 249)(1595) 941 --> (1595) 941:PUNB, pass, PEGB6
			9'd257 : rdata = 43'b1100011011111000000000000000000000011100000;
			// PEs: 17 -> 0
			// srcs: (374, 256)(1750) 917 --> (1750) 917:PEGB1, pass, PUGB0
			9'd258 : rdata = 43'b1100011100010000000000000000000000000001000;
			// PEs: 8 -> 17
			// srcs: (510, 252)(1636) 1847 --> (1636) 1847:PUNB, pass, PENB
			9'd259 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 8 -> 17
			// srcs: (512, 253)(1692) 1410 --> (1692) 1410:PUNB, pass, PENB
			9'd260 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 8 -> 17
			// srcs: (513, 254)(1711) 1614 --> (1711) 1614:PUNB, pass, PENB
			9'd261 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 17 -> 56
			// srcs: (518, 286)(1639) 3149 --> (1639) 3149:PEGB1, pass, PUGB7
			9'd262 : rdata = 43'b1100011100010000000000000000000000000001111;
			// PEs: 17 -> 24
			// srcs: (519, 289)(1696) 2251 --> (1696) 2251:PEGB1, pass, PUNB
			9'd263 : rdata = 43'b1100011100010000000000000000000001000000000;
			// PEs: 17 -> 24
			// srcs: (520, 290)(1715) 3592 --> (1715) 3592:PEGB1, pass, PUNB
			9'd264 : rdata = 43'b1100011100010000000000000000000001000000000;
			// PEs: 8 -> 17
			// srcs: (998, 255)(1730) 2549 --> (1730) 2549:PUNB, pass, PENB
			9'd265 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 8 -> 17
			// srcs: (999, 257)(1768) 3151 --> (1768) 3151:PUNB, pass, PENB
			9'd266 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 8 -> 17
			// srcs: (1000, 258)(1787) 2303 --> (1787) 2303:PUNB, pass, PENB
			9'd267 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 24 -> 16
			// srcs: (1001, 259)(1333) 532 --> (1333) 532:PUGB3, pass, NI0
			9'd268 : rdata = 43'b1100011100111000000001000000000000000000000;
			// PEs: 56 -> 17
			// srcs: (1002, 260)(1334) 3857 --> (1334) 3857:PUGB7, pass, PENB
			9'd269 : rdata = 43'b1100011101111000000000000000000000100000000;
			// PEs: 17 -> 0
			// srcs: (1007, 291)(1791) 3445 --> (1791) 3445:PEGB1, pass, PUGB0
			9'd270 : rdata = 43'b1100011100010000000000000000000000000001000;
			// PEs: 16 -> 17
			// srcs: (1008, 261)(1333) 532 --> (1333) 532:NI0, pass, PENB
			9'd271 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 24 -> 16
			// srcs: (1009, 262)(1523) 1890 --> (1523) 1890:PUGB3, pass, NI0
			9'd272 : rdata = 43'b1100011100111000000001000000000000000000000;
			// PEs: 32 -> 17
			// srcs: (1010, 263)(1524) 4683 --> (1524) 4683:PUGB4, pass, PENB
			9'd273 : rdata = 43'b1100011101001000000000000000000000100000000;
			// PEs: 17 -> 40
			// srcs: (1015, 279)(1336) 4389 --> (1336) 4389:PEGB1, pass, PUGB5
			9'd274 : rdata = 43'b1100011100010000000000000000000000000001101;
			// PEs: 16 -> 17
			// srcs: (1016, 264)(1523) 1890 --> (1523) 1890:NI0, pass, PENB
			9'd275 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 24 -> 16
			// srcs: (1017, 265)(1542) 2466 --> (1542) 2466:PUGB3, pass, NI0
			9'd276 : rdata = 43'b1100011100111000000001000000000000000000000;
			// PEs: 40 -> 17
			// srcs: (1018, 266)(1543) 4164 --> (1543) 4164:PUGB5, pass, PENB
			9'd277 : rdata = 43'b1100011101011000000000000000000000100000000;
			// PEs: 23 -> 40
			// srcs: (1023, 281)(1468) 3219 --> (1468) 3219:PENB, pass, PUGB5
			9'd278 : rdata = 43'b1100011011110000000000000000000000000001101;
			// PEs: 16 -> 17
			// srcs: (1024, 267)(1542) 2466 --> (1542) 2466:NI0, pass, PENB
			9'd279 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 24 -> 16
			// srcs: (1025, 268)(1580) 2614 --> (1580) 2614:PUGB3, pass, NI0
			9'd280 : rdata = 43'b1100011100111000000001000000000000000000000;
			// PEs: 56 -> 17
			// srcs: (1026, 269)(1581) 6146 --> (1581) 6146:PUGB7, pass, PENB
			9'd281 : rdata = 43'b1100011101111000000000000000000000100000000;
			// PEs: 17 -> 48
			// srcs: (1027, 282)(1526) 6573 --> (1526) 6573:PEGB1, pass, PUGB6
			9'd282 : rdata = 43'b1100011100010000000000000000000000000001110;
			// PEs: 17 -> 48
			// srcs: (1031, 283)(1545) 6630 --> (1545) 6630:PEGB1, pass, PUGB6
			9'd283 : rdata = 43'b1100011100010000000000000000000000000001110;
			// PEs: 16 -> 17
			// srcs: (1032, 270)(1580) 2614 --> (1580) 2614:NI0, pass, PENB
			9'd284 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 8 -> 17
			// srcs: (1033, 271)(1599) 2075 --> (1599) 2075:PUNB, pass, PENB
			9'd285 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 8 -> 17
			// srcs: (1034, 274)(1733) 5670 --> (1733) 5670:PUNB, pass, PENB
			9'd286 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 8 -> 17
			// srcs: (1035, 276)(1771) 6226 --> (1771) 6226:PUNB, pass, PENB
			9'd287 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 17 -> 48
			// srcs: (1039, 284)(1583) 8760 --> (1583) 8760:PEGB1, pass, PUGB6
			9'd288 : rdata = 43'b1100011100010000000000000000000000000001110;
			// PEs: 18 -> 48
			// srcs: (1040, 285)(1620) 2914 --> (1620) 2914:PEGB2, pass, PUGB6
			9'd289 : rdata = 43'b1100011100100000000000000000000000000001110;
			// PEs: 18 -> 56
			// srcs: (1041, 287)(1658) 5192 --> (1658) 5192:PEGB2, pass, PUGB7
			9'd290 : rdata = 43'b1100011100100000000000000000000000000001111;
			// PEs: 17 -> 56
			// srcs: (1049, 288)(1677) 3421 --> (1677) 3421:PEGB1, pass, PUGB7
			9'd291 : rdata = 43'b1100011100010000000000000000000000000001111;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 17) begin
	always @(*) begin
		case(address)
			// PEs: 17, 17 -> 23
			// srcs: (1, 0)(444) 0, (18) 36 --> (1044) 0:NW0, ND0, *, PEGB7
			9'd0 : rdata = 43'b0001101000000011000000000000000000011110000;
			// PEs: 17, 17 -> 23
			// srcs: (2, 1)(445) 15, (18) 36 --> (1045) 540:NW1, ND0, *, PEGB7
			9'd1 : rdata = 43'b0001101000001011000000000000000000011110000;
			// PEs: 17, 17 -> 16
			// srcs: (3, 2)(446) 32, (18) 36 --> (1046) 1152:NW2, ND0, *, PEGB0
			9'd2 : rdata = 43'b0001101000010011000000000000000000010000000;
			// PEs: 17, 17 -> 16
			// srcs: (4, 3)(447) 29, (18) 36 --> (1047) 1044:NW3, ND0, *, PEGB0
			9'd3 : rdata = 43'b0001101000011011000000000000000000010000000;
			// PEs: 17, 17 -> 23
			// srcs: (5, 4)(448) 14, (18) 36 --> (1048) 504:NW4, ND0, *, PEGB7
			9'd4 : rdata = 43'b0001101000100011000000000000000000011110000;
			// PEs: 17, 17 -> 23
			// srcs: (6, 5)(449) 11, (18) 36 --> (1049) 396:NW5, ND0, *, PEGB7
			9'd5 : rdata = 43'b0001101000101011000000000000000000011110000;
			// PEs: 17, 17 -> 16
			// srcs: (7, 6)(450) 37, (18) 36 --> (1050) 1332:NW6, ND0, *, PEGB0
			9'd6 : rdata = 43'b0001101000110011000000000000000000010000000;
			// PEs: 17, 17 -> 16
			// srcs: (8, 7)(451) 3, (18) 36 --> (1051) 108:NW7, ND0, *, PEGB0
			9'd7 : rdata = 43'b0001101000111011000000000000000000010000000;
			// PEs: 17, 17 -> 23
			// srcs: (9, 8)(452) 4, (18) 36 --> (1052) 144:NW8, ND0, *, PEGB7
			9'd8 : rdata = 43'b0001101001000011000000000000000000011110000;
			// PEs: 17, 17 -> 23
			// srcs: (10, 9)(453) 31, (18) 36 --> (1053) 1116:NW9, ND0, *, PEGB7
			9'd9 : rdata = 43'b0001101001001011000000000000000000011110000;
			// PEs: 17, 17 -> 16
			// srcs: (11, 10)(454) 33, (18) 36 --> (1054) 1188:NW10, ND0, *, PEGB0
			9'd10 : rdata = 43'b0001101001010011000000000000000000010000000;
			// PEs: 17, 17 -> 23
			// srcs: (12, 11)(455) 39, (18) 36 --> (1055) 1404:NW11, ND0, *, PEGB7
			9'd11 : rdata = 43'b0001101001011011000000000000000000011110000;
			// PEs: 17, 17 -> 23
			// srcs: (13, 12)(456) 21, (18) 36 --> (1056) 756:NW12, ND0, *, PEGB7
			9'd12 : rdata = 43'b0001101001100011000000000000000000011110000;
			// PEs: 17, 17 -> 16
			// srcs: (14, 13)(457) 30, (18) 36 --> (1057) 1080:NW13, ND0, *, PEGB0
			9'd13 : rdata = 43'b0001101001101011000000000000000000010000000;
			// PEs: 17, 17 -> 23
			// srcs: (15, 14)(458) 35, (18) 36 --> (1058) 1260:NW14, ND0, *, PEGB7
			9'd14 : rdata = 43'b0001101001110011000000000000000000011110000;
			// PEs: 17, 17 -> 23
			// srcs: (16, 15)(459) 5, (18) 36 --> (1059) 180:NW15, ND0, *, PEGB7
			9'd15 : rdata = 43'b0001101001111011000000000000000000011110000;
			// PEs: 17, 17 -> 16
			// srcs: (17, 16)(460) 20, (18) 36 --> (1060) 720:NW16, ND0, *, PEGB0
			9'd16 : rdata = 43'b0001101010000011000000000000000000010000000;
			// PEs: 17, 17 -> 16
			// srcs: (18, 17)(461) 14, (18) 36 --> (1061) 504:NW17, ND0, *, PEGB0
			9'd17 : rdata = 43'b0001101010001011000000000000000000010000000;
			// PEs: 17, 17 -> 16
			// srcs: (19, 18)(462) 17, (18) 36 --> (1062) 612:NW18, ND0, *, PEGB0
			9'd18 : rdata = 43'b0001101010010011000000000000000000010000000;
			// PEs: 17, 17 -> 23
			// srcs: (20, 19)(463) 0, (18) 36 --> (1063) 0:NW19, ND0, *, PEGB7
			9'd19 : rdata = 43'b0001101010011011000000000000000000011110000;
			// PEs: 17, 17 -> 23
			// srcs: (21, 20)(464) 9, (18) 36 --> (1064) 324:NW20, ND0, *, PEGB7
			9'd20 : rdata = 43'b0001101010100011000000000000000000011110000;
			// PEs: 17, 17 -> 16
			// srcs: (22, 21)(465) 24, (18) 36 --> (1065) 864:NW21, ND0, *, PEGB0
			9'd21 : rdata = 43'b0001101010101011000000000000000000010000000;
			// PEs: 17, 17 -> 23
			// srcs: (23, 22)(466) 24, (18) 36 --> (1066) 864:NW22, ND0, *, PEGB7
			9'd22 : rdata = 43'b0001101010110011000000000000000000011110000;
			// PEs: 17, 17 -> 23
			// srcs: (24, 23)(467) 31, (18) 36 --> (1067) 1116:NW23, ND0, *, PEGB7
			9'd23 : rdata = 43'b0001101010111011000000000000000000011110000;
			// PEs: 17, 17 -> 17
			// srcs: (25, 24)(468) 5, (18) 36 --> (1068) 180:NW24, ND0, *, NI0
			9'd24 : rdata = 43'b0001101011000011000001000000000000000000000;
			// PEs: 17, 17 -> 17
			// srcs: (26, 25)(469) 45, (18) 36 --> (1069) 1620:NW25, ND0, *, NI1
			9'd25 : rdata = 43'b0001101011001011000001000010000000000000000;
			// PEs: 17, 17 -> 17
			// srcs: (27, 26)(470) 1, (18) 36 --> (1070) 36:NW26, ND0, *, NI2
			9'd26 : rdata = 43'b0001101011010011000001000100000000000000000;
			// PEs: 17, 17 -> 22
			// srcs: (28, 27)(471) 0, (18) 36 --> (1071) 0:NW27, ND0, *, PEGB6
			9'd27 : rdata = 43'b0001101011011011000000000000000000011100000;
			// PEs: 17, 17 -> 17
			// srcs: (29, 28)(472) -1, (18) 36 --> (1072) -36:NW28, ND0, *, NI3
			9'd28 : rdata = 43'b0001101011100011000001000110000000000000000;
			// PEs: 17, 17 -> 17
			// srcs: (30, 29)(473) -3, (18) 36 --> (1073) -108:NW29, ND0, *, NI4
			9'd29 : rdata = 43'b0001101011101011000001001000000000000000000;
			// PEs: 17, 18 -> 17
			// srcs: (31, 54)(1068) 180, (1098) -63 --> (1687) 117:NI0, PEGB2, +, NI5
			9'd30 : rdata = 43'b0000110100000111001001001010000000000000000;
			// PEs: 17, 18 -> 17
			// srcs: (32, 55)(1069) 1620, (1099) 0 --> (1706) 1620:NI1, PEGB2, +, NI0
			9'd31 : rdata = 43'b0000110100001111001001000000000000000000000;
			// PEs: 17, 18 -> 17
			// srcs: (33, 56)(1070) 36, (1100) 504 --> (1725) 540:NI2, PEGB2, +, NI1
			9'd32 : rdata = 43'b0000110100010111001001000010000000000000000;
			// PEs: 17, 18 -> 17
			// srcs: (35, 57)(1072) -36, (1102) -63 --> (1763) -99:NI3, PEGB2, +, NI2
			9'd33 : rdata = 43'b0000110100011111001001000100000000000000000;
			// PEs: 17, 18 -> 17
			// srcs: (36, 58)(1073) -108, (1103) 714 --> (1782) 606:NI4, PEGB2, +, NI3
			9'd34 : rdata = 43'b0000110100100111001001000110000000000000000;
			// PEs: 22 -> 17
			// srcs: (37, 79)(1746) 906 --> (1746) 906:PEGB6, pass, NI4
			9'd35 : rdata = 43'b1100011101100000000001001000000000000000000;
			// PEs: 19 -> 17
			// srcs: (38, 77)(1689) 199 --> (1689) 199:PEGB3, pass, NI6
			9'd36 : rdata = 43'b1100011100110000000001001100000000000000000;
			// PEs: 20, 17 -> 16
			// srcs: (39, 80)(1745) 1099, (1746) 906 --> (1751) 2005:PEGB4, NI4, +, PEGB0
			9'd37 : rdata = 43'b0000111101000101001000000000000000010000000;
			// PEs: 18, 17 -> 16
			// srcs: (41, 78)(1688) 641, (1689) 199 --> (1694) 840:PEGB2, NI6, +, PEGB0
			9'd38 : rdata = 43'b0000111100100101001100000000000000010000000;
			// PEs: 18 -> 
			// srcs: (44, 81)(1764) 283 --> (1764) 283:PEGB2, pass, 
			9'd39 : rdata = 43'b1100011100100000000000000000000000000000000;
			// PEs: 17, 22 -> 17
			// srcs: (47, 82)(1764) 283, (1765) 90 --> (1770) 373:ALU, PEGB6, +, NI4
			9'd40 : rdata = 43'b0000100111111111011001001000000000000000000;
			// PEs: 23 -> 
			// srcs: (72, 59)(1249) 96 --> (1249) 96:PEGB7, pass, 
			9'd41 : rdata = 43'b1100011101110000000000000000000000000000000;
			// PEs: 17, 23 -> 
			// srcs: (82, 60)(1249) 96, (1250) 813 --> (1256) 909:ALU, PEGB7, +, 
			9'd42 : rdata = 43'b0000100111111111011100000000000000000000000;
			// PEs: 23, 17 -> 16
			// srcs: (96, 83)(1255) 2389, (1256) 909 --> (1259) 3298:PEGB7, ALU, +, PEGB0
			9'd43 : rdata = 43'b0000111101110001111110000000000000010000000;
			// PEs: 16 -> 
			// srcs: (268, 30)(914) -19 --> (914) -19:PENB, pass, 
			9'd44 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 16, 17 -> 17
			// srcs: (274, 31)(884) 640, (914) -19 --> (1608) 621:PENB, ALU, +, NI6
			9'd45 : rdata = 43'b0000111011110001111111001100000000000000000;
			// PEs: 16 -> 
			// srcs: (277, 32)(974) 759 --> (974) 759:PENB, pass, 
			9'd46 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 16, 17 -> 17
			// srcs: (283, 33)(944) 580, (974) 759 --> (1609) 1339:PENB, ALU, +, NI7
			9'd47 : rdata = 43'b0000111011110001111111001110000000000000000;
			// PEs: 16 -> 17
			// srcs: (285, 34)(1034) 220 --> (1034) 220:PENB, pass, NI8
			9'd48 : rdata = 43'b1100011011110000000001010000000000000000000;
			// PEs: 17 -> 17
			// srcs: (286, 107)(1608) 621 --> (1608) 621:NI6, pass, NI6
			9'd49 : rdata = 43'b1100010100110000000001001100000000000000000;
			// PEs: 17, 17 -> 17
			// srcs: (286, 64)(1608) 621, (1609) 1339 --> (1616) 1960:ALU, NI7, +, NI9
			9'd50 : rdata = 43'b0000100111111101001111010010000000000000000;
			// PEs: 16, 17 -> 17
			// srcs: (291, 35)(1004) 32, (1034) 220 --> (1610) 252:PENB, NI8, +, NI6
			9'd51 : rdata = 43'b0000111011110101010001001100000000000000000;
			// PEs: 16 -> 
			// srcs: (293, 36)(915) -2 --> (915) -2:PENB, pass, 
			9'd52 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 16, 17 -> 17
			// srcs: (299, 37)(885) 128, (915) -2 --> (1627) 126:PENB, ALU, +, NI7
			9'd53 : rdata = 43'b0000111011110001111111001110000000000000000;
			// PEs: 16 -> 17
			// srcs: (301, 38)(975) 1089 --> (975) 1089:PENB, pass, NI8
			9'd54 : rdata = 43'b1100011011110000000001010000000000000000000;
			// PEs: 17, 23 -> 18
			// srcs: (304, 65)(1610) 252, (1611) 702 --> (1617) 954:NI6, PEGB7, +, PENB
			9'd55 : rdata = 43'b0000110100110111011100000000000000100000000;
			// PEs: 16, 17 -> 17
			// srcs: (307, 39)(945) 87, (975) 1089 --> (1628) 1176:PENB, NI8, +, NI6
			9'd56 : rdata = 43'b0000111011110101010001001100000000000000000;
			// PEs: 16 -> 17
			// srcs: (309, 40)(1035) 330 --> (1035) 330:PENB, pass, NI8
			9'd57 : rdata = 43'b1100011011110000000001010000000000000000000;
			// PEs: 17 -> 17
			// srcs: (310, 108)(1627) 126 --> (1627) 126:NI7, pass, NI7
			9'd58 : rdata = 43'b1100010100111000000001001110000000000000000;
			// PEs: 17, 17 -> 17
			// srcs: (310, 66)(1627) 126, (1628) 1176 --> (1635) 1302:ALU, NI6, +, NI10
			9'd59 : rdata = 43'b0000100111111101001101010100000000000000000;
			// PEs: 17 -> 18
			// srcs: (311, 84)(1616) 1960 --> (1616) 1960:NI9, pass, PENB
			9'd60 : rdata = 43'b1100010101001000000000000000000000100000000;
			// PEs: 16, 17 -> 16
			// srcs: (315, 41)(1005) 44, (1035) 330 --> (1629) 374:PENB, NI8, +, PEGB0
			9'd61 : rdata = 43'b0000111011110101010000000000000000010000000;
			// PEs: 16 -> 
			// srcs: (317, 42)(916) -23 --> (916) -23:PENB, pass, 
			9'd62 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 16, 17 -> 17
			// srcs: (323, 43)(886) 1024, (916) -23 --> (1646) 1001:PENB, ALU, +, NI6
			9'd63 : rdata = 43'b0000111011110001111111001100000000000000000;
			// PEs: 16 -> 
			// srcs: (325, 44)(976) 891 --> (976) 891:PENB, pass, 
			9'd64 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 16, 17 -> 17
			// srcs: (331, 45)(946) 1421, (976) 891 --> (1647) 2312:PENB, ALU, +, NI7
			9'd65 : rdata = 43'b0000111011110001111111001110000000000000000;
			// PEs: 16 -> 17
			// srcs: (333, 46)(1036) 0 --> (1036) 0:PENB, pass, NI8
			9'd66 : rdata = 43'b1100011011110000000001010000000000000000000;
			// PEs: 17 -> 17
			// srcs: (334, 109)(1646) 1001 --> (1646) 1001:NI6, pass, NI6
			9'd67 : rdata = 43'b1100010100110000000001001100000000000000000;
			// PEs: 17, 17 -> 17
			// srcs: (334, 67)(1646) 1001, (1647) 2312 --> (1654) 3313:ALU, NI7, +, NI9
			9'd68 : rdata = 43'b0000100111111101001111010010000000000000000;
			// PEs: 16, 17 -> 17
			// srcs: (339, 47)(1006) 70, (1036) 0 --> (1648) 70:PENB, NI8, +, NI6
			9'd69 : rdata = 43'b0000111011110101010001001100000000000000000;
			// PEs: 16 -> 
			// srcs: (341, 48)(917) -39 --> (917) -39:PENB, pass, 
			9'd70 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 16, 17 -> 17
			// srcs: (347, 49)(887) 128, (917) -39 --> (1665) 89:PENB, ALU, +, NI7
			9'd71 : rdata = 43'b0000111011110001111111001110000000000000000;
			// PEs: 16 -> 17
			// srcs: (349, 50)(977) 132 --> (977) 132:PENB, pass, NI8
			9'd72 : rdata = 43'b1100011011110000000001010000000000000000000;
			// PEs: 17, 23 -> 18
			// srcs: (352, 68)(1648) 70, (1649) 1809 --> (1655) 1879:NI6, PEGB7, +, PENB
			9'd73 : rdata = 43'b0000110100110111011100000000000000100000000;
			// PEs: 16, 17 -> 17
			// srcs: (355, 51)(947) 1015, (977) 132 --> (1666) 1147:PENB, NI8, +, NI6
			9'd74 : rdata = 43'b0000111011110101010001001100000000000000000;
			// PEs: 16 -> 17
			// srcs: (357, 52)(1037) 220 --> (1037) 220:PENB, pass, NI8
			9'd75 : rdata = 43'b1100011011110000000001010000000000000000000;
			// PEs: 17 -> 17
			// srcs: (358, 110)(1665) 89 --> (1665) 89:NI7, pass, NI7
			9'd76 : rdata = 43'b1100010100111000000001001110000000000000000;
			// PEs: 17, 17 -> 17
			// srcs: (358, 69)(1665) 89, (1666) 1147 --> (1673) 1236:ALU, NI6, +, NI11
			9'd77 : rdata = 43'b0000100111111101001101010110000000000000000;
			// PEs: 17 -> 18
			// srcs: (359, 86)(1654) 3313 --> (1654) 3313:NI9, pass, PENB
			9'd78 : rdata = 43'b1100010101001000000000000000000000100000000;
			// PEs: 16, 17 -> 17
			// srcs: (363, 53)(1007) 72, (1037) 220 --> (1667) 292:PENB, NI8, +, NI6
			9'd79 : rdata = 43'b0000111011110101010001001100000000000000000;
			// PEs: 16, 18 -> 22
			// srcs: (364, 61)(1587) 23, (1588) 780 --> (1596) 803:PENB, PEGB2, +, PEGB6
			9'd80 : rdata = 43'b0000111011110111001000000000000000011100000;
			// PEs: 18 -> 17
			// srcs: (365, 62)(1591) 732 --> (1591) 732:PEGB2, pass, NI7
			9'd81 : rdata = 43'b1100011100100000000001001110000000000000000;
			// PEs: 16, 17 -> 17
			// srcs: (366, 71)(1686) 724, (1687) 117 --> (1693) 841:PENB, NI5, +, NI8
			9'd82 : rdata = 43'b0000111011110101001011010000000000000000000;
			// PEs: 16, 17 -> 17
			// srcs: (367, 72)(1705) 358, (1706) 1620 --> (1712) 1978:PENB, NI0, +, NI5
			9'd83 : rdata = 43'b0000111011110101000001001010000000000000000;
			// PEs: 16, 17 -> 17
			// srcs: (368, 73)(1724) 482, (1725) 540 --> (1731) 1022:PENB, NI1, +, NI0
			9'd84 : rdata = 43'b0000111011110101000011000000000000000000000;
			// PEs: 16, 22 -> 16
			// srcs: (369, 74)(1743) 560, (1744) 357 --> (1750) 917:PENB, PEGB6, +, PEGB0
			9'd85 : rdata = 43'b0000111011110111011000000000000000010000000;
			// PEs: 16, 17 -> 17
			// srcs: (370, 75)(1762) 102, (1763) -99 --> (1769) 3:PENB, NI2, +, NI1
			9'd86 : rdata = 43'b0000111011110101000101000010000000000000000;
			// PEs: 16, 17 -> 17
			// srcs: (371, 76)(1781) 536, (1782) 606 --> (1788) 1142:PENB, NI3, +, NI2
			9'd87 : rdata = 43'b0000111011110101000111000100000000000000000;
			// PEs: 17, 23 -> 18
			// srcs: (374, 63)(1591) 732, (1592) 21 --> (1598) 753:NI7, PEGB7, +, PENB
			9'd88 : rdata = 43'b0000110100111111011100000000000000100000000;
			// PEs: 17, 23 -> 
			// srcs: (376, 70)(1667) 292, (1668) 1893 --> (1674) 2185:NI6, PEGB7, +, 
			9'd89 : rdata = 43'b0000110100110111011100000000000000000000000;
			// PEs: 17, 17 -> 17
			// srcs: (379, 87)(1673) 1236, (1674) 2185 --> (1677) 3421:NI11, ALU, +, NI3
			9'd90 : rdata = 43'b0000110101011001111111000110000000000000000;
			// PEs: 17, 16 -> 16
			// srcs: (513, 85)(1635) 1302, (1636) 1847 --> (1639) 3149:NI10, PENB, +, PEGB0
			9'd91 : rdata = 43'b0000110101010110111100000000000000010000000;
			// PEs: 16, 17 -> 16
			// srcs: (514, 88)(1692) 1410, (1693) 841 --> (1696) 2251:PENB, NI8, +, PEGB0
			9'd92 : rdata = 43'b0000111011110101010000000000000000010000000;
			// PEs: 16, 17 -> 16
			// srcs: (515, 89)(1711) 1614, (1712) 1978 --> (1715) 3592:PENB, NI5, +, PEGB0
			9'd93 : rdata = 43'b0000111011110101001010000000000000010000000;
			// PEs: 16, 17 -> 17
			// srcs: (1000, 90)(1730) 2549, (1731) 1022 --> (1734) 3571:PENB, NI0, +, NI5
			9'd94 : rdata = 43'b0000111011110101000001001010000000000000000;
			// PEs: 16, 17 -> 17
			// srcs: (1001, 91)(1768) 3151, (1769) 3 --> (1772) 3154:PENB, NI1, +, NI0
			9'd95 : rdata = 43'b0000111011110101000011000000000000000000000;
			// PEs: 16, 17 -> 16
			// srcs: (1002, 92)(1787) 2303, (1788) 1142 --> (1791) 3445:PENB, NI2, +, PEGB0
			9'd96 : rdata = 43'b0000111011110101000100000000000000010000000;
			// PEs: 16 -> 
			// srcs: (1004, 93)(1334) 3857 --> (1334) 3857:PENB, pass, 
			9'd97 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 16, 17 -> 16
			// srcs: (1010, 94)(1333) 532, (1334) 3857 --> (1336) 4389:PENB, ALU, +, PEGB0
			9'd98 : rdata = 43'b0000111011110001111110000000000000010000000;
			// PEs: 16 -> 
			// srcs: (1012, 95)(1524) 4683 --> (1524) 4683:PENB, pass, 
			9'd99 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 16, 17 -> 16
			// srcs: (1018, 96)(1523) 1890, (1524) 4683 --> (1526) 6573:PENB, ALU, +, PEGB0
			9'd100 : rdata = 43'b0000111011110001111110000000000000010000000;
			// PEs: 16 -> 
			// srcs: (1020, 97)(1543) 4164 --> (1543) 4164:PENB, pass, 
			9'd101 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 16, 17 -> 16
			// srcs: (1026, 98)(1542) 2466, (1543) 4164 --> (1545) 6630:PENB, ALU, +, PEGB0
			9'd102 : rdata = 43'b0000111011110001111110000000000000010000000;
			// PEs: 16 -> 
			// srcs: (1028, 99)(1581) 6146 --> (1581) 6146:PENB, pass, 
			9'd103 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 16, 17 -> 16
			// srcs: (1034, 100)(1580) 2614, (1581) 6146 --> (1583) 8760:PENB, ALU, +, PEGB0
			9'd104 : rdata = 43'b0000111011110001111110000000000000010000000;
			// PEs: 16, 22 -> 18
			// srcs: (1035, 101)(1599) 2075, (1600) 1744 --> (1602) 3819:PENB, PEGB6, +, PENB
			9'd105 : rdata = 43'b0000111011110111011000000000000000100000000;
			// PEs: 21, 16 -> 17
			// srcs: (1036, 102)(1732) 1727, (1733) 5670 --> (1735) 7397:PEGB5, PENB, +, NI1
			9'd106 : rdata = 43'b0000111101010110111101000010000000000000000;
			// PEs: 17, 16 -> 17
			// srcs: (1037, 103)(1770) 373, (1771) 6226 --> (1773) 6599:NI4, PENB, +, NI2
			9'd107 : rdata = 43'b0000110100100110111101000100000000000000000;
			// PEs: 17 -> 17
			// srcs: (1039, 111)(1734) 3571 --> (1734) 3571:NI5, pass, NI5
			9'd108 : rdata = 43'b1100010100101000000001001010000000000000000;
			// PEs: 17, 17 -> 17
			// srcs: (1039, 105)(1734) 3571, (1735) 7397 --> (1736) 10968:ALU, NI1, +, NW30
			9'd109 : rdata = 43'b0000100111111101000010000001111100000000000;
			// PEs: 17 -> 17
			// srcs: (1041, 112)(1772) 3154 --> (1772) 3154:NI0, pass, NI0
			9'd110 : rdata = 43'b1100010100000000000001000000000000000000000;
			// PEs: 17, 17 -> 17
			// srcs: (1040, 106)(1772) 3154, (1773) 6599 --> (1774) 9753:ALU, NI2, +, NW31
			9'd111 : rdata = 43'b0000100111111101000100000001111110000000000;
			// PEs: 17 -> 16
			// srcs: (1044, 104)(1677) 3421 --> (1677) 3421:NI3, pass, PEGB0
			9'd112 : rdata = 43'b1100010100011000000000000000000000010000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 18) begin
	always @(*) begin
		case(address)
			// PEs: 18, 18 -> 23
			// srcs: (1, 0)(474) 36, (19) 21 --> (1074) 756:NW0, ND0, *, PEGB7
			9'd0 : rdata = 43'b0001101000000011000000000000000000011110000;
			// PEs: 18, 18 -> 23
			// srcs: (2, 1)(475) 13, (19) 21 --> (1075) 273:NW1, ND0, *, PEGB7
			9'd1 : rdata = 43'b0001101000001011000000000000000000011110000;
			// PEs: 18, 18 -> 16
			// srcs: (3, 2)(476) 13, (19) 21 --> (1076) 273:NW2, ND0, *, PEGB0
			9'd2 : rdata = 43'b0001101000010011000000000000000000010000000;
			// PEs: 18, 18 -> 16
			// srcs: (4, 3)(477) 42, (19) 21 --> (1077) 882:NW3, ND0, *, PEGB0
			9'd3 : rdata = 43'b0001101000011011000000000000000000010000000;
			// PEs: 18, 18 -> 23
			// srcs: (5, 4)(478) 38, (19) 21 --> (1078) 798:NW4, ND0, *, PEGB7
			9'd4 : rdata = 43'b0001101000100011000000000000000000011110000;
			// PEs: 18, 18 -> 23
			// srcs: (6, 5)(479) 35, (19) 21 --> (1079) 735:NW5, ND0, *, PEGB7
			9'd5 : rdata = 43'b0001101000101011000000000000000000011110000;
			// PEs: 18, 18 -> 16
			// srcs: (7, 6)(480) 23, (19) 21 --> (1080) 483:NW6, ND0, *, PEGB0
			9'd6 : rdata = 43'b0001101000110011000000000000000000010000000;
			// PEs: 18, 18 -> 16
			// srcs: (8, 7)(481) 11, (19) 21 --> (1081) 231:NW7, ND0, *, PEGB0
			9'd7 : rdata = 43'b0001101000111011000000000000000000010000000;
			// PEs: 18, 18 -> 23
			// srcs: (9, 8)(482) 47, (19) 21 --> (1082) 987:NW8, ND0, *, PEGB7
			9'd8 : rdata = 43'b0001101001000011000000000000000000011110000;
			// PEs: 18, 18 -> 23
			// srcs: (10, 9)(483) -3, (19) 21 --> (1083) -63:NW9, ND0, *, PEGB7
			9'd9 : rdata = 43'b0001101001001011000000000000000000011110000;
			// PEs: 18, 18 -> 16
			// srcs: (11, 10)(484) 25, (19) 21 --> (1084) 525:NW10, ND0, *, PEGB0
			9'd10 : rdata = 43'b0001101001010011000000000000000000010000000;
			// PEs: 18, 18 -> 23
			// srcs: (12, 11)(485) 8, (19) 21 --> (1085) 168:NW11, ND0, *, PEGB7
			9'd11 : rdata = 43'b0001101001011011000000000000000000011110000;
			// PEs: 18, 18 -> 23
			// srcs: (13, 12)(486) -3, (19) 21 --> (1086) -63:NW12, ND0, *, PEGB7
			9'd12 : rdata = 43'b0001101001100011000000000000000000011110000;
			// PEs: 18, 18 -> 16
			// srcs: (14, 13)(487) 43, (19) 21 --> (1087) 903:NW13, ND0, *, PEGB0
			9'd13 : rdata = 43'b0001101001101011000000000000000000010000000;
			// PEs: 18, 18 -> 23
			// srcs: (15, 14)(488) 24, (19) 21 --> (1088) 504:NW14, ND0, *, PEGB7
			9'd14 : rdata = 43'b0001101001110011000000000000000000011110000;
			// PEs: 18, 18 -> 23
			// srcs: (16, 15)(489) 14, (19) 21 --> (1089) 294:NW15, ND0, *, PEGB7
			9'd15 : rdata = 43'b0001101001111011000000000000000000011110000;
			// PEs: 18, 18 -> 16
			// srcs: (17, 16)(490) 28, (19) 21 --> (1090) 588:NW16, ND0, *, PEGB0
			9'd16 : rdata = 43'b0001101010000011000000000000000000010000000;
			// PEs: 18, 18 -> 16
			// srcs: (18, 17)(491) 6, (19) 21 --> (1091) 126:NW17, ND0, *, PEGB0
			9'd17 : rdata = 43'b0001101010001011000000000000000000010000000;
			// PEs: 18, 18 -> 16
			// srcs: (19, 18)(492) 32, (19) 21 --> (1092) 672:NW18, ND0, *, PEGB0
			9'd18 : rdata = 43'b0001101010010011000000000000000000010000000;
			// PEs: 18, 18 -> 23
			// srcs: (20, 19)(493) 1, (19) 21 --> (1093) 21:NW19, ND0, *, PEGB7
			9'd19 : rdata = 43'b0001101010011011000000000000000000011110000;
			// PEs: 18, 18 -> 23
			// srcs: (21, 20)(494) 18, (19) 21 --> (1094) 378:NW20, ND0, *, PEGB7
			9'd20 : rdata = 43'b0001101010100011000000000000000000011110000;
			// PEs: 18, 18 -> 16
			// srcs: (22, 21)(495) 29, (19) 21 --> (1095) 609:NW21, ND0, *, PEGB0
			9'd21 : rdata = 43'b0001101010101011000000000000000000010000000;
			// PEs: 18, 18 -> 23
			// srcs: (23, 22)(496) 45, (19) 21 --> (1096) 945:NW22, ND0, *, PEGB7
			9'd22 : rdata = 43'b0001101010110011000000000000000000011110000;
			// PEs: 18, 18 -> 23
			// srcs: (24, 23)(497) 37, (19) 21 --> (1097) 777:NW23, ND0, *, PEGB7
			9'd23 : rdata = 43'b0001101010111011000000000000000000011110000;
			// PEs: 18, 18 -> 17
			// srcs: (25, 24)(498) -3, (19) 21 --> (1098) -63:NW24, ND0, *, PEGB1
			9'd24 : rdata = 43'b0001101011000011000000000000000000010010000;
			// PEs: 18, 18 -> 17
			// srcs: (26, 25)(499) 0, (19) 21 --> (1099) 0:NW25, ND0, *, PEGB1
			9'd25 : rdata = 43'b0001101011001011000000000000000000010010000;
			// PEs: 18, 18 -> 17
			// srcs: (27, 26)(500) 24, (19) 21 --> (1100) 504:NW26, ND0, *, PEGB1
			9'd26 : rdata = 43'b0001101011010011000000000000000000010010000;
			// PEs: 18, 18 -> 22
			// srcs: (28, 27)(501) 17, (19) 21 --> (1101) 357:NW27, ND0, *, PEGB6
			9'd27 : rdata = 43'b0001101011011011000000000000000000011100000;
			// PEs: 18, 18 -> 17
			// srcs: (29, 28)(502) -3, (19) 21 --> (1102) -63:NW28, ND0, *, PEGB1
			9'd28 : rdata = 43'b0001101011100011000000000000000000010010000;
			// PEs: 18, 18 -> 17
			// srcs: (30, 29)(503) 34, (19) 21 --> (1103) 714:NW29, ND0, *, PEGB1
			9'd29 : rdata = 43'b0001101011101011000000000000000000010010000;
			// PEs: 20 -> 18
			// srcs: (31, 38)(1158) -26 --> (1158) -26:PEGB4, pass, NI0
			9'd30 : rdata = 43'b1100011101000000000001000000000000000000000;
			// PEs: 20 -> 18
			// srcs: (32, 40)(1159) 637 --> (1159) 637:PEGB4, pass, NI1
			9'd31 : rdata = 43'b1100011101000000000001000010000000000000000;
			// PEs: 19, 18 -> 17
			// srcs: (33, 39)(1128) 667, (1158) -26 --> (1688) 641:PEGB3, NI0, +, PEGB1
			9'd32 : rdata = 43'b0000111100110101000000000000000000010010000;
			// PEs: 20 -> 18
			// srcs: (34, 42)(1162) -39 --> (1162) -39:PEGB4, pass, NI0
			9'd33 : rdata = 43'b1100011101000000000001000000000000000000000;
			// PEs: 19, 18 -> 19
			// srcs: (36, 41)(1129) 276, (1159) 637 --> (1707) 913:PEGB3, NI1, +, PENB
			9'd34 : rdata = 43'b0000111100110101000010000000000000100000000;
			// PEs: 19, 18 -> 17
			// srcs: (39, 43)(1132) 322, (1162) -39 --> (1764) 283:PEGB3, NI0, +, PEGB1
			9'd35 : rdata = 43'b0000111100110101000000000000000000010010000;
			// PEs: 16 -> 
			// srcs: (236, 30)(853) 160 --> (853) 160:PEGB0, pass, 
			9'd36 : rdata = 43'b1100011100000000000000000000000000000000000;
			// PEs: 16, 18 -> 17
			// srcs: (245, 31)(823) 620, (853) 160 --> (1588) 780:PEGB0, ALU, +, PEGB1
			9'd37 : rdata = 43'b0000111100000001111110000000000000010010000;
			// PEs: 16 -> 
			// srcs: (247, 32)(913) -30 --> (913) -30:PEGB0, pass, 
			9'd38 : rdata = 43'b1100011100000000000000000000000000000000000;
			// PEs: 16, 18 -> 18
			// srcs: (256, 33)(883) -96, (913) -30 --> (1589) -126:PEGB0, ALU, +, NI0
			9'd39 : rdata = 43'b0000111100000001111111000000000000000000000;
			// PEs: 16 -> 
			// srcs: (258, 34)(973) 363 --> (973) 363:PEGB0, pass, 
			9'd40 : rdata = 43'b1100011100000000000000000000000000000000000;
			// PEs: 16, 18 -> 18
			// srcs: (267, 35)(943) 203, (973) 363 --> (1590) 566:PEGB0, ALU, +, NI1
			9'd41 : rdata = 43'b0000111100000001111111000010000000000000000;
			// PEs: 16 -> 18
			// srcs: (269, 36)(1033) 638 --> (1033) 638:PEGB0, pass, NI2
			9'd42 : rdata = 43'b1100011100000000000001000100000000000000000;
			// PEs: 18 -> 18
			// srcs: (270, 51)(1589) -126 --> (1589) -126:NI0, pass, NI0
			9'd43 : rdata = 43'b1100010100000000000001000000000000000000000;
			// PEs: 18, 18 -> 18
			// srcs: (270, 44)(1589) -126, (1590) 566 --> (1597) 440:ALU, NI1, +, NI3
			9'd44 : rdata = 43'b0000100111111101000011000110000000000000000;
			// PEs: 16, 18 -> 17
			// srcs: (278, 37)(1003) 94, (1033) 638 --> (1591) 732:PEGB0, NI2, +, PEGB1
			9'd45 : rdata = 43'b0000111100000101000100000000000000010010000;
			// PEs: 17 -> 
			// srcs: (306, 46)(1617) 954 --> (1617) 954:PENB, pass, 
			9'd46 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 17, 18 -> 16
			// srcs: (313, 47)(1616) 1960, (1617) 954 --> (1620) 2914:PENB, ALU, +, PEGB0
			9'd47 : rdata = 43'b0000111011110001111110000000000000010000000;
			// PEs: 17 -> 
			// srcs: (354, 48)(1655) 1879 --> (1655) 1879:PENB, pass, 
			9'd48 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 17, 18 -> 16
			// srcs: (361, 49)(1654) 3313, (1655) 1879 --> (1658) 5192:PENB, ALU, +, PEGB0
			9'd49 : rdata = 43'b0000111011110001111110000000000000010000000;
			// PEs: 18, 17 -> 
			// srcs: (377, 45)(1597) 440, (1598) 753 --> (1601) 1193:NI3, PENB, +, 
			9'd50 : rdata = 43'b0000110100011110111100000000000000000000000;
			// PEs: 18, 17 -> 18
			// srcs: (1038, 50)(1601) 1193, (1602) 3819 --> (1603) 5012:ALU, PENB, +, NW30
			9'd51 : rdata = 43'b0000100111111110111100000001111100000000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 19) begin
	always @(*) begin
		case(address)
			// PEs: 19, 19 -> 23
			// srcs: (1, 0)(504) 21, (20) 23 --> (1104) 483:NW0, ND0, *, PEGB7
			9'd0 : rdata = 43'b0001101000000011000000000000000000011110000;
			// PEs: 19, 19 -> 16
			// srcs: (2, 1)(505) 39, (20) 23 --> (1105) 897:NW1, ND0, *, PEGB0
			9'd1 : rdata = 43'b0001101000001011000000000000000000010000000;
			// PEs: 19, 19 -> 16
			// srcs: (3, 2)(506) 19, (20) 23 --> (1106) 437:NW2, ND0, *, PEGB0
			9'd2 : rdata = 43'b0001101000010011000000000000000000010000000;
			// PEs: 19, 19 -> 16
			// srcs: (4, 3)(507) 35, (20) 23 --> (1107) 805:NW3, ND0, *, PEGB0
			9'd3 : rdata = 43'b0001101000011011000000000000000000010000000;
			// PEs: 19, 19 -> 16
			// srcs: (5, 4)(508) 46, (20) 23 --> (1108) 1058:NW4, ND0, *, PEGB0
			9'd4 : rdata = 43'b0001101000100011000000000000000000010000000;
			// PEs: 19, 19 -> 16
			// srcs: (6, 5)(509) 2, (20) 23 --> (1109) 46:NW5, ND0, *, PEGB0
			9'd5 : rdata = 43'b0001101000101011000000000000000000010000000;
			// PEs: 19, 19 -> 16
			// srcs: (7, 6)(510) 17, (20) 23 --> (1110) 391:NW6, ND0, *, PEGB0
			9'd6 : rdata = 43'b0001101000110011000000000000000000010000000;
			// PEs: 19, 19 -> 16
			// srcs: (8, 7)(511) 19, (20) 23 --> (1111) 437:NW7, ND0, *, PEGB0
			9'd7 : rdata = 43'b0001101000111011000000000000000000010000000;
			// PEs: 19, 19 -> 16
			// srcs: (9, 8)(512) 7, (20) 23 --> (1112) 161:NW8, ND0, *, PEGB0
			9'd8 : rdata = 43'b0001101001000011000000000000000000010000000;
			// PEs: 19, 19 -> 16
			// srcs: (10, 9)(513) 13, (20) 23 --> (1113) 299:NW9, ND0, *, PEGB0
			9'd9 : rdata = 43'b0001101001001011000000000000000000010000000;
			// PEs: 19, 19 -> 16
			// srcs: (11, 10)(514) 21, (20) 23 --> (1114) 483:NW10, ND0, *, PEGB0
			9'd10 : rdata = 43'b0001101001010011000000000000000000010000000;
			// PEs: 19, 19 -> 16
			// srcs: (12, 11)(515) 3, (20) 23 --> (1115) 69:NW11, ND0, *, PEGB0
			9'd11 : rdata = 43'b0001101001011011000000000000000000010000000;
			// PEs: 19, 19 -> 16
			// srcs: (13, 12)(516) 26, (20) 23 --> (1116) 598:NW12, ND0, *, PEGB0
			9'd12 : rdata = 43'b0001101001100011000000000000000000010000000;
			// PEs: 19, 19 -> 16
			// srcs: (14, 13)(517) 45, (20) 23 --> (1117) 1035:NW13, ND0, *, PEGB0
			9'd13 : rdata = 43'b0001101001101011000000000000000000010000000;
			// PEs: 19, 19 -> 16
			// srcs: (15, 14)(518) 17, (20) 23 --> (1118) 391:NW14, ND0, *, PEGB0
			9'd14 : rdata = 43'b0001101001110011000000000000000000010000000;
			// PEs: 19, 19 -> 16
			// srcs: (16, 15)(519) 14, (20) 23 --> (1119) 322:NW15, ND0, *, PEGB0
			9'd15 : rdata = 43'b0001101001111011000000000000000000010000000;
			// PEs: 19, 19 -> 16
			// srcs: (17, 16)(520) 19, (20) 23 --> (1120) 437:NW16, ND0, *, PEGB0
			9'd16 : rdata = 43'b0001101010000011000000000000000000010000000;
			// PEs: 19, 19 -> 16
			// srcs: (18, 17)(521) 42, (20) 23 --> (1121) 966:NW17, ND0, *, PEGB0
			9'd17 : rdata = 43'b0001101010001011000000000000000000010000000;
			// PEs: 19, 19 -> 16
			// srcs: (19, 18)(522) 40, (20) 23 --> (1122) 920:NW18, ND0, *, PEGB0
			9'd18 : rdata = 43'b0001101010010011000000000000000000010000000;
			// PEs: 19, 19 -> 16
			// srcs: (20, 19)(523) 37, (20) 23 --> (1123) 851:NW19, ND0, *, PEGB0
			9'd19 : rdata = 43'b0001101010011011000000000000000000010000000;
			// PEs: 19, 19 -> 16
			// srcs: (21, 20)(524) 49, (20) 23 --> (1124) 1127:NW20, ND0, *, PEGB0
			9'd20 : rdata = 43'b0001101010100011000000000000000000010000000;
			// PEs: 19, 19 -> 16
			// srcs: (22, 21)(525) 6, (20) 23 --> (1125) 138:NW21, ND0, *, PEGB0
			9'd21 : rdata = 43'b0001101010101011000000000000000000010000000;
			// PEs: 19, 19 -> 16
			// srcs: (23, 22)(526) 39, (20) 23 --> (1126) 897:NW22, ND0, *, PEGB0
			9'd22 : rdata = 43'b0001101010110011000000000000000000010000000;
			// PEs: 19, 19 -> 16
			// srcs: (24, 23)(527) 43, (20) 23 --> (1127) 989:NW23, ND0, *, PEGB0
			9'd23 : rdata = 43'b0001101010111011000000000000000000010000000;
			// PEs: 19, 19 -> 18
			// srcs: (25, 24)(528) 29, (20) 23 --> (1128) 667:NW24, ND0, *, PEGB2
			9'd24 : rdata = 43'b0001101011000011000000000000000000010100000;
			// PEs: 19, 19 -> 18
			// srcs: (26, 25)(529) 12, (20) 23 --> (1129) 276:NW25, ND0, *, PEGB2
			9'd25 : rdata = 43'b0001101011001011000000000000000000010100000;
			// PEs: 19, 19 -> 21
			// srcs: (27, 26)(530) -3, (20) 23 --> (1130) -69:NW26, ND0, *, PEGB5
			9'd26 : rdata = 43'b0001101011010011000000000000000000011010000;
			// PEs: 19, 19 -> 20
			// srcs: (28, 27)(531) 28, (20) 23 --> (1131) 644:NW27, ND0, *, PENB
			9'd27 : rdata = 43'b0001101011011011000000000000000000100000000;
			// PEs: 19, 19 -> 18
			// srcs: (29, 28)(532) 14, (20) 23 --> (1132) 322:NW28, ND0, *, PEGB2
			9'd28 : rdata = 43'b0001101011100011000000000000000000010100000;
			// PEs: 19, 19 -> 20
			// srcs: (30, 29)(533) 11, (20) 23 --> (1133) 253:NW29, ND0, *, PENB
			9'd29 : rdata = 43'b0001101011101011000000000000000000100000000;
			// PEs: 22 -> 19
			// srcs: (31, 30)(1218) 217 --> (1218) 217:PEGB6, pass, NI0
			9'd30 : rdata = 43'b1100011101100000000001000000000000000000000;
			// PEs: 22 -> 19
			// srcs: (32, 32)(1219) 837 --> (1219) 837:PEGB6, pass, NI1
			9'd31 : rdata = 43'b1100011101100000000001000010000000000000000;
			// PEs: 21, 19 -> 17
			// srcs: (33, 31)(1188) -18, (1218) 217 --> (1689) 199:PEGB5, NI0, +, PEGB1
			9'd32 : rdata = 43'b0000111101010101000000000000000000010010000;
			// PEs: 21, 19 -> 
			// srcs: (36, 33)(1189) 423, (1219) 837 --> (1708) 1260:PEGB5, NI1, +, 
			9'd33 : rdata = 43'b0000111101010101000010000000000000000000000;
			// PEs: 18, 19 -> 16
			// srcs: (39, 34)(1707) 913, (1708) 1260 --> (1713) 2173:PENB, ALU, +, PEGB0
			9'd34 : rdata = 43'b0000111011110001111110000000000000010000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 20) begin
	always @(*) begin
		case(address)
			// PEs: 20, 20 -> 23
			// srcs: (1, 0)(534) 10, (21) 13 --> (1134) 130:NW0, ND0, *, PEGB7
			9'd0 : rdata = 43'b0001101000000011000000000000000000011110000;
			// PEs: 20, 20 -> 16
			// srcs: (2, 1)(535) -3, (21) 13 --> (1135) -39:NW1, ND0, *, PEGB0
			9'd1 : rdata = 43'b0001101000001011000000000000000000010000000;
			// PEs: 20, 20 -> 16
			// srcs: (3, 2)(536) 36, (21) 13 --> (1136) 468:NW2, ND0, *, PEGB0
			9'd2 : rdata = 43'b0001101000010011000000000000000000010000000;
			// PEs: 20, 20 -> 16
			// srcs: (4, 3)(537) 46, (21) 13 --> (1137) 598:NW3, ND0, *, PEGB0
			9'd3 : rdata = 43'b0001101000011011000000000000000000010000000;
			// PEs: 20, 20 -> 16
			// srcs: (5, 4)(538) 33, (21) 13 --> (1138) 429:NW4, ND0, *, PEGB0
			9'd4 : rdata = 43'b0001101000100011000000000000000000010000000;
			// PEs: 20, 20 -> 16
			// srcs: (6, 5)(539) 11, (21) 13 --> (1139) 143:NW5, ND0, *, PEGB0
			9'd5 : rdata = 43'b0001101000101011000000000000000000010000000;
			// PEs: 20, 20 -> 16
			// srcs: (7, 6)(540) 3, (21) 13 --> (1140) 39:NW6, ND0, *, PEGB0
			9'd6 : rdata = 43'b0001101000110011000000000000000000010000000;
			// PEs: 20, 20 -> 16
			// srcs: (8, 7)(541) 7, (21) 13 --> (1141) 91:NW7, ND0, *, PEGB0
			9'd7 : rdata = 43'b0001101000111011000000000000000000010000000;
			// PEs: 20, 20 -> 16
			// srcs: (9, 8)(542) 7, (21) 13 --> (1142) 91:NW8, ND0, *, PEGB0
			9'd8 : rdata = 43'b0001101001000011000000000000000000010000000;
			// PEs: 20, 20 -> 16
			// srcs: (10, 9)(543) 30, (21) 13 --> (1143) 390:NW9, ND0, *, PEGB0
			9'd9 : rdata = 43'b0001101001001011000000000000000000010000000;
			// PEs: 20, 20 -> 16
			// srcs: (11, 10)(544) 1, (21) 13 --> (1144) 13:NW10, ND0, *, PEGB0
			9'd10 : rdata = 43'b0001101001010011000000000000000000010000000;
			// PEs: 20, 20 -> 16
			// srcs: (12, 11)(545) 24, (21) 13 --> (1145) 312:NW11, ND0, *, PEGB0
			9'd11 : rdata = 43'b0001101001011011000000000000000000010000000;
			// PEs: 20, 20 -> 16
			// srcs: (13, 12)(546) 15, (21) 13 --> (1146) 195:NW12, ND0, *, PEGB0
			9'd12 : rdata = 43'b0001101001100011000000000000000000010000000;
			// PEs: 20, 20 -> 16
			// srcs: (14, 13)(547) 29, (21) 13 --> (1147) 377:NW13, ND0, *, PEGB0
			9'd13 : rdata = 43'b0001101001101011000000000000000000010000000;
			// PEs: 20, 20 -> 16
			// srcs: (15, 14)(548) 21, (21) 13 --> (1148) 273:NW14, ND0, *, PEGB0
			9'd14 : rdata = 43'b0001101001110011000000000000000000010000000;
			// PEs: 20, 20 -> 16
			// srcs: (16, 15)(549) 33, (21) 13 --> (1149) 429:NW15, ND0, *, PEGB0
			9'd15 : rdata = 43'b0001101001111011000000000000000000010000000;
			// PEs: 20, 20 -> 16
			// srcs: (17, 16)(550) 43, (21) 13 --> (1150) 559:NW16, ND0, *, PEGB0
			9'd16 : rdata = 43'b0001101010000011000000000000000000010000000;
			// PEs: 20, 20 -> 16
			// srcs: (18, 17)(551) 41, (21) 13 --> (1151) 533:NW17, ND0, *, PEGB0
			9'd17 : rdata = 43'b0001101010001011000000000000000000010000000;
			// PEs: 20, 20 -> 16
			// srcs: (19, 18)(552) 24, (21) 13 --> (1152) 312:NW18, ND0, *, PEGB0
			9'd18 : rdata = 43'b0001101010010011000000000000000000010000000;
			// PEs: 20, 20 -> 16
			// srcs: (20, 19)(553) 29, (21) 13 --> (1153) 377:NW19, ND0, *, PEGB0
			9'd19 : rdata = 43'b0001101010011011000000000000000000010000000;
			// PEs: 20, 20 -> 16
			// srcs: (21, 20)(554) 21, (21) 13 --> (1154) 273:NW20, ND0, *, PEGB0
			9'd20 : rdata = 43'b0001101010100011000000000000000000010000000;
			// PEs: 20, 20 -> 16
			// srcs: (22, 21)(555) 0, (21) 13 --> (1155) 0:NW21, ND0, *, PEGB0
			9'd21 : rdata = 43'b0001101010101011000000000000000000010000000;
			// PEs: 20, 20 -> 16
			// srcs: (23, 22)(556) 3, (21) 13 --> (1156) 39:NW22, ND0, *, PEGB0
			9'd22 : rdata = 43'b0001101010110011000000000000000000010000000;
			// PEs: 20, 20 -> 16
			// srcs: (24, 23)(557) 15, (21) 13 --> (1157) 195:NW23, ND0, *, PEGB0
			9'd23 : rdata = 43'b0001101010111011000000000000000000010000000;
			// PEs: 20, 20 -> 18
			// srcs: (25, 24)(558) -2, (21) 13 --> (1158) -26:NW24, ND0, *, PEGB2
			9'd24 : rdata = 43'b0001101011000011000000000000000000010100000;
			// PEs: 20, 20 -> 18
			// srcs: (26, 25)(559) 49, (21) 13 --> (1159) 637:NW25, ND0, *, PEGB2
			9'd25 : rdata = 43'b0001101011001011000000000000000000010100000;
			// PEs: 20, 20 -> 21
			// srcs: (27, 26)(560) 44, (21) 13 --> (1160) 572:NW26, ND0, *, PENB
			9'd26 : rdata = 43'b0001101011010011000000000000000000100000000;
			// PEs: 20, 20 -> 20
			// srcs: (28, 27)(561) 35, (21) 13 --> (1161) 455:NW27, ND0, *, NI0
			9'd27 : rdata = 43'b0001101011011011000001000000000000000000000;
			// PEs: 20, 20 -> 18
			// srcs: (29, 28)(562) -3, (21) 13 --> (1162) -39:NW28, ND0, *, PEGB2
			9'd28 : rdata = 43'b0001101011100011000000000000000000010100000;
			// PEs: 20, 20 -> 20
			// srcs: (30, 29)(563) 33, (21) 13 --> (1163) 429:NW29, ND0, *, NI1
			9'd29 : rdata = 43'b0001101011101011000001000010000000000000000;
			// PEs: 19, 20 -> 17
			// srcs: (31, 32)(1131) 644, (1161) 455 --> (1745) 1099:PENB, NI0, +, PEGB1
			9'd30 : rdata = 43'b0000111011110101000000000000000000010010000;
			// PEs: 22 -> 20
			// srcs: (32, 30)(1220) 1116 --> (1220) 1116:PEGB6, pass, NI0
			9'd31 : rdata = 43'b1100011101100000000001000000000000000000000;
			// PEs: 19, 20 -> 20
			// srcs: (33, 33)(1133) 253, (1163) 429 --> (1783) 682:PENB, NI1, +, NI2
			9'd32 : rdata = 43'b0000111011110101000011000100000000000000000;
			// PEs: 21, 20 -> 21
			// srcs: (35, 31)(1190) 108, (1220) 1116 --> (1727) 1224:PEGB5, NI0, +, PENB
			9'd33 : rdata = 43'b0000111101010101000000000000000000100000000;
			// PEs: 22 -> 
			// srcs: (36, 34)(1223) 1147 --> (1223) 1147:PEGB6, pass, 
			9'd34 : rdata = 43'b1100011101100000000000000000000000000000000;
			// PEs: 21, 20 -> 
			// srcs: (38, 35)(1193) 288, (1223) 1147 --> (1784) 1435:PEGB5, ALU, +, 
			9'd35 : rdata = 43'b0000111101010001111110000000000000000000000;
			// PEs: 20, 20 -> 16
			// srcs: (41, 36)(1783) 682, (1784) 1435 --> (1789) 2117:NI2, ALU, +, PEGB0
			9'd36 : rdata = 43'b0000110100010001111110000000000000010000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 21) begin
	always @(*) begin
		case(address)
			// PEs: 21, 21 -> 16
			// srcs: (1, 0)(564) -1, (22) 9 --> (1164) -9:NW0, ND0, *, PEGB0
			9'd0 : rdata = 43'b0001101000000011000000000000000000010000000;
			// PEs: 21, 21 -> 16
			// srcs: (2, 1)(565) 13, (22) 9 --> (1165) 117:NW1, ND0, *, PEGB0
			9'd1 : rdata = 43'b0001101000001011000000000000000000010000000;
			// PEs: 21, 21 -> 16
			// srcs: (3, 2)(566) 18, (22) 9 --> (1166) 162:NW2, ND0, *, PEGB0
			9'd2 : rdata = 43'b0001101000010011000000000000000000010000000;
			// PEs: 21, 21 -> 16
			// srcs: (4, 3)(567) 18, (22) 9 --> (1167) 162:NW3, ND0, *, PEGB0
			9'd3 : rdata = 43'b0001101000011011000000000000000000010000000;
			// PEs: 21, 21 -> 16
			// srcs: (5, 4)(568) 5, (22) 9 --> (1168) 45:NW4, ND0, *, PEGB0
			9'd4 : rdata = 43'b0001101000100011000000000000000000010000000;
			// PEs: 21, 21 -> 16
			// srcs: (6, 5)(569) 45, (22) 9 --> (1169) 405:NW5, ND0, *, PEGB0
			9'd5 : rdata = 43'b0001101000101011000000000000000000010000000;
			// PEs: 21, 21 -> 16
			// srcs: (7, 6)(570) -1, (22) 9 --> (1170) -9:NW6, ND0, *, PEGB0
			9'd6 : rdata = 43'b0001101000110011000000000000000000010000000;
			// PEs: 21, 21 -> 16
			// srcs: (8, 7)(571) 41, (22) 9 --> (1171) 369:NW7, ND0, *, PEGB0
			9'd7 : rdata = 43'b0001101000111011000000000000000000010000000;
			// PEs: 21, 21 -> 16
			// srcs: (9, 8)(572) 41, (22) 9 --> (1172) 369:NW8, ND0, *, PEGB0
			9'd8 : rdata = 43'b0001101001000011000000000000000000010000000;
			// PEs: 21, 21 -> 16
			// srcs: (10, 9)(573) 4, (22) 9 --> (1173) 36:NW9, ND0, *, PEGB0
			9'd9 : rdata = 43'b0001101001001011000000000000000000010000000;
			// PEs: 21, 21 -> 16
			// srcs: (11, 10)(574) 18, (22) 9 --> (1174) 162:NW10, ND0, *, PEGB0
			9'd10 : rdata = 43'b0001101001010011000000000000000000010000000;
			// PEs: 21, 21 -> 16
			// srcs: (12, 11)(575) 22, (22) 9 --> (1175) 198:NW11, ND0, *, PEGB0
			9'd11 : rdata = 43'b0001101001011011000000000000000000010000000;
			// PEs: 21, 21 -> 16
			// srcs: (13, 12)(576) 40, (22) 9 --> (1176) 360:NW12, ND0, *, PEGB0
			9'd12 : rdata = 43'b0001101001100011000000000000000000010000000;
			// PEs: 21, 21 -> 16
			// srcs: (14, 13)(577) 44, (22) 9 --> (1177) 396:NW13, ND0, *, PEGB0
			9'd13 : rdata = 43'b0001101001101011000000000000000000010000000;
			// PEs: 21, 21 -> 16
			// srcs: (15, 14)(578) 9, (22) 9 --> (1178) 81:NW14, ND0, *, PEGB0
			9'd14 : rdata = 43'b0001101001110011000000000000000000010000000;
			// PEs: 21, 21 -> 16
			// srcs: (16, 15)(579) 37, (22) 9 --> (1179) 333:NW15, ND0, *, PEGB0
			9'd15 : rdata = 43'b0001101001111011000000000000000000010000000;
			// PEs: 21, 21 -> 16
			// srcs: (17, 16)(580) 29, (22) 9 --> (1180) 261:NW16, ND0, *, PEGB0
			9'd16 : rdata = 43'b0001101010000011000000000000000000010000000;
			// PEs: 21, 21 -> 16
			// srcs: (18, 17)(581) 42, (22) 9 --> (1181) 378:NW17, ND0, *, PEGB0
			9'd17 : rdata = 43'b0001101010001011000000000000000000010000000;
			// PEs: 21, 21 -> 16
			// srcs: (19, 18)(582) 33, (22) 9 --> (1182) 297:NW18, ND0, *, PEGB0
			9'd18 : rdata = 43'b0001101010010011000000000000000000010000000;
			// PEs: 21, 21 -> 16
			// srcs: (20, 19)(583) 8, (22) 9 --> (1183) 72:NW19, ND0, *, PEGB0
			9'd19 : rdata = 43'b0001101010011011000000000000000000010000000;
			// PEs: 21, 21 -> 16
			// srcs: (21, 20)(584) 9, (22) 9 --> (1184) 81:NW20, ND0, *, PEGB0
			9'd20 : rdata = 43'b0001101010100011000000000000000000010000000;
			// PEs: 21, 21 -> 16
			// srcs: (22, 21)(585) 16, (22) 9 --> (1185) 144:NW21, ND0, *, PEGB0
			9'd21 : rdata = 43'b0001101010101011000000000000000000010000000;
			// PEs: 21, 21 -> 16
			// srcs: (23, 22)(586) 22, (22) 9 --> (1186) 198:NW22, ND0, *, PEGB0
			9'd22 : rdata = 43'b0001101010110011000000000000000000010000000;
			// PEs: 21, 21 -> 16
			// srcs: (24, 23)(587) 49, (22) 9 --> (1187) 441:NW23, ND0, *, PEGB0
			9'd23 : rdata = 43'b0001101010111011000000000000000000010000000;
			// PEs: 21, 21 -> 19
			// srcs: (25, 24)(588) -2, (22) 9 --> (1188) -18:NW24, ND0, *, PEGB3
			9'd24 : rdata = 43'b0001101011000011000000000000000000010110000;
			// PEs: 21, 21 -> 19
			// srcs: (26, 25)(589) 47, (22) 9 --> (1189) 423:NW25, ND0, *, PEGB3
			9'd25 : rdata = 43'b0001101011001011000000000000000000010110000;
			// PEs: 21, 21 -> 20
			// srcs: (27, 26)(590) 12, (22) 9 --> (1190) 108:NW26, ND0, *, PEGB4
			9'd26 : rdata = 43'b0001101011010011000000000000000000011000000;
			// PEs: 21, 21 -> 22
			// srcs: (28, 27)(591) 49, (22) 9 --> (1191) 441:NW27, ND0, *, PENB
			9'd27 : rdata = 43'b0001101011011011000000000000000000100000000;
			// PEs: 21, 21 -> 22
			// srcs: (29, 28)(592) 10, (22) 9 --> (1192) 90:NW28, ND0, *, PENB
			9'd28 : rdata = 43'b0001101011100011000000000000000000100000000;
			// PEs: 21, 21 -> 20
			// srcs: (30, 29)(593) 32, (22) 9 --> (1193) 288:NW29, ND0, *, PEGB4
			9'd29 : rdata = 43'b0001101011101011000000000000000000011000000;
			// PEs: 19, 20 -> 
			// srcs: (33, 30)(1130) -69, (1160) 572 --> (1726) 503:PEGB3, PENB, +, 
			9'd30 : rdata = 43'b0000111100110110111100000000000000000000000;
			// PEs: 21, 20 -> 17
			// srcs: (38, 31)(1726) 503, (1727) 1224 --> (1732) 1727:ALU, PENB, +, PEGB1
			9'd31 : rdata = 43'b0000100111111110111100000000000000010010000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 22) begin
	always @(*) begin
		case(address)
			// PEs: 22, 22 -> 16
			// srcs: (1, 0)(594) 11, (23) 31 --> (1194) 341:NW0, ND0, *, PEGB0
			9'd0 : rdata = 43'b0001101000000011000000000000000000010000000;
			// PEs: 22, 22 -> 16
			// srcs: (2, 1)(595) 3, (23) 31 --> (1195) 93:NW1, ND0, *, PEGB0
			9'd1 : rdata = 43'b0001101000001011000000000000000000010000000;
			// PEs: 22, 22 -> 16
			// srcs: (3, 2)(596) 40, (23) 31 --> (1196) 1240:NW2, ND0, *, PEGB0
			9'd2 : rdata = 43'b0001101000010011000000000000000000010000000;
			// PEs: 22, 22 -> 16
			// srcs: (4, 3)(597) 32, (23) 31 --> (1197) 992:NW3, ND0, *, PEGB0
			9'd3 : rdata = 43'b0001101000011011000000000000000000010000000;
			// PEs: 22, 22 -> 16
			// srcs: (5, 4)(598) 48, (23) 31 --> (1198) 1488:NW4, ND0, *, PEGB0
			9'd4 : rdata = 43'b0001101000100011000000000000000000010000000;
			// PEs: 22, 22 -> 16
			// srcs: (6, 5)(599) -2, (23) 31 --> (1199) -62:NW5, ND0, *, PEGB0
			9'd5 : rdata = 43'b0001101000101011000000000000000000010000000;
			// PEs: 22, 22 -> 16
			// srcs: (7, 6)(600) 14, (23) 31 --> (1200) 434:NW6, ND0, *, PEGB0
			9'd6 : rdata = 43'b0001101000110011000000000000000000010000000;
			// PEs: 22, 22 -> 16
			// srcs: (8, 7)(601) 6, (23) 31 --> (1201) 186:NW7, ND0, *, PEGB0
			9'd7 : rdata = 43'b0001101000111011000000000000000000010000000;
			// PEs: 22, 22 -> 16
			// srcs: (9, 8)(602) 43, (23) 31 --> (1202) 1333:NW8, ND0, *, PEGB0
			9'd8 : rdata = 43'b0001101001000011000000000000000000010000000;
			// PEs: 22, 22 -> 16
			// srcs: (10, 9)(603) 17, (23) 31 --> (1203) 527:NW9, ND0, *, PEGB0
			9'd9 : rdata = 43'b0001101001001011000000000000000000010000000;
			// PEs: 22, 22 -> 16
			// srcs: (11, 10)(604) 42, (23) 31 --> (1204) 1302:NW10, ND0, *, PEGB0
			9'd10 : rdata = 43'b0001101001010011000000000000000000010000000;
			// PEs: 22, 22 -> 16
			// srcs: (12, 11)(605) 1, (23) 31 --> (1205) 31:NW11, ND0, *, PEGB0
			9'd11 : rdata = 43'b0001101001011011000000000000000000010000000;
			// PEs: 22, 22 -> 16
			// srcs: (13, 12)(606) 38, (23) 31 --> (1206) 1178:NW12, ND0, *, PEGB0
			9'd12 : rdata = 43'b0001101001100011000000000000000000010000000;
			// PEs: 22, 22 -> 16
			// srcs: (14, 13)(607) 12, (23) 31 --> (1207) 372:NW13, ND0, *, PEGB0
			9'd13 : rdata = 43'b0001101001101011000000000000000000010000000;
			// PEs: 22, 22 -> 16
			// srcs: (15, 14)(608) -2, (23) 31 --> (1208) -62:NW14, ND0, *, PEGB0
			9'd14 : rdata = 43'b0001101001110011000000000000000000010000000;
			// PEs: 22, 22 -> 16
			// srcs: (16, 15)(609) 26, (23) 31 --> (1209) 806:NW15, ND0, *, PEGB0
			9'd15 : rdata = 43'b0001101001111011000000000000000000010000000;
			// PEs: 22, 22 -> 16
			// srcs: (17, 16)(610) 39, (23) 31 --> (1210) 1209:NW16, ND0, *, PEGB0
			9'd16 : rdata = 43'b0001101010000011000000000000000000010000000;
			// PEs: 22, 22 -> 16
			// srcs: (18, 17)(611) 43, (23) 31 --> (1211) 1333:NW17, ND0, *, PEGB0
			9'd17 : rdata = 43'b0001101010001011000000000000000000010000000;
			// PEs: 22, 22 -> 16
			// srcs: (19, 18)(612) 35, (23) 31 --> (1212) 1085:NW18, ND0, *, PEGB0
			9'd18 : rdata = 43'b0001101010010011000000000000000000010000000;
			// PEs: 22, 22 -> 16
			// srcs: (20, 19)(613) 25, (23) 31 --> (1213) 775:NW19, ND0, *, PEGB0
			9'd19 : rdata = 43'b0001101010011011000000000000000000010000000;
			// PEs: 22, 22 -> 16
			// srcs: (21, 20)(614) -1, (23) 31 --> (1214) -31:NW20, ND0, *, PEGB0
			9'd20 : rdata = 43'b0001101010100011000000000000000000010000000;
			// PEs: 22, 22 -> 16
			// srcs: (22, 21)(615) -3, (23) 31 --> (1215) -93:NW21, ND0, *, PEGB0
			9'd21 : rdata = 43'b0001101010101011000000000000000000010000000;
			// PEs: 22, 22 -> 16
			// srcs: (23, 22)(616) 11, (23) 31 --> (1216) 341:NW22, ND0, *, PEGB0
			9'd22 : rdata = 43'b0001101010110011000000000000000000010000000;
			// PEs: 22, 22 -> 16
			// srcs: (24, 23)(617) 10, (23) 31 --> (1217) 310:NW23, ND0, *, PEGB0
			9'd23 : rdata = 43'b0001101010111011000000000000000000010000000;
			// PEs: 22, 22 -> 19
			// srcs: (25, 24)(618) 7, (23) 31 --> (1218) 217:NW24, ND0, *, PEGB3
			9'd24 : rdata = 43'b0001101011000011000000000000000000010110000;
			// PEs: 22, 22 -> 19
			// srcs: (26, 25)(619) 27, (23) 31 --> (1219) 837:NW25, ND0, *, PEGB3
			9'd25 : rdata = 43'b0001101011001011000000000000000000010110000;
			// PEs: 22, 22 -> 20
			// srcs: (27, 26)(620) 36, (23) 31 --> (1220) 1116:NW26, ND0, *, PEGB4
			9'd26 : rdata = 43'b0001101011010011000000000000000000011000000;
			// PEs: 22, 22 -> 22
			// srcs: (28, 27)(621) 15, (23) 31 --> (1221) 465:NW27, ND0, *, NI0
			9'd27 : rdata = 43'b0001101011011011000001000000000000000000000;
			// PEs: 22, 22 -> 22
			// srcs: (29, 28)(622) 0, (23) 31 --> (1222) 0:NW28, ND0, *, NI1
			9'd28 : rdata = 43'b0001101011100011000001000010000000000000000;
			// PEs: 22, 22 -> 20
			// srcs: (30, 29)(623) 37, (23) 31 --> (1223) 1147:NW29, ND0, *, PEGB4
			9'd29 : rdata = 43'b0001101011101011000000000000000000011000000;
			// PEs: 21, 22 -> 17
			// srcs: (31, 32)(1191) 441, (1221) 465 --> (1746) 906:PENB, NI0, +, PEGB1
			9'd30 : rdata = 43'b0000111011110101000000000000000000010010000;
			// PEs: 21, 22 -> 17
			// srcs: (32, 33)(1192) 90, (1222) 0 --> (1765) 90:PENB, NI1, +, PEGB1
			9'd31 : rdata = 43'b0000111011110101000010000000000000010010000;
			// PEs: 18 -> 
			// srcs: (33, 30)(1101) 357 --> (1101) 357:PEGB2, pass, 
			9'd32 : rdata = 43'b1100011100100000000000000000000000000000000;
			// PEs: 17, 22 -> 17
			// srcs: (36, 31)(1071) 0, (1101) 357 --> (1744) 357:PEGB1, ALU, +, PEGB1
			9'd33 : rdata = 43'b0000111100010001111110000000000000010010000;
			// PEs: 16 -> 
			// srcs: (374, 34)(1595) 941 --> (1595) 941:PEGB0, pass, 
			9'd34 : rdata = 43'b1100011100000000000000000000000000000000000;
			// PEs: 22, 17 -> 17
			// srcs: (379, 35)(1595) 941, (1596) 803 --> (1600) 1744:ALU, PEGB1, +, PEGB1
			9'd35 : rdata = 43'b0000100111111111000100000000000000010010000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 23) begin
	always @(*) begin
		case(address)
			// PEs: 18 -> 23
			// srcs: (6, 2)(1074) 756 --> (1074) 756:PEGB2, pass, NI0
			9'd0 : rdata = 43'b1100011100100000000001000000000000000000000;
			// PEs: 20 -> 23
			// srcs: (7, 4)(1134) 130 --> (1134) 130:PEGB4, pass, NI1
			9'd1 : rdata = 43'b1100011101000000000001000010000000000000000;
			// PEs: 18 -> 23
			// srcs: (8, 14)(1075) 273 --> (1075) 273:PEGB2, pass, NI2
			9'd2 : rdata = 43'b1100011100100000000001000100000000000000000;
			// PEs: 17, 23 -> 23
			// srcs: (9, 3)(1044) 0, (1074) 756 --> (1231) 756:PEGB1, NI0, +, NI3
			9'd3 : rdata = 43'b0000111100010101000001000110000000000000000;
			// PEs: 19, 23 -> 23
			// srcs: (10, 5)(1104) 483, (1134) 130 --> (1232) 613:PEGB3, NI1, +, NI0
			9'd4 : rdata = 43'b0000111100110101000011000000000000000000000;
			// PEs: 18 -> 23
			// srcs: (11, 16)(1078) 798 --> (1078) 798:PEGB2, pass, NI1
			9'd5 : rdata = 43'b1100011100100000000001000010000000000000000;
			// PEs: 18 -> 23
			// srcs: (12, 18)(1079) 735 --> (1079) 735:PEGB2, pass, NI4
			9'd6 : rdata = 43'b1100011100100000000001001000000000000000000;
			// PEs: 17, 23 -> 23
			// srcs: (13, 15)(1045) 540, (1075) 273 --> (1250) 813:PEGB1, NI2, +, NI5
			9'd7 : rdata = 43'b0000111100010101000101001010000000000000000;
			// PEs: 16 -> 23
			// srcs: (14, 0)(834) 992 --> (834) 992:PEGB0, pass, NI2
			9'd8 : rdata = 43'b1100011100000000000001000100000000000000000;
			// PEs: 18 -> 23
			// srcs: (15, 36)(1082) 987 --> (1082) 987:PEGB2, pass, NI6
			9'd9 : rdata = 43'b1100011100100000000001001100000000000000000;
			// PEs: 18 -> 23
			// srcs: (16, 38)(1083) -63 --> (1083) -63:PEGB2, pass, NI7
			9'd10 : rdata = 43'b1100011100100000000001001110000000000000000;
			// PEs: 17, 23 -> 23
			// srcs: (17, 17)(1048) 504, (1078) 798 --> (1307) 1302:PEGB1, NI1, +, NI8
			9'd11 : rdata = 43'b0000111100010101000011010000000000000000000;
			// PEs: 18 -> 23
			// srcs: (18, 40)(1085) 168 --> (1085) 168:PEGB2, pass, NI1
			9'd12 : rdata = 43'b1100011100100000000001000010000000000000000;
			// PEs: 18 -> 23
			// srcs: (19, 50)(1086) -63 --> (1086) -63:PEGB2, pass, NI9
			9'd13 : rdata = 43'b1100011100100000000001010010000000000000000;
			// PEs: 17, 23 -> 23
			// srcs: (20, 19)(1049) 396, (1079) 735 --> (1326) 1131:PEGB1, NI4, +, NI10
			9'd14 : rdata = 43'b0000111100010101001001010100000000000000000;
			// PEs: 18 -> 23
			// srcs: (21, 60)(1088) 504 --> (1088) 504:PEGB2, pass, NI4
			9'd15 : rdata = 43'b1100011100100000000001001000000000000000000;
			// PEs: 18 -> 23
			// srcs: (22, 62)(1089) 294 --> (1089) 294:PEGB2, pass, NI11
			9'd16 : rdata = 43'b1100011100100000000001010110000000000000000;
			// PEs: 16, 23 -> 16
			// srcs: (23, 1)(804) 1395, (834) 992 --> (1227) 2387:PEGB0, NI2, +, PENB
			9'd17 : rdata = 43'b0000111100000101000100000000000000100000000;
			// PEs: 17, 23 -> 23
			// srcs: (24, 37)(1052) 144, (1082) 987 --> (1383) 1131:PEGB1, NI6, +, NI2
			9'd18 : rdata = 43'b0000111100010101001101000100000000000000000;
			// PEs: 16 -> 23
			// srcs: (25, 6)(835) 32 --> (835) 32:PEGB0, pass, NI6
			9'd19 : rdata = 43'b1100011100000000000001001100000000000000000;
			// PEs: 18 -> 23
			// srcs: (26, 64)(1093) 21 --> (1093) 21:PEGB2, pass, NI12
			9'd20 : rdata = 43'b1100011100100000000001011000000000000000000;
			// PEs: 18 -> 23
			// srcs: (27, 66)(1094) 378 --> (1094) 378:PEGB2, pass, NI13
			9'd21 : rdata = 43'b1100011100100000000001011010000000000000000;
			// PEs: 17, 23 -> 23
			// srcs: (28, 39)(1053) 1116, (1083) -63 --> (1402) 1053:PEGB1, NI7, +, NI14
			9'd22 : rdata = 43'b0000111100010101001111011100000000000000000;
			// PEs: 18 -> 23
			// srcs: (29, 68)(1096) 945 --> (1096) 945:PEGB2, pass, NI7
			9'd23 : rdata = 43'b1100011100100000000001001110000000000000000;
			// PEs: 18 -> 23
			// srcs: (30, 70)(1097) 777 --> (1097) 777:PEGB2, pass, NI15
			9'd24 : rdata = 43'b1100011100100000000001011110000000000000000;
			// PEs: 17, 23 -> 23
			// srcs: (31, 41)(1055) 1404, (1085) 168 --> (1440) 1572:PEGB1, NI1, +, NI16
			9'd25 : rdata = 43'b0000111100010101000011100000000000000000000;
			// PEs: 16, 23 -> 16
			// srcs: (34, 7)(805) 930, (835) 32 --> (1246) 962:PEGB0, NI6, +, PENB
			9'd26 : rdata = 43'b0000111100000101001100000000000000100000000;
			// PEs: 17, 23 -> 23
			// srcs: (35, 51)(1056) 756, (1086) -63 --> (1459) 693:PEGB1, NI9, +, NI1
			9'd27 : rdata = 43'b0000111100010101010011000010000000000000000;
			// PEs: 16 -> 23
			// srcs: (36, 8)(895) -23 --> (895) -23:PEGB0, pass, NI6
			9'd28 : rdata = 43'b1100011100000000000001001100000000000000000;
			// PEs: 17, 23 -> 23
			// srcs: (39, 61)(1058) 1260, (1088) 504 --> (1497) 1764:PEGB1, NI4, +, NI9
			9'd29 : rdata = 43'b0000111100010101001001010010000000000000000;
			// PEs: 17, 23 -> 23
			// srcs: (42, 63)(1059) 180, (1089) 294 --> (1516) 474:PEGB1, NI11, +, NI4
			9'd30 : rdata = 43'b0000111100010101010111001000000000000000000;
			// PEs: 16, 23 -> 23
			// srcs: (45, 9)(865) 1312, (895) -23 --> (1247) 1289:PEGB0, NI6, +, NI11
			9'd31 : rdata = 43'b0000111100000101001101010110000000000000000;
			// PEs: 17, 23 -> 23
			// srcs: (46, 65)(1063) 0, (1093) 21 --> (1592) 21:PEGB1, NI12, +, NI6
			9'd32 : rdata = 43'b0000111100010101011001001100000000000000000;
			// PEs: 16 -> 23
			// srcs: (47, 10)(955) 462 --> (955) 462:PEGB0, pass, NI12
			9'd33 : rdata = 43'b1100011100000000000001011000000000000000000;
			// PEs: 17, 23 -> 23
			// srcs: (50, 67)(1064) 324, (1094) 378 --> (1611) 702:PEGB1, NI13, +, NI17
			9'd34 : rdata = 43'b0000111100010101011011100010000000000000000;
			// PEs: 17, 23 -> 23
			// srcs: (53, 69)(1066) 864, (1096) 945 --> (1649) 1809:PEGB1, NI7, +, NI13
			9'd35 : rdata = 43'b0000111100010101001111011010000000000000000;
			// PEs: 16, 23 -> 23
			// srcs: (56, 11)(925) 638, (955) 462 --> (1248) 1100:PEGB0, NI12, +, NI7
			9'd36 : rdata = 43'b0000111100000101011001001110000000000000000;
			// PEs: 17, 23 -> 23
			// srcs: (57, 71)(1067) 1116, (1097) 777 --> (1668) 1893:PEGB1, NI15, +, NI12
			9'd37 : rdata = 43'b0000111100010101011111011000000000000000000;
			// PEs: 16 -> 23
			// srcs: (58, 12)(1015) 44 --> (1015) 44:PEGB0, pass, NI15
			9'd38 : rdata = 43'b1100011100000000000001011110000000000000000;
			// PEs: 23 -> 23
			// srcs: (59, 99)(1247) 1289 --> (1247) 1289:NI11, pass, NI11
			9'd39 : rdata = 43'b1100010101011000000001010110000000000000000;
			// PEs: 23, 23 -> 23
			// srcs: (59, 73)(1247) 1289, (1248) 1100 --> (1255) 2389:ALU, NI7, +, NI18
			9'd40 : rdata = 43'b0000100111111101001111100100000000000000000;
			// PEs: 16, 23 -> 17
			// srcs: (67, 13)(985) 52, (1015) 44 --> (1249) 96:PEGB0, NI15, +, PEGB1
			9'd41 : rdata = 43'b0000111100000101011110000000000000010010000;
			// PEs: 16 -> 23
			// srcs: (70, 20)(841) -96 --> (841) -96:PEGB0, pass, NI7
			9'd42 : rdata = 43'b1100011100000000000001001110000000000000000;
			// PEs: 23 -> 17
			// srcs: (77, 74)(1250) 813 --> (1250) 813:NI5, pass, PEGB1
			9'd43 : rdata = 43'b1100010100101000000000000000000000010010000;
			// PEs: 16, 23 -> 16
			// srcs: (79, 21)(811) 279, (841) -96 --> (1360) 183:PEGB0, NI7, +, PENB
			9'd44 : rdata = 43'b0000111100000101001110000000000000100000000;
			// PEs: 16 -> 
			// srcs: (81, 22)(901) -47 --> (901) -47:PEGB0, pass, 
			9'd45 : rdata = 43'b1100011100000000000000000000000000000000000;
			// PEs: 16, 23 -> 23
			// srcs: (90, 23)(871) 928, (901) -47 --> (1361) 881:PEGB0, ALU, +, NI5
			9'd46 : rdata = 43'b0000111100000001111111001010000000000000000;
			// PEs: 23 -> 17
			// srcs: (91, 92)(1255) 2389 --> (1255) 2389:NI18, pass, PEGB1
			9'd47 : rdata = 43'b1100010110010000000000000000000000010010000;
			// PEs: 16 -> 
			// srcs: (92, 24)(961) 363 --> (961) 363:PEGB0, pass, 
			9'd48 : rdata = 43'b1100011100000000000000000000000000000000000;
			// PEs: 16, 23 -> 23
			// srcs: (101, 25)(931) 464, (961) 363 --> (1362) 827:PEGB0, ALU, +, NI7
			9'd49 : rdata = 43'b0000111100000001111111001110000000000000000;
			// PEs: 16 -> 23
			// srcs: (103, 26)(1021) 880 --> (1021) 880:PEGB0, pass, NI11
			9'd50 : rdata = 43'b1100011100000000000001010110000000000000000;
			// PEs: 23 -> 23
			// srcs: (104, 100)(1361) 881 --> (1361) 881:NI5, pass, NI5
			9'd51 : rdata = 43'b1100010100101000000001001010000000000000000;
			// PEs: 23, 23 -> 23
			// srcs: (104, 77)(1361) 881, (1362) 827 --> (1369) 1708:ALU, NI7, +, NI15
			9'd52 : rdata = 43'b0000100111111101001111011110000000000000000;
			// PEs: 16, 23 -> 16
			// srcs: (112, 27)(991) 50, (1021) 880 --> (1363) 930:PEGB0, NI11, +, PENB
			9'd53 : rdata = 43'b0000111100000101010110000000000000100000000;
			// PEs: 16 -> 
			// srcs: (114, 28)(842) 416 --> (842) 416:PEGB0, pass, 
			9'd54 : rdata = 43'b1100011100000000000000000000000000000000000;
			// PEs: 16, 23 -> 16
			// srcs: (123, 29)(812) 1457, (842) 416 --> (1379) 1873:PEGB0, ALU, +, PENB
			9'd55 : rdata = 43'b0000111100000001111110000000000000100000000;
			// PEs: 16 -> 
			// srcs: (125, 30)(902) -45 --> (902) -45:PEGB0, pass, 
			9'd56 : rdata = 43'b1100011100000000000000000000000000000000000;
			// PEs: 16, 23 -> 23
			// srcs: (134, 31)(872) 1024, (902) -45 --> (1380) 979:PEGB0, ALU, +, NI5
			9'd57 : rdata = 43'b0000111100000001111111001010000000000000000;
			// PEs: 16 -> 
			// srcs: (136, 32)(962) 99 --> (962) 99:PEGB0, pass, 
			9'd58 : rdata = 43'b1100011100000000000000000000000000000000000;
			// PEs: 16, 23 -> 23
			// srcs: (145, 33)(932) 580, (962) 99 --> (1381) 679:PEGB0, ALU, +, NI7
			9'd59 : rdata = 43'b0000111100000001111111001110000000000000000;
			// PEs: 16 -> 23
			// srcs: (147, 34)(1022) 66 --> (1022) 66:PEGB0, pass, NI11
			9'd60 : rdata = 43'b1100011100000000000001010110000000000000000;
			// PEs: 23 -> 23
			// srcs: (148, 101)(1380) 979 --> (1380) 979:NI5, pass, NI5
			9'd61 : rdata = 43'b1100010100101000000001001010000000000000000;
			// PEs: 23, 23 -> 23
			// srcs: (148, 78)(1380) 979, (1381) 679 --> (1388) 1658:ALU, NI7, +, NI18
			9'd62 : rdata = 43'b0000100111111101001111100100000000000000000;
			// PEs: 16, 23 -> 23
			// srcs: (156, 35)(992) 50, (1022) 66 --> (1382) 116:PEGB0, NI11, +, NI5
			9'd63 : rdata = 43'b0000111100000101010111001010000000000000000;
			// PEs: 16 -> 23
			// srcs: (158, 42)(846) 448 --> (846) 448:PEGB0, pass, NI7
			9'd64 : rdata = 43'b1100011100000000000001001110000000000000000;
			// PEs: 23 -> 23
			// srcs: (159, 102)(1382) 116 --> (1382) 116:NI5, pass, NI5
			9'd65 : rdata = 43'b1100010100101000000001001010000000000000000;
			// PEs: 23, 23 -> 
			// srcs: (159, 79)(1382) 116, (1383) 1131 --> (1389) 1247:ALU, NI2, +, 
			9'd66 : rdata = 43'b0000100111111101000100000000000000000000000;
			// PEs: 23, 23 -> 23
			// srcs: (162, 94)(1388) 1658, (1389) 1247 --> (1392) 2905:NI18, ALU, +, NI2
			9'd67 : rdata = 43'b0000110110010001111111000100000000000000000;
			// PEs: 16, 23 -> 16
			// srcs: (167, 43)(816) 341, (846) 448 --> (1455) 789:PEGB0, NI7, +, PENB
			9'd68 : rdata = 43'b0000111100000101001110000000000000100000000;
			// PEs: 23 -> 16
			// srcs: (168, 72)(1231) 756 --> (1231) 756:NI3, pass, PENB
			9'd69 : rdata = 43'b1100010100011000000000000000000000100000000;
			// PEs: 16 -> 23
			// srcs: (169, 44)(906) -28 --> (906) -28:PEGB0, pass, NI3
			9'd70 : rdata = 43'b1100011100000000000001000110000000000000000;
			// PEs: 23 -> 16
			// srcs: (170, 75)(1307) 1302 --> (1307) 1302:NI8, pass, PENB
			9'd71 : rdata = 43'b1100010101000000000000000000000000100000000;
			// PEs: 23 -> 16
			// srcs: (171, 76)(1326) 1131 --> (1326) 1131:NI10, pass, PENB
			9'd72 : rdata = 43'b1100010101010000000000000000000000100000000;
			// PEs: 23 -> 16
			// srcs: (173, 80)(1402) 1053 --> (1402) 1053:NI14, pass, PENB
			9'd73 : rdata = 43'b1100010101110000000000000000000000100000000;
			// PEs: 23 -> 16
			// srcs: (174, 81)(1440) 1572 --> (1440) 1572:NI16, pass, PENB
			9'd74 : rdata = 43'b1100010110000000000000000000000000100000000;
			// PEs: 16, 23 -> 23
			// srcs: (178, 45)(876) 704, (906) -28 --> (1456) 676:PEGB0, NI3, +, NI5
			9'd75 : rdata = 43'b0000111100000101000111001010000000000000000;
			// PEs: 16 -> 23
			// srcs: (180, 46)(966) 1518 --> (966) 1518:PEGB0, pass, NI3
			9'd76 : rdata = 43'b1100011100000000000001000110000000000000000;
			// PEs: 23 -> 16
			// srcs: (181, 85)(1497) 1764 --> (1497) 1764:NI9, pass, PENB
			9'd77 : rdata = 43'b1100010101001000000000000000000000100000000;
			// PEs: 23 -> 16
			// srcs: (182, 86)(1516) 474 --> (1516) 474:NI4, pass, PENB
			9'd78 : rdata = 43'b1100010100100000000000000000000000100000000;
			// PEs: 16, 23 -> 23
			// srcs: (189, 47)(936) 290, (966) 1518 --> (1457) 1808:PEGB0, NI3, +, NI4
			9'd79 : rdata = 43'b0000111100000101000111001000000000000000000;
			// PEs: 16 -> 23
			// srcs: (191, 48)(1026) -22 --> (1026) -22:PEGB0, pass, NI3
			9'd80 : rdata = 43'b1100011100000000000001000110000000000000000;
			// PEs: 23 -> 23
			// srcs: (192, 103)(1456) 676 --> (1456) 676:NI5, pass, NI5
			9'd81 : rdata = 43'b1100010100101000000001001010000000000000000;
			// PEs: 23, 23 -> 23
			// srcs: (192, 82)(1456) 676, (1457) 1808 --> (1464) 2484:ALU, NI4, +, NI7
			9'd82 : rdata = 43'b0000100111111101001001001110000000000000000;
			// PEs: 16, 23 -> 23
			// srcs: (200, 49)(996) 64, (1026) -22 --> (1458) 42:PEGB0, NI3, +, NI4
			9'd83 : rdata = 43'b0000111100000101000111001000000000000000000;
			// PEs: 16 -> 23
			// srcs: (202, 52)(847) 1568 --> (847) 1568:PEGB0, pass, NI3
			9'd84 : rdata = 43'b1100011100000000000001000110000000000000000;
			// PEs: 23 -> 23
			// srcs: (203, 104)(1458) 42 --> (1458) 42:NI4, pass, NI4
			9'd85 : rdata = 43'b1100010100100000000001001000000000000000000;
			// PEs: 23, 23 -> 
			// srcs: (203, 83)(1458) 42, (1459) 693 --> (1465) 735:ALU, NI1, +, 
			9'd86 : rdata = 43'b0000100111111101000010000000000000000000000;
			// PEs: 23, 23 -> 23
			// srcs: (206, 95)(1464) 2484, (1465) 735 --> (1468) 3219:NI7, ALU, +, NI1
			9'd87 : rdata = 43'b0000110100111001111111000010000000000000000;
			// PEs: 16, 23 -> 16
			// srcs: (211, 53)(817) 372, (847) 1568 --> (1474) 1940:PEGB0, NI3, +, PENB
			9'd88 : rdata = 43'b0000111100000101000110000000000000100000000;
			// PEs: 16 -> 
			// srcs: (213, 54)(907) -13 --> (907) -13:PEGB0, pass, 
			9'd89 : rdata = 43'b1100011100000000000000000000000000000000000;
			// PEs: 16, 23 -> 23
			// srcs: (222, 55)(877) 1024, (907) -13 --> (1475) 1011:PEGB0, ALU, +, NI3
			9'd90 : rdata = 43'b0000111100000001111111000110000000000000000;
			// PEs: 16 -> 
			// srcs: (224, 56)(967) 1485 --> (967) 1485:PEGB0, pass, 
			9'd91 : rdata = 43'b1100011100000000000000000000000000000000000;
			// PEs: 16, 23 -> 23
			// srcs: (233, 57)(937) 551, (967) 1485 --> (1476) 2036:PEGB0, ALU, +, NI4
			9'd92 : rdata = 43'b0000111100000001111111001000000000000000000;
			// PEs: 16 -> 23
			// srcs: (235, 58)(1027) 792 --> (1027) 792:PEGB0, pass, NI5
			9'd93 : rdata = 43'b1100011100000000000001001010000000000000000;
			// PEs: 23 -> 23
			// srcs: (236, 105)(1475) 1011 --> (1475) 1011:NI3, pass, NI3
			9'd94 : rdata = 43'b1100010100011000000001000110000000000000000;
			// PEs: 23, 23 -> 23
			// srcs: (236, 84)(1475) 1011, (1476) 2036 --> (1483) 3047:ALU, NI4, +, NI7
			9'd95 : rdata = 43'b0000100111111101001001001110000000000000000;
			// PEs: 16, 23 -> 16
			// srcs: (244, 59)(997) 78, (1027) 792 --> (1477) 870:PEGB0, NI5, +, PENB
			9'd96 : rdata = 43'b0000111100000101001010000000000000100000000;
			// PEs: 23 -> 16
			// srcs: (249, 91)(1232) 613 --> (1232) 613:NI0, pass, PENB
			9'd97 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 23 -> 16
			// srcs: (257, 93)(1369) 1708 --> (1369) 1708:NI15, pass, PENB
			9'd98 : rdata = 43'b1100010101111000000000000000000000100000000;
			// PEs: 23 -> 16
			// srcs: (262, 96)(1483) 3047 --> (1483) 3047:NI7, pass, PENB
			9'd99 : rdata = 43'b1100010100111000000000000000000000100000000;
			// PEs: 23 -> 17
			// srcs: (299, 88)(1611) 702 --> (1611) 702:NI17, pass, PEGB1
			9'd100 : rdata = 43'b1100010110001000000000000000000000010010000;
			// PEs: 23 -> 16
			// srcs: (326, 97)(1392) 2905 --> (1392) 2905:NI2, pass, PENB
			9'd101 : rdata = 43'b1100010100010000000000000000000000100000000;
			// PEs: 23 -> 17
			// srcs: (347, 89)(1649) 1809 --> (1649) 1809:NI13, pass, PEGB1
			9'd102 : rdata = 43'b1100010101101000000000000000000000010010000;
			// PEs: 23 -> 17
			// srcs: (369, 87)(1592) 21 --> (1592) 21:NI6, pass, PEGB1
			9'd103 : rdata = 43'b1100010100110000000000000000000000010010000;
			// PEs: 23 -> 17
			// srcs: (371, 90)(1668) 1893 --> (1668) 1893:NI12, pass, PEGB1
			9'd104 : rdata = 43'b1100010101100000000000000000000000010010000;
			// PEs: 23 -> 16
			// srcs: (1021, 98)(1468) 3219 --> (1468) 3219:NI1, pass, PENB
			9'd105 : rdata = 43'b1100010100001000000000000000000000100000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 24) begin
	always @(*) begin
		case(address)
			// PEs: 0 -> 24
			// srcs: (11, 0)(624) 84 --> (624) 84:PUGB0, pass, NI0
			9'd0 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 0 -> 25
			// srcs: (12, 1)(654) 11 --> (654) 11:PUGB0, pass, PENB
			9'd1 : rdata = 43'b1100011100001000000000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (18, 2)(624) 84 --> (624) 84:NI0, pass, PENB
			9'd2 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 16 -> 24
			// srcs: (19, 3)(1164) -9 --> (1164) -9:PUNB, pass, NI0
			9'd3 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 16 -> 25
			// srcs: (20, 4)(1194) 341 --> (1194) 341:PUNB, pass, PENB
			9'd4 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 25 -> 48
			// srcs: (25, 195)(1224) 95 --> (1224) 95:PEGB1, pass, PUGB6
			9'd5 : rdata = 43'b1100011100010000000000000000000000000001110;
			// PEs: 24 -> 25
			// srcs: (26, 5)(1164) -9 --> (1164) -9:NI0, pass, PENB
			9'd6 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 24
			// srcs: (27, 6)(625) 560 --> (625) 560:PUGB0, pass, NI0
			9'd7 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 0 -> 25
			// srcs: (28, 7)(655) 176 --> (655) 176:PUGB0, pass, PENB
			9'd8 : rdata = 43'b1100011100001000000000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (34, 8)(625) 560 --> (625) 560:NI0, pass, PENB
			9'd9 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 24
			// srcs: (35, 9)(685) 864 --> (685) 864:PUGB0, pass, NI0
			9'd10 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 0 -> 25
			// srcs: (36, 10)(715) 1104 --> (715) 1104:PUGB0, pass, PENB
			9'd11 : rdata = 43'b1100011100001000000000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (42, 11)(685) 864 --> (685) 864:NI0, pass, PENB
			9'd12 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 24
			// srcs: (43, 12)(745) 1008 --> (745) 1008:PUGB0, pass, NI0
			9'd13 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 0 -> 25
			// srcs: (44, 13)(775) 551 --> (775) 551:PUGB0, pass, PENB
			9'd14 : rdata = 43'b1100011100001000000000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (50, 14)(745) 1008 --> (745) 1008:NI0, pass, PENB
			9'd15 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 16 -> 24
			// srcs: (51, 15)(1105) 897 --> (1105) 897:PUNB, pass, NI0
			9'd16 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 16 -> 25
			// srcs: (52, 16)(1135) -39 --> (1135) -39:PUNB, pass, PENB
			9'd17 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (58, 17)(1105) 897 --> (1105) 897:NI0, pass, PENB
			9'd18 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 16 -> 24
			// srcs: (59, 18)(1165) 117 --> (1165) 117:PUNB, pass, NI0
			9'd19 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 16 -> 25
			// srcs: (60, 19)(1195) 93 --> (1195) 93:PUNB, pass, PENB
			9'd20 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (66, 20)(1165) 117 --> (1165) 117:NI0, pass, PENB
			9'd21 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 24
			// srcs: (67, 21)(626) 364 --> (626) 364:PUGB0, pass, NI0
			9'd22 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 0 -> 25
			// srcs: (68, 22)(656) 121 --> (656) 121:PUGB0, pass, PENB
			9'd23 : rdata = 43'b1100011100001000000000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (74, 23)(626) 364 --> (626) 364:NI0, pass, PENB
			9'd24 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 24
			// srcs: (75, 24)(686) 816 --> (686) 816:PUGB0, pass, NI0
			9'd25 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 0 -> 25
			// srcs: (76, 25)(716) 644 --> (716) 644:PUGB0, pass, PENB
			9'd26 : rdata = 43'b1100011100001000000000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (82, 26)(686) 816 --> (686) 816:NI0, pass, PENB
			9'd27 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 24
			// srcs: (83, 27)(746) 792 --> (746) 792:PUGB0, pass, NI0
			9'd28 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 0 -> 25
			// srcs: (84, 28)(776) 361 --> (776) 361:PUGB0, pass, PENB
			9'd29 : rdata = 43'b1100011100001000000000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (90, 29)(746) 792 --> (746) 792:NI0, pass, PENB
			9'd30 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 24
			// srcs: (91, 30)(806) 372 --> (806) 372:PUGB0, pass, NI0
			9'd31 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 8 -> 25
			// srcs: (92, 31)(836) 672 --> (836) 672:PUGB1, pass, PENB
			9'd32 : rdata = 43'b1100011100011000000000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (98, 32)(806) 372 --> (806) 372:NI0, pass, PENB
			9'd33 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 8 -> 24
			// srcs: (99, 33)(866) 416 --> (866) 416:PUGB1, pass, NI0
			9'd34 : rdata = 43'b1100011100011000000001000000000000000000000;
			// PEs: 8 -> 25
			// srcs: (100, 34)(896) -5 --> (896) -5:PUGB1, pass, PENB
			9'd35 : rdata = 43'b1100011100011000000000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (106, 35)(866) 416 --> (866) 416:NI0, pass, PENB
			9'd36 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 16 -> 24
			// srcs: (107, 36)(1046) 1152 --> (1046) 1152:PUNB, pass, NI0
			9'd37 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 16 -> 25
			// srcs: (108, 37)(1076) 273 --> (1076) 273:PUNB, pass, PENB
			9'd38 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 25 -> 56
			// srcs: (113, 197)(1266) 411 --> (1266) 411:PEGB1, pass, PUGB7
			9'd39 : rdata = 43'b1100011100010000000000000000000000000001111;
			// PEs: 24 -> 25
			// srcs: (114, 38)(1046) 1152 --> (1046) 1152:NI0, pass, PENB
			9'd40 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 16 -> 24
			// srcs: (115, 39)(1106) 437 --> (1106) 437:PUNB, pass, NI0
			9'd41 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 16 -> 25
			// srcs: (116, 40)(1136) 468 --> (1136) 468:PUNB, pass, PENB
			9'd42 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 25 -> 56
			// srcs: (121, 198)(1269) 1425 --> (1269) 1425:PEGB1, pass, PUGB7
			9'd43 : rdata = 43'b1100011100010000000000000000000000000001111;
			// PEs: 24 -> 25
			// srcs: (122, 41)(1106) 437 --> (1106) 437:NI0, pass, PENB
			9'd44 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 16 -> 24
			// srcs: (123, 42)(1166) 162 --> (1166) 162:PUNB, pass, NI0
			9'd45 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 16 -> 25
			// srcs: (124, 43)(1196) 1240 --> (1196) 1240:PUNB, pass, PENB
			9'd46 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (130, 44)(1166) 162 --> (1166) 162:NI0, pass, PENB
			9'd47 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 16 -> 24
			// srcs: (131, 45)(1108) 1058 --> (1108) 1058:PUNB, pass, NI0
			9'd48 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 16 -> 25
			// srcs: (132, 46)(1138) 429 --> (1138) 429:PUNB, pass, PENB
			9'd49 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (138, 47)(1108) 1058 --> (1108) 1058:NI0, pass, PENB
			9'd50 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 16 -> 24
			// srcs: (139, 48)(1168) 45 --> (1168) 45:PUNB, pass, NI0
			9'd51 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 16 -> 25
			// srcs: (140, 49)(1198) 1488 --> (1198) 1488:PUNB, pass, PENB
			9'd52 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (146, 50)(1168) 45 --> (1168) 45:NI0, pass, PENB
			9'd53 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 16 -> 24
			// srcs: (147, 51)(1109) 46 --> (1109) 46:PUNB, pass, NI0
			9'd54 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 16 -> 25
			// srcs: (148, 52)(1139) 143 --> (1139) 143:PUNB, pass, PENB
			9'd55 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (154, 53)(1109) 46 --> (1109) 46:NI0, pass, PENB
			9'd56 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 16 -> 24
			// srcs: (155, 54)(1169) 405 --> (1169) 405:PUNB, pass, NI0
			9'd57 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 16 -> 25
			// srcs: (156, 55)(1199) -62 --> (1199) -62:PUNB, pass, PENB
			9'd58 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (162, 56)(1169) 405 --> (1169) 405:NI0, pass, PENB
			9'd59 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 16 -> 24
			// srcs: (163, 57)(1050) 1332 --> (1050) 1332:PUNB, pass, NI0
			9'd60 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 16 -> 25
			// srcs: (164, 58)(1080) 483 --> (1080) 483:PUNB, pass, PENB
			9'd61 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (170, 59)(1050) 1332 --> (1050) 1332:NI0, pass, PENB
			9'd62 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 16 -> 24
			// srcs: (171, 60)(1110) 391 --> (1110) 391:PUNB, pass, NI0
			9'd63 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 16 -> 25
			// srcs: (172, 61)(1140) 39 --> (1140) 39:PUNB, pass, PENB
			9'd64 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 25 -> 16
			// srcs: (173, 223)(1333) 532 --> (1333) 532:PEGB1, pass, PUGB2
			9'd65 : rdata = 43'b1100011100010000000000000000000000000001010;
			// PEs: 25 -> 8
			// srcs: (177, 199)(1345) 1815 --> (1345) 1815:PEGB1, pass, PUGB1
			9'd66 : rdata = 43'b1100011100010000000000000000000000000001001;
			// PEs: 24 -> 25
			// srcs: (178, 62)(1110) 391 --> (1110) 391:NI0, pass, PENB
			9'd67 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 16 -> 24
			// srcs: (179, 63)(1170) -9 --> (1170) -9:PUNB, pass, NI0
			9'd68 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 16 -> 25
			// srcs: (180, 64)(1200) 434 --> (1200) 434:PUNB, pass, PENB
			9'd69 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (186, 65)(1170) -9 --> (1170) -9:NI0, pass, PENB
			9'd70 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 24
			// srcs: (187, 66)(631) 28 --> (631) 28:PUGB0, pass, NI0
			9'd71 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 0 -> 25
			// srcs: (188, 67)(661) 99 --> (661) 99:PUGB0, pass, PENB
			9'd72 : rdata = 43'b1100011100001000000000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (194, 68)(631) 28 --> (631) 28:NI0, pass, PENB
			9'd73 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 24
			// srcs: (195, 69)(691) 240 --> (691) 240:PUGB0, pass, NI0
			9'd74 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 0 -> 25
			// srcs: (196, 70)(721) 506 --> (721) 506:PUGB0, pass, PENB
			9'd75 : rdata = 43'b1100011100001000000000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (202, 71)(691) 240 --> (691) 240:NI0, pass, PENB
			9'd76 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 24
			// srcs: (203, 72)(751) 552 --> (751) 552:PUGB0, pass, NI0
			9'd77 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 0 -> 25
			// srcs: (204, 73)(781) 114 --> (781) 114:PUGB0, pass, PENB
			9'd78 : rdata = 43'b1100011100001000000000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (210, 74)(751) 552 --> (751) 552:NI0, pass, PENB
			9'd79 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 16 -> 24
			// srcs: (211, 75)(1051) 108 --> (1051) 108:PUNB, pass, NI0
			9'd80 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 16 -> 25
			// srcs: (212, 76)(1081) 231 --> (1081) 231:PUNB, pass, PENB
			9'd81 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (218, 77)(1051) 108 --> (1051) 108:NI0, pass, PENB
			9'd82 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 16 -> 24
			// srcs: (219, 78)(1111) 437 --> (1111) 437:PUNB, pass, NI0
			9'd83 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 16 -> 25
			// srcs: (220, 79)(1141) 91 --> (1141) 91:PUNB, pass, PENB
			9'd84 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (226, 80)(1111) 437 --> (1111) 437:NI0, pass, PENB
			9'd85 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 16 -> 24
			// srcs: (227, 81)(1171) 369 --> (1171) 369:PUNB, pass, NI0
			9'd86 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 16 -> 25
			// srcs: (228, 82)(1201) 186 --> (1201) 186:PUNB, pass, PENB
			9'd87 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (234, 83)(1171) 369 --> (1171) 369:NI0, pass, PENB
			9'd88 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 16 -> 24
			// srcs: (235, 84)(1112) 161 --> (1112) 161:PUNB, pass, NI0
			9'd89 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 16 -> 25
			// srcs: (236, 85)(1142) 91 --> (1142) 91:PUNB, pass, PENB
			9'd90 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (242, 86)(1112) 161 --> (1112) 161:NI0, pass, PENB
			9'd91 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 16 -> 24
			// srcs: (243, 87)(1172) 369 --> (1172) 369:PUNB, pass, NI0
			9'd92 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 16 -> 25
			// srcs: (244, 88)(1202) 1333 --> (1202) 1333:PUNB, pass, PENB
			9'd93 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (250, 89)(1172) 369 --> (1172) 369:NI0, pass, PENB
			9'd94 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 16 -> 24
			// srcs: (251, 90)(1054) 1188 --> (1054) 1188:PUNB, pass, NI0
			9'd95 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 16 -> 25
			// srcs: (252, 91)(1084) 525 --> (1084) 525:PUNB, pass, PENB
			9'd96 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (258, 92)(1054) 1188 --> (1054) 1188:NI0, pass, PENB
			9'd97 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 16 -> 24
			// srcs: (259, 93)(1114) 483 --> (1114) 483:PUNB, pass, NI0
			9'd98 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 16 -> 25
			// srcs: (260, 94)(1144) 13 --> (1144) 13:PUNB, pass, PENB
			9'd99 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (266, 95)(1114) 483 --> (1114) 483:NI0, pass, PENB
			9'd100 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 16 -> 24
			// srcs: (267, 96)(1174) 162 --> (1174) 162:PUNB, pass, NI0
			9'd101 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 16 -> 25
			// srcs: (268, 97)(1204) 1302 --> (1204) 1302:PUNB, pass, PENB
			9'd102 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (274, 98)(1174) 162 --> (1174) 162:NI0, pass, PENB
			9'd103 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 24
			// srcs: (275, 99)(696) 792 --> (696) 792:PUGB0, pass, NI0
			9'd104 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 0 -> 25
			// srcs: (276, 100)(726) 1242 --> (726) 1242:PUGB0, pass, PENB
			9'd105 : rdata = 43'b1100011100001000000000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (282, 101)(696) 792 --> (696) 792:NI0, pass, PENB
			9'd106 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 24
			// srcs: (283, 102)(756) 72 --> (756) 72:PUGB0, pass, NI0
			9'd107 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 0 -> 25
			// srcs: (284, 103)(786) 266 --> (786) 266:PUGB0, pass, PENB
			9'd108 : rdata = 43'b1100011100001000000000000000000000100000000;
			// PEs: 25 -> 32
			// srcs: (289, 203)(1453) 2034 --> (1453) 2034:PEGB1, pass, PUNB
			9'd109 : rdata = 43'b1100011100010000000000000000000001000000000;
			// PEs: 24 -> 25
			// srcs: (290, 104)(756) 72 --> (756) 72:NI0, pass, PENB
			9'd110 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 16 -> 24
			// srcs: (291, 105)(1116) 598 --> (1116) 598:PUNB, pass, NI0
			9'd111 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 16 -> 25
			// srcs: (292, 106)(1146) 195 --> (1146) 195:PUNB, pass, PENB
			9'd112 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (298, 107)(1116) 598 --> (1116) 598:NI0, pass, PENB
			9'd113 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 16 -> 24
			// srcs: (299, 108)(1176) 360 --> (1176) 360:PUNB, pass, NI0
			9'd114 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 16 -> 25
			// srcs: (300, 109)(1206) 1178 --> (1206) 1178:PUNB, pass, PENB
			9'd115 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (306, 110)(1176) 360 --> (1176) 360:NI0, pass, PENB
			9'd116 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 24
			// srcs: (307, 111)(637) 84 --> (637) 84:PUGB0, pass, NI0
			9'd117 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 0 -> 25
			// srcs: (308, 112)(667) 0 --> (667) 0:PUGB0, pass, PENB
			9'd118 : rdata = 43'b1100011100001000000000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (314, 113)(637) 84 --> (637) 84:NI0, pass, PENB
			9'd119 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 24
			// srcs: (315, 114)(697) 1176 --> (697) 1176:PUGB0, pass, NI0
			9'd120 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 0 -> 25
			// srcs: (316, 115)(727) 184 --> (727) 184:PUGB0, pass, PENB
			9'd121 : rdata = 43'b1100011100001000000000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (322, 116)(697) 1176 --> (697) 1176:NI0, pass, PENB
			9'd122 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 24
			// srcs: (323, 117)(757) 888 --> (757) 888:PUGB0, pass, NI0
			9'd123 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 0 -> 25
			// srcs: (324, 118)(787) 741 --> (787) 741:PUGB0, pass, PENB
			9'd124 : rdata = 43'b1100011100001000000000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (330, 119)(757) 888 --> (757) 888:NI0, pass, PENB
			9'd125 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 16 -> 24
			// srcs: (331, 120)(1057) 1080 --> (1057) 1080:PUNB, pass, NI0
			9'd126 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 16 -> 25
			// srcs: (332, 121)(1087) 903 --> (1087) 903:PUNB, pass, PENB
			9'd127 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (338, 122)(1057) 1080 --> (1057) 1080:NI0, pass, PENB
			9'd128 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 16 -> 24
			// srcs: (339, 123)(1117) 1035 --> (1117) 1035:PUNB, pass, NI0
			9'd129 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 16 -> 25
			// srcs: (340, 124)(1147) 377 --> (1147) 377:PUNB, pass, PENB
			9'd130 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (346, 125)(1117) 1035 --> (1117) 1035:NI0, pass, PENB
			9'd131 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 16 -> 24
			// srcs: (347, 126)(1177) 396 --> (1177) 396:PUNB, pass, NI0
			9'd132 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 16 -> 25
			// srcs: (348, 127)(1207) 372 --> (1207) 372:PUNB, pass, PENB
			9'd133 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (354, 128)(1177) 396 --> (1177) 396:NI0, pass, PENB
			9'd134 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 16 -> 24
			// srcs: (355, 129)(1118) 391 --> (1118) 391:PUNB, pass, NI0
			9'd135 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 16 -> 25
			// srcs: (356, 130)(1148) 273 --> (1148) 273:PUNB, pass, PENB
			9'd136 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (362, 131)(1118) 391 --> (1118) 391:NI0, pass, PENB
			9'd137 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 16 -> 24
			// srcs: (363, 132)(1178) 81 --> (1178) 81:PUNB, pass, NI0
			9'd138 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 16 -> 25
			// srcs: (364, 133)(1208) -62 --> (1208) -62:PUNB, pass, PENB
			9'd139 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (370, 134)(1178) 81 --> (1178) 81:NI0, pass, PENB
			9'd140 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 24
			// srcs: (371, 135)(639) 56 --> (639) 56:PUGB0, pass, NI0
			9'd141 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 0 -> 25
			// srcs: (372, 136)(669) 187 --> (669) 187:PUGB0, pass, PENB
			9'd142 : rdata = 43'b1100011100001000000000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (378, 137)(639) 56 --> (639) 56:NI0, pass, PENB
			9'd143 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 24
			// srcs: (379, 138)(699) 408 --> (699) 408:PUGB0, pass, NI0
			9'd144 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 0 -> 25
			// srcs: (380, 139)(729) 1472 --> (729) 1472:PUGB0, pass, PENB
			9'd145 : rdata = 43'b1100011100001000000000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (386, 140)(699) 408 --> (699) 408:NI0, pass, PENB
			9'd146 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 24
			// srcs: (387, 141)(759) 840 --> (759) 840:PUGB0, pass, NI0
			9'd147 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 0 -> 25
			// srcs: (388, 142)(789) 532 --> (789) 532:PUGB0, pass, PENB
			9'd148 : rdata = 43'b1100011100001000000000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (394, 143)(759) 840 --> (759) 840:NI0, pass, PENB
			9'd149 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 16 -> 24
			// srcs: (395, 144)(1119) 322 --> (1119) 322:PUNB, pass, NI0
			9'd150 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 16 -> 25
			// srcs: (396, 145)(1149) 429 --> (1149) 429:PUNB, pass, PENB
			9'd151 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 25 -> 32
			// srcs: (401, 207)(1511) 1372 --> (1511) 1372:PEGB1, pass, PUNB
			9'd152 : rdata = 43'b1100011100010000000000000000000001000000000;
			// PEs: 24 -> 25
			// srcs: (402, 146)(1119) 322 --> (1119) 322:NI0, pass, PENB
			9'd153 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 16 -> 24
			// srcs: (403, 147)(1179) 333 --> (1179) 333:PUNB, pass, NI0
			9'd154 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 16 -> 25
			// srcs: (404, 148)(1209) 806 --> (1209) 806:PUNB, pass, PENB
			9'd155 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (410, 149)(1179) 333 --> (1179) 333:NI0, pass, PENB
			9'd156 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 16 -> 24
			// srcs: (411, 150)(1060) 720 --> (1060) 720:PUNB, pass, NI0
			9'd157 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 16 -> 25
			// srcs: (412, 151)(1090) 588 --> (1090) 588:PUNB, pass, PENB
			9'd158 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (418, 152)(1060) 720 --> (1060) 720:NI0, pass, PENB
			9'd159 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 16 -> 24
			// srcs: (419, 153)(1120) 437 --> (1120) 437:PUNB, pass, NI0
			9'd160 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 16 -> 25
			// srcs: (420, 154)(1150) 559 --> (1150) 559:PUNB, pass, PENB
			9'd161 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 25 -> 16
			// srcs: (421, 229)(1523) 1890 --> (1523) 1890:PEGB1, pass, PUGB2
			9'd162 : rdata = 43'b1100011100010000000000000000000000000001010;
			// PEs: 25 -> 48
			// srcs: (425, 208)(1535) 1308 --> (1535) 1308:PEGB1, pass, PUGB6
			9'd163 : rdata = 43'b1100011100010000000000000000000000000001110;
			// PEs: 24 -> 25
			// srcs: (426, 155)(1120) 437 --> (1120) 437:NI0, pass, PENB
			9'd164 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 16 -> 24
			// srcs: (427, 156)(1180) 261 --> (1180) 261:PUNB, pass, NI0
			9'd165 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 16 -> 25
			// srcs: (428, 157)(1210) 1209 --> (1210) 1209:PUNB, pass, PENB
			9'd166 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (434, 158)(1180) 261 --> (1180) 261:NI0, pass, PENB
			9'd167 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 16 -> 24
			// srcs: (435, 159)(1062) 612 --> (1062) 612:PUNB, pass, NI0
			9'd168 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 16 -> 25
			// srcs: (436, 160)(1092) 672 --> (1092) 672:PUNB, pass, PENB
			9'd169 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (442, 161)(1062) 612 --> (1062) 612:NI0, pass, PENB
			9'd170 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 16 -> 24
			// srcs: (443, 162)(1122) 920 --> (1122) 920:PUNB, pass, NI0
			9'd171 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 16 -> 25
			// srcs: (444, 163)(1152) 312 --> (1152) 312:PUNB, pass, PENB
			9'd172 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 25 -> 16
			// srcs: (445, 230)(1542) 2466 --> (1542) 2466:PEGB1, pass, PUGB2
			9'd173 : rdata = 43'b1100011100010000000000000000000000000001010;
			// PEs: 25 -> 56
			// srcs: (449, 209)(1573) 1284 --> (1573) 1284:PEGB1, pass, PUGB7
			9'd174 : rdata = 43'b1100011100010000000000000000000000000001111;
			// PEs: 24 -> 25
			// srcs: (450, 164)(1122) 920 --> (1122) 920:NI0, pass, PENB
			9'd175 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 16 -> 24
			// srcs: (451, 165)(1182) 297 --> (1182) 297:PUNB, pass, NI0
			9'd176 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 16 -> 25
			// srcs: (452, 166)(1212) 1085 --> (1212) 1085:PUNB, pass, PENB
			9'd177 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (458, 167)(1182) 297 --> (1182) 297:NI0, pass, PENB
			9'd178 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 16 -> 24
			// srcs: (459, 168)(1124) 1127 --> (1124) 1127:PUNB, pass, NI0
			9'd179 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 16 -> 25
			// srcs: (460, 169)(1154) 273 --> (1154) 273:PUNB, pass, PENB
			9'd180 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (466, 170)(1124) 1127 --> (1124) 1127:NI0, pass, PENB
			9'd181 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 16 -> 24
			// srcs: (467, 171)(1184) 81 --> (1184) 81:PUNB, pass, NI0
			9'd182 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 16 -> 25
			// srcs: (468, 172)(1214) -31 --> (1214) -31:PUNB, pass, PENB
			9'd183 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 25 -> 16
			// srcs: (469, 231)(1580) 2614 --> (1580) 2614:PEGB1, pass, PUGB2
			9'd184 : rdata = 43'b1100011100010000000000000000000000000001010;
			// PEs: 24 -> 25
			// srcs: (474, 173)(1184) 81 --> (1184) 81:NI0, pass, PENB
			9'd185 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 16 -> 24
			// srcs: (475, 174)(1065) 864 --> (1065) 864:PUNB, pass, NI0
			9'd186 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 16 -> 25
			// srcs: (476, 175)(1095) 609 --> (1095) 609:PUNB, pass, PENB
			9'd187 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (482, 176)(1065) 864 --> (1065) 864:NI0, pass, PENB
			9'd188 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 16 -> 24
			// srcs: (483, 177)(1125) 138 --> (1125) 138:PUNB, pass, NI0
			9'd189 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 16 -> 25
			// srcs: (484, 178)(1155) 0 --> (1155) 0:PUNB, pass, PENB
			9'd190 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 25 -> 8
			// srcs: (489, 210)(1630) 1473 --> (1630) 1473:PEGB1, pass, PUGB1
			9'd191 : rdata = 43'b1100011100010000000000000000000000000001001;
			// PEs: 24 -> 25
			// srcs: (490, 179)(1125) 138 --> (1125) 138:NI0, pass, PENB
			9'd192 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 16 -> 24
			// srcs: (491, 180)(1185) 144 --> (1185) 144:PUNB, pass, NI0
			9'd193 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 16 -> 25
			// srcs: (492, 181)(1215) -93 --> (1215) -93:PUNB, pass, PENB
			9'd194 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (498, 182)(1185) 144 --> (1185) 144:NI0, pass, PENB
			9'd195 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 16 -> 24
			// srcs: (499, 183)(1126) 897 --> (1126) 897:PUNB, pass, NI0
			9'd196 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 16 -> 25
			// srcs: (500, 184)(1156) 39 --> (1156) 39:PUNB, pass, PENB
			9'd197 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 25 -> 8
			// srcs: (501, 222)(1314) 3020 --> (1314) 3020:PEGB1, pass, PUGB1
			9'd198 : rdata = 43'b1100011100010000000000000000000000000001001;
			// PEs: 24 -> 25
			// srcs: (506, 185)(1126) 897 --> (1126) 897:NI0, pass, PENB
			9'd199 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 16 -> 24
			// srcs: (507, 186)(1186) 198 --> (1186) 198:PUNB, pass, NI0
			9'd200 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 16 -> 25
			// srcs: (508, 187)(1216) 341 --> (1216) 341:PUNB, pass, PENB
			9'd201 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 25 -> 8
			// srcs: (509, 225)(1390) 1954 --> (1390) 1954:PEGB1, pass, PUGB1
			9'd202 : rdata = 43'b1100011100010000000000000000000000000001001;
			// PEs: 24 -> 25
			// srcs: (514, 188)(1186) 198 --> (1186) 198:NI0, pass, PENB
			9'd203 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 16 -> 24
			// srcs: (515, 189)(1127) 989 --> (1127) 989:PUNB, pass, NI0
			9'd204 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 16 -> 25
			// srcs: (516, 190)(1157) 195 --> (1157) 195:PUNB, pass, PENB
			9'd205 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 25 -> 8
			// srcs: (517, 226)(1428) 1960 --> (1428) 1960:PEGB1, pass, PUGB1
			9'd206 : rdata = 43'b1100011100010000000000000000000000000001001;
			// PEs: 24 -> 25
			// srcs: (522, 191)(1127) 989 --> (1127) 989:NI0, pass, PENB
			9'd207 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 16 -> 24
			// srcs: (523, 192)(1187) 441 --> (1187) 441:PUNB, pass, NI0
			9'd208 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 16 -> 25
			// srcs: (524, 193)(1217) 310 --> (1217) 310:PUNB, pass, PENB
			9'd209 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (530, 194)(1187) 441 --> (1187) 441:NI0, pass, PENB
			9'd210 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 16 -> 25
			// srcs: (531, 196)(1246) 962 --> (1246) 962:PUNB, pass, PENB
			9'd211 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 16 -> 25
			// srcs: (532, 200)(1360) 183 --> (1360) 183:PUNB, pass, PENB
			9'd212 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 16 -> 25
			// srcs: (533, 201)(1363) 930 --> (1363) 930:PUNB, pass, PENB
			9'd213 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 48 -> 25
			// srcs: (534, 202)(1420) 858 --> (1420) 858:PUGB6, pass, PENB
			9'd214 : rdata = 43'b1100011101101000000000000000000000100000000;
			// PEs: 16 -> 25
			// srcs: (535, 204)(1455) 789 --> (1455) 789:PUNB, pass, PENB
			9'd215 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 16 -> 25
			// srcs: (536, 205)(1474) 1940 --> (1474) 1940:PUNB, pass, PENB
			9'd216 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 16 -> 25
			// srcs: (537, 206)(1477) 870 --> (1477) 870:PUNB, pass, PENB
			9'd217 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 0 -> 24
			// srcs: (538, 211)(1701) 1049 --> (1701) 1049:PUGB0, pass, NI0
			9'd218 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 8 -> 25
			// srcs: (539, 212)(1702) 1312 --> (1702) 1312:PUGB1, pass, PENB
			9'd219 : rdata = 43'b1100011100011000000000000000000000100000000;
			// PEs: 25 -> 48
			// srcs: (541, 219)(1427) 2571 --> (1427) 2571:PEGB1, pass, PUGB6
			9'd220 : rdata = 43'b1100011100010000000000000000000000000001110;
			// PEs: 25 -> 32
			// srcs: (542, 215)(1463) 1127 --> (1463) 1127:PEGB1, pass, PUNB
			9'd221 : rdata = 43'b1100011100010000000000000000000001000000000;
			// PEs: 24 -> 25
			// srcs: (545, 213)(1701) 1049 --> (1701) 1049:NI0, pass, PENB
			9'd222 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 16 -> 25
			// srcs: (546, 214)(1232) 613 --> (1232) 613:PUNB, pass, PENB
			9'd223 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 16 -> 27
			// srcs: (547, 218)(1369) 1708 --> (1369) 1708:PUNB, pass, PEGB3
			9'd224 : rdata = 43'b1100011011111000000000000000000000010110000;
			// PEs: 16 -> 26
			// srcs: (548, 220)(1483) 3047 --> (1483) 3047:PUNB, pass, PEGB2
			9'd225 : rdata = 43'b1100011011111000000000000000000000010100000;
			// PEs: 16 -> 24
			// srcs: (549, 236)(1694) 840 --> (1694) 840:PUNB, pass, NI0
			9'd226 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 25 -> 32
			// srcs: (551, 216)(1519) 2123 --> (1519) 2123:PEGB1, pass, PUNB
			9'd227 : rdata = 43'b1100011100010000000000000000000001000000000;
			// PEs: 25 -> 32
			// srcs: (552, 217)(1710) 2361 --> (1710) 2361:PEGB1, pass, PUNB
			9'd228 : rdata = 43'b1100011100010000000000000000000001000000000;
			// PEs: 25 -> 0
			// srcs: (553, 221)(1238) 945 --> (1238) 945:PEGB1, pass, PUGB0
			9'd229 : rdata = 43'b1100011100010000000000000000000000000001000;
			// PEs: 25 -> 32
			// srcs: (561, 224)(1352) 855 --> (1352) 855:PEGB1, pass, PUNB
			9'd230 : rdata = 43'b1100011100010000000000000000000001000000000;
			// PEs: 25 -> 32
			// srcs: (569, 227)(1466) 2331 --> (1466) 2331:PEGB1, pass, PUNB
			9'd231 : rdata = 43'b1100011100010000000000000000000001000000000;
			// PEs: 25 -> 32
			// srcs: (577, 228)(1504) 683 --> (1504) 683:PEGB1, pass, PUNB
			9'd232 : rdata = 43'b1100011100010000000000000000000001000000000;
			// PEs: 25 -> 32
			// srcs: (585, 232)(1618) 1450 --> (1618) 1450:PEGB1, pass, PUNB
			9'd233 : rdata = 43'b1100011100010000000000000000000001000000000;
			// PEs: 25 -> 32
			// srcs: (593, 233)(1637) 189 --> (1637) 189:PEGB1, pass, PUNB
			9'd234 : rdata = 43'b1100011100010000000000000000000001000000000;
			// PEs: 25 -> 32
			// srcs: (601, 234)(1656) 1475 --> (1656) 1475:PEGB1, pass, PUNB
			9'd235 : rdata = 43'b1100011100010000000000000000000001000000000;
			// PEs: 26 -> 32
			// srcs: (602, 235)(1675) 1935 --> (1675) 1935:PEGB2, pass, PUNB
			9'd236 : rdata = 43'b1100011100100000000000000000000001000000000;
			// PEs: 25 -> 32
			// srcs: (610, 243)(1279) 6449 --> (1279) 6449:PEGB1, pass, PUNB
			9'd237 : rdata = 43'b1100011100010000000000000000000001000000000;
			// PEs: 32 -> 25
			// srcs: (725, 237)(1695) 8048 --> (1695) 8048:PUGB4, pass, PENB
			9'd238 : rdata = 43'b1100011101001000000000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (732, 238)(1694) 840 --> (1694) 840:NI0, pass, PENB
			9'd239 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 16 -> 24
			// srcs: (733, 239)(1713) 2173 --> (1713) 2173:PUNB, pass, NI0
			9'd240 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 32 -> 25
			// srcs: (734, 240)(1714) 3029 --> (1714) 3029:PUGB4, pass, PENB
			9'd241 : rdata = 43'b1100011101001000000000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (740, 241)(1713) 2173 --> (1713) 2173:NI0, pass, PENB
			9'd242 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 16 -> 25
			// srcs: (741, 242)(1259) 3298 --> (1259) 3298:PUNB, pass, PENB
			9'd243 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 16 -> 25
			// srcs: (742, 244)(1696) 2251 --> (1696) 2251:PUNB, pass, PENB
			9'd244 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 16 -> 25
			// srcs: (743, 245)(1715) 3592 --> (1715) 3592:PUNB, pass, PENB
			9'd245 : rdata = 43'b1100011011111000000000000000000000100000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 25) begin
	always @(*) begin
		case(address)
			// PEs: 24 -> 
			// srcs: (14, 0)(654) 11 --> (654) 11:PENB, pass, 
			9'd0 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 24, 25 -> 24
			// srcs: (20, 1)(624) 84, (654) 11 --> (1224) 95:PENB, ALU, +, PEGB0
			9'd1 : rdata = 43'b0000111011110001111110000000000000010000000;
			// PEs: 24 -> 
			// srcs: (22, 2)(1194) 341 --> (1194) 341:PENB, pass, 
			9'd2 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 24, 25 -> 25
			// srcs: (28, 3)(1164) -9, (1194) 341 --> (1233) 332:PENB, ALU, +, NI0
			9'd3 : rdata = 43'b0000111011110001111111000000000000000000000;
			// PEs: 24 -> 
			// srcs: (30, 4)(655) 176 --> (655) 176:PENB, pass, 
			9'd4 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 24, 25 -> 25
			// srcs: (36, 5)(625) 560, (655) 176 --> (1243) 736:PENB, ALU, +, NI1
			9'd5 : rdata = 43'b0000111011110001111111000010000000000000000;
			// PEs: 24 -> 
			// srcs: (38, 6)(715) 1104 --> (715) 1104:PENB, pass, 
			9'd6 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 24, 25 -> 25
			// srcs: (44, 7)(685) 864, (715) 1104 --> (1244) 1968:PENB, ALU, +, NI2
			9'd7 : rdata = 43'b0000111011110001111111000100000000000000000;
			// PEs: 24 -> 25
			// srcs: (46, 8)(775) 551 --> (775) 551:PENB, pass, NI3
			9'd8 : rdata = 43'b1100011011110000000001000110000000000000000;
			// PEs: 25 -> 25
			// srcs: (47, 191)(1243) 736 --> (1243) 736:NI1, pass, NI1
			9'd9 : rdata = 43'b1100010100001000000001000010000000000000000;
			// PEs: 25, 25 -> 25
			// srcs: (47, 130)(1243) 736, (1244) 1968 --> (1253) 2704:ALU, NI2, +, NI4
			9'd10 : rdata = 43'b0000100111111101000101001000000000000000000;
			// PEs: 24, 25 -> 25
			// srcs: (52, 9)(745) 1008, (775) 551 --> (1245) 1559:PENB, NI3, +, NI1
			9'd11 : rdata = 43'b0000111011110101000111000010000000000000000;
			// PEs: 24 -> 
			// srcs: (54, 10)(1135) -39 --> (1135) -39:PENB, pass, 
			9'd12 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 24, 25 -> 25
			// srcs: (60, 11)(1105) 897, (1135) -39 --> (1251) 858:PENB, ALU, +, NI2
			9'd13 : rdata = 43'b0000111011110001111111000100000000000000000;
			// PEs: 24 -> 
			// srcs: (62, 12)(1195) 93 --> (1195) 93:PENB, pass, 
			9'd14 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 24, 25 -> 25
			// srcs: (68, 13)(1165) 117, (1195) 93 --> (1252) 210:PENB, ALU, +, NI3
			9'd15 : rdata = 43'b0000111011110001111111000110000000000000000;
			// PEs: 24 -> 25
			// srcs: (70, 14)(656) 121 --> (656) 121:PENB, pass, NI5
			9'd16 : rdata = 43'b1100011011110000000001001010000000000000000;
			// PEs: 25 -> 25
			// srcs: (71, 192)(1251) 858 --> (1251) 858:NI2, pass, NI2
			9'd17 : rdata = 43'b1100010100010000000001000100000000000000000;
			// PEs: 25, 25 -> 25
			// srcs: (71, 146)(1251) 858, (1252) 210 --> (1257) 1068:ALU, NI3, +, NI6
			9'd18 : rdata = 43'b0000100111111101000111001100000000000000000;
			// PEs: 24, 25 -> 25
			// srcs: (76, 15)(626) 364, (656) 121 --> (1262) 485:PENB, NI5, +, NI2
			9'd19 : rdata = 43'b0000111011110101001011000100000000000000000;
			// PEs: 24 -> 
			// srcs: (78, 16)(716) 644 --> (716) 644:PENB, pass, 
			9'd20 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 24, 25 -> 25
			// srcs: (84, 17)(686) 816, (716) 644 --> (1263) 1460:PENB, ALU, +, NI3
			9'd21 : rdata = 43'b0000111011110001111111000110000000000000000;
			// PEs: 24 -> 25
			// srcs: (86, 18)(776) 361 --> (776) 361:PENB, pass, NI5
			9'd22 : rdata = 43'b1100011011110000000001001010000000000000000;
			// PEs: 25 -> 25
			// srcs: (87, 193)(1262) 485 --> (1262) 485:NI2, pass, NI2
			9'd23 : rdata = 43'b1100010100010000000001000100000000000000000;
			// PEs: 25, 25 -> 25
			// srcs: (87, 132)(1262) 485, (1263) 1460 --> (1272) 1945:ALU, NI3, +, NI7
			9'd24 : rdata = 43'b0000100111111101000111001110000000000000000;
			// PEs: 24, 25 -> 25
			// srcs: (92, 19)(746) 792, (776) 361 --> (1264) 1153:PENB, NI5, +, NI2
			9'd25 : rdata = 43'b0000111011110101001011000100000000000000000;
			// PEs: 24 -> 
			// srcs: (94, 20)(836) 672 --> (836) 672:PENB, pass, 
			9'd26 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 24, 25 -> 25
			// srcs: (100, 21)(806) 372, (836) 672 --> (1265) 1044:PENB, ALU, +, NI3
			9'd27 : rdata = 43'b0000111011110001111111000110000000000000000;
			// PEs: 24 -> 25
			// srcs: (102, 22)(896) -5 --> (896) -5:PENB, pass, NI5
			9'd28 : rdata = 43'b1100011011110000000001001010000000000000000;
			// PEs: 25 -> 25
			// srcs: (103, 194)(1264) 1153 --> (1264) 1153:NI2, pass, NI2
			9'd29 : rdata = 43'b1100010100010000000001000100000000000000000;
			// PEs: 25, 25 -> 
			// srcs: (103, 133)(1264) 1153, (1265) 1044 --> (1273) 2197:ALU, NI3, +, 
			9'd30 : rdata = 43'b0000100111111101000110000000000000000000000;
			// PEs: 25, 25 -> 25
			// srcs: (106, 165)(1272) 1945, (1273) 2197 --> (1277) 4142:NI7, ALU, +, NI2
			9'd31 : rdata = 43'b0000110100111001111111000100000000000000000;
			// PEs: 24, 25 -> 24
			// srcs: (108, 23)(866) 416, (896) -5 --> (1266) 411:PENB, NI5, +, PEGB0
			9'd32 : rdata = 43'b0000111011110101001010000000000000010000000;
			// PEs: 24 -> 
			// srcs: (110, 24)(1076) 273 --> (1076) 273:PENB, pass, 
			9'd33 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 24, 25 -> 24
			// srcs: (116, 25)(1046) 1152, (1076) 273 --> (1269) 1425:PENB, ALU, +, PEGB0
			9'd34 : rdata = 43'b0000111011110001111110000000000000010000000;
			// PEs: 24 -> 
			// srcs: (118, 26)(1136) 468 --> (1136) 468:PENB, pass, 
			9'd35 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 24, 25 -> 25
			// srcs: (124, 27)(1106) 437, (1136) 468 --> (1270) 905:PENB, ALU, +, NI3
			9'd36 : rdata = 43'b0000111011110001111111000110000000000000000;
			// PEs: 24 -> 
			// srcs: (126, 28)(1196) 1240 --> (1196) 1240:PENB, pass, 
			9'd37 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 24, 25 -> 25
			// srcs: (132, 29)(1166) 162, (1196) 1240 --> (1271) 1402:PENB, ALU, +, NI5
			9'd38 : rdata = 43'b0000111011110001111111001010000000000000000;
			// PEs: 24 -> 25
			// srcs: (134, 30)(1138) 429 --> (1138) 429:PENB, pass, NI7
			9'd39 : rdata = 43'b1100011011110000000001001110000000000000000;
			// PEs: 25 -> 25
			// srcs: (135, 195)(1270) 905 --> (1270) 905:NI3, pass, NI3
			9'd40 : rdata = 43'b1100010100011000000001000110000000000000000;
			// PEs: 25, 25 -> 
			// srcs: (135, 147)(1270) 905, (1271) 1402 --> (1276) 2307:ALU, NI5, +, 
			9'd41 : rdata = 43'b0000100111111101001010000000000000000000000;
			// PEs: 25, 25 -> 25
			// srcs: (138, 171)(1276) 2307, (1277) 4142 --> (1279) 6449:ALU, NI2, +, NI3
			9'd42 : rdata = 43'b0000100111111101000101000110000000000000000;
			// PEs: 24, 25 -> 25
			// srcs: (140, 31)(1108) 1058, (1138) 429 --> (1308) 1487:PENB, NI7, +, NI2
			9'd43 : rdata = 43'b0000111011110101001111000100000000000000000;
			// PEs: 24 -> 
			// srcs: (142, 32)(1198) 1488 --> (1198) 1488:PENB, pass, 
			9'd44 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 24, 25 -> 25
			// srcs: (148, 33)(1168) 45, (1198) 1488 --> (1309) 1533:PENB, ALU, +, NI5
			9'd45 : rdata = 43'b0000111011110001111111001010000000000000000;
			// PEs: 24 -> 25
			// srcs: (150, 34)(1139) 143 --> (1139) 143:PENB, pass, NI7
			9'd46 : rdata = 43'b1100011011110000000001001110000000000000000;
			// PEs: 25 -> 25
			// srcs: (151, 196)(1308) 1487 --> (1308) 1487:NI2, pass, NI2
			9'd47 : rdata = 43'b1100010100010000000001000100000000000000000;
			// PEs: 25, 25 -> 25
			// srcs: (151, 148)(1308) 1487, (1309) 1533 --> (1314) 3020:ALU, NI5, +, NI8
			9'd48 : rdata = 43'b0000100111111101001011010000000000000000000;
			// PEs: 24, 25 -> 25
			// srcs: (156, 35)(1109) 46, (1139) 143 --> (1327) 189:PENB, NI7, +, NI2
			9'd49 : rdata = 43'b0000111011110101001111000100000000000000000;
			// PEs: 24 -> 
			// srcs: (158, 36)(1199) -62 --> (1199) -62:PENB, pass, 
			9'd50 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 24, 25 -> 25
			// srcs: (164, 37)(1169) 405, (1199) -62 --> (1328) 343:PENB, ALU, +, NI5
			9'd51 : rdata = 43'b0000111011110001111111001010000000000000000;
			// PEs: 24 -> 25
			// srcs: (166, 38)(1080) 483 --> (1080) 483:PENB, pass, NI7
			9'd52 : rdata = 43'b1100011011110000000001001110000000000000000;
			// PEs: 25 -> 25
			// srcs: (167, 197)(1327) 189 --> (1327) 189:NI2, pass, NI2
			9'd53 : rdata = 43'b1100010100010000000001000100000000000000000;
			// PEs: 25, 25 -> 24
			// srcs: (167, 149)(1327) 189, (1328) 343 --> (1333) 532:ALU, NI5, +, PEGB0
			9'd54 : rdata = 43'b0000100111111101001010000000000000010000000;
			// PEs: 24, 25 -> 24
			// srcs: (172, 39)(1050) 1332, (1080) 483 --> (1345) 1815:PENB, NI7, +, PEGB0
			9'd55 : rdata = 43'b0000111011110101001110000000000000010000000;
			// PEs: 24 -> 
			// srcs: (174, 40)(1140) 39 --> (1140) 39:PENB, pass, 
			9'd56 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 24, 25 -> 25
			// srcs: (180, 41)(1110) 391, (1140) 39 --> (1346) 430:PENB, ALU, +, NI2
			9'd57 : rdata = 43'b0000111011110001111111000100000000000000000;
			// PEs: 24 -> 
			// srcs: (182, 42)(1200) 434 --> (1200) 434:PENB, pass, 
			9'd58 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 24, 25 -> 25
			// srcs: (188, 43)(1170) -9, (1200) 434 --> (1347) 425:PENB, ALU, +, NI5
			9'd59 : rdata = 43'b0000111011110001111111001010000000000000000;
			// PEs: 24 -> 25
			// srcs: (190, 44)(661) 99 --> (661) 99:PENB, pass, NI7
			9'd60 : rdata = 43'b1100011011110000000001001110000000000000000;
			// PEs: 25 -> 25
			// srcs: (191, 198)(1346) 430 --> (1346) 430:NI2, pass, NI2
			9'd61 : rdata = 43'b1100010100010000000001000100000000000000000;
			// PEs: 25, 25 -> 25
			// srcs: (191, 150)(1346) 430, (1347) 425 --> (1352) 855:ALU, NI5, +, NI9
			9'd62 : rdata = 43'b0000100111111101001011010010000000000000000;
			// PEs: 24, 25 -> 25
			// srcs: (196, 45)(631) 28, (661) 99 --> (1357) 127:PENB, NI7, +, NI2
			9'd63 : rdata = 43'b0000111011110101001111000100000000000000000;
			// PEs: 24 -> 
			// srcs: (198, 46)(721) 506 --> (721) 506:PENB, pass, 
			9'd64 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 24, 25 -> 25
			// srcs: (204, 47)(691) 240, (721) 506 --> (1358) 746:PENB, ALU, +, NI5
			9'd65 : rdata = 43'b0000111011110001111111001010000000000000000;
			// PEs: 24 -> 25
			// srcs: (206, 48)(781) 114 --> (781) 114:PENB, pass, NI7
			9'd66 : rdata = 43'b1100011011110000000001001110000000000000000;
			// PEs: 25 -> 25
			// srcs: (207, 199)(1357) 127 --> (1357) 127:NI2, pass, NI2
			9'd67 : rdata = 43'b1100010100010000000001000100000000000000000;
			// PEs: 25, 25 -> 25
			// srcs: (207, 134)(1357) 127, (1358) 746 --> (1367) 873:ALU, NI5, +, NI10
			9'd68 : rdata = 43'b0000100111111101001011010100000000000000000;
			// PEs: 24, 25 -> 25
			// srcs: (212, 49)(751) 552, (781) 114 --> (1359) 666:PENB, NI7, +, NI2
			9'd69 : rdata = 43'b0000111011110101001111000100000000000000000;
			// PEs: 24 -> 
			// srcs: (214, 50)(1081) 231 --> (1081) 231:PENB, pass, 
			9'd70 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 24, 25 -> 25
			// srcs: (220, 51)(1051) 108, (1081) 231 --> (1364) 339:PENB, ALU, +, NI5
			9'd71 : rdata = 43'b0000111011110001111111001010000000000000000;
			// PEs: 24 -> 
			// srcs: (222, 52)(1141) 91 --> (1141) 91:PENB, pass, 
			9'd72 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 24, 25 -> 25
			// srcs: (228, 53)(1111) 437, (1141) 91 --> (1365) 528:PENB, ALU, +, NI7
			9'd73 : rdata = 43'b0000111011110001111111001110000000000000000;
			// PEs: 24 -> 
			// srcs: (230, 54)(1201) 186 --> (1201) 186:PENB, pass, 
			9'd74 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 24, 25 -> 25
			// srcs: (236, 55)(1171) 369, (1201) 186 --> (1366) 555:PENB, ALU, +, NI11
			9'd75 : rdata = 43'b0000111011110001111111010110000000000000000;
			// PEs: 24 -> 25
			// srcs: (238, 56)(1142) 91 --> (1142) 91:PENB, pass, NI12
			9'd76 : rdata = 43'b1100011011110000000001011000000000000000000;
			// PEs: 25 -> 25
			// srcs: (239, 200)(1365) 528 --> (1365) 528:NI7, pass, NI7
			9'd77 : rdata = 43'b1100010100111000000001001110000000000000000;
			// PEs: 25, 25 -> 25
			// srcs: (239, 151)(1365) 528, (1366) 555 --> (1371) 1083:ALU, NI11, +, NI13
			9'd78 : rdata = 43'b0000100111111101010111011010000000000000000;
			// PEs: 24, 25 -> 25
			// srcs: (244, 57)(1112) 161, (1142) 91 --> (1384) 252:PENB, NI12, +, NI7
			9'd79 : rdata = 43'b0000111011110101011001001110000000000000000;
			// PEs: 24 -> 
			// srcs: (246, 58)(1202) 1333 --> (1202) 1333:PENB, pass, 
			9'd80 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 24, 25 -> 25
			// srcs: (252, 59)(1172) 369, (1202) 1333 --> (1385) 1702:PENB, ALU, +, NI11
			9'd81 : rdata = 43'b0000111011110001111111010110000000000000000;
			// PEs: 24 -> 25
			// srcs: (254, 60)(1084) 525 --> (1084) 525:PENB, pass, NI12
			9'd82 : rdata = 43'b1100011011110000000001011000000000000000000;
			// PEs: 25 -> 25
			// srcs: (255, 201)(1384) 252 --> (1384) 252:NI7, pass, NI7
			9'd83 : rdata = 43'b1100010100111000000001001110000000000000000;
			// PEs: 25, 25 -> 25
			// srcs: (255, 152)(1384) 252, (1385) 1702 --> (1390) 1954:ALU, NI11, +, NI14
			9'd84 : rdata = 43'b0000100111111101010111011100000000000000000;
			// PEs: 24, 25 -> 25
			// srcs: (260, 61)(1054) 1188, (1084) 525 --> (1421) 1713:PENB, NI12, +, NI7
			9'd85 : rdata = 43'b0000111011110101011001001110000000000000000;
			// PEs: 24 -> 
			// srcs: (262, 62)(1144) 13 --> (1144) 13:PENB, pass, 
			9'd86 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 24, 25 -> 25
			// srcs: (268, 63)(1114) 483, (1144) 13 --> (1422) 496:PENB, ALU, +, NI11
			9'd87 : rdata = 43'b0000111011110001111111010110000000000000000;
			// PEs: 24 -> 
			// srcs: (270, 64)(1204) 1302 --> (1204) 1302:PENB, pass, 
			9'd88 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 24, 25 -> 25
			// srcs: (276, 65)(1174) 162, (1204) 1302 --> (1423) 1464:PENB, ALU, +, NI12
			9'd89 : rdata = 43'b0000111011110001111111011000000000000000000;
			// PEs: 24 -> 25
			// srcs: (278, 66)(726) 1242 --> (726) 1242:PENB, pass, NI15
			9'd90 : rdata = 43'b1100011011110000000001011110000000000000000;
			// PEs: 25 -> 25
			// srcs: (279, 202)(1422) 496 --> (1422) 496:NI11, pass, NI11
			9'd91 : rdata = 43'b1100010101011000000001010110000000000000000;
			// PEs: 25, 25 -> 25
			// srcs: (279, 153)(1422) 496, (1423) 1464 --> (1428) 1960:ALU, NI12, +, NI16
			9'd92 : rdata = 43'b0000100111111101011001100000000000000000000;
			// PEs: 24, 25 -> 24
			// srcs: (284, 67)(696) 792, (726) 1242 --> (1453) 2034:PENB, NI15, +, PEGB0
			9'd93 : rdata = 43'b0000111011110101011110000000000000010000000;
			// PEs: 24 -> 
			// srcs: (286, 68)(786) 266 --> (786) 266:PENB, pass, 
			9'd94 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 24, 25 -> 25
			// srcs: (292, 69)(756) 72, (786) 266 --> (1454) 338:PENB, ALU, +, NI11
			9'd95 : rdata = 43'b0000111011110001111111010110000000000000000;
			// PEs: 24 -> 
			// srcs: (294, 70)(1146) 195 --> (1146) 195:PENB, pass, 
			9'd96 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 24, 25 -> 25
			// srcs: (300, 71)(1116) 598, (1146) 195 --> (1460) 793:PENB, ALU, +, NI12
			9'd97 : rdata = 43'b0000111011110001111111011000000000000000000;
			// PEs: 24 -> 
			// srcs: (302, 72)(1206) 1178 --> (1206) 1178:PENB, pass, 
			9'd98 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 24, 25 -> 25
			// srcs: (308, 73)(1176) 360, (1206) 1178 --> (1461) 1538:PENB, ALU, +, NI15
			9'd99 : rdata = 43'b0000111011110001111111011110000000000000000;
			// PEs: 24 -> 25
			// srcs: (310, 74)(667) 0 --> (667) 0:PENB, pass, NI17
			9'd100 : rdata = 43'b1100011011110000000001100010000000000000000;
			// PEs: 25 -> 25
			// srcs: (311, 203)(1460) 793 --> (1460) 793:NI12, pass, NI12
			9'd101 : rdata = 43'b1100010101100000000001011000000000000000000;
			// PEs: 25, 25 -> 25
			// srcs: (311, 154)(1460) 793, (1461) 1538 --> (1466) 2331:ALU, NI15, +, NI18
			9'd102 : rdata = 43'b0000100111111101011111100100000000000000000;
			// PEs: 24, 25 -> 25
			// srcs: (316, 75)(637) 84, (667) 0 --> (1471) 84:PENB, NI17, +, NI12
			9'd103 : rdata = 43'b0000111011110101100011011000000000000000000;
			// PEs: 24 -> 
			// srcs: (318, 76)(727) 184 --> (727) 184:PENB, pass, 
			9'd104 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 24, 25 -> 25
			// srcs: (324, 77)(697) 1176, (727) 184 --> (1472) 1360:PENB, ALU, +, NI15
			9'd105 : rdata = 43'b0000111011110001111111011110000000000000000;
			// PEs: 24 -> 25
			// srcs: (326, 78)(787) 741 --> (787) 741:PENB, pass, NI17
			9'd106 : rdata = 43'b1100011011110000000001100010000000000000000;
			// PEs: 25 -> 25
			// srcs: (327, 204)(1471) 84 --> (1471) 84:NI12, pass, NI12
			9'd107 : rdata = 43'b1100010101100000000001011000000000000000000;
			// PEs: 25, 25 -> 25
			// srcs: (327, 139)(1471) 84, (1472) 1360 --> (1481) 1444:ALU, NI15, +, NI19
			9'd108 : rdata = 43'b0000100111111101011111100110000000000000000;
			// PEs: 24, 25 -> 25
			// srcs: (332, 79)(757) 888, (787) 741 --> (1473) 1629:PENB, NI17, +, NI12
			9'd109 : rdata = 43'b0000111011110101100011011000000000000000000;
			// PEs: 24 -> 
			// srcs: (334, 80)(1087) 903 --> (1087) 903:PENB, pass, 
			9'd110 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 24, 25 -> 25
			// srcs: (340, 81)(1057) 1080, (1087) 903 --> (1478) 1983:PENB, ALU, +, NI15
			9'd111 : rdata = 43'b0000111011110001111111011110000000000000000;
			// PEs: 24 -> 
			// srcs: (342, 82)(1147) 377 --> (1147) 377:PENB, pass, 
			9'd112 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 24, 25 -> 25
			// srcs: (348, 83)(1117) 1035, (1147) 377 --> (1479) 1412:PENB, ALU, +, NI17
			9'd113 : rdata = 43'b0000111011110001111111100010000000000000000;
			// PEs: 24 -> 
			// srcs: (350, 84)(1207) 372 --> (1207) 372:PENB, pass, 
			9'd114 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 24, 25 -> 25
			// srcs: (356, 85)(1177) 396, (1207) 372 --> (1480) 768:PENB, ALU, +, NI20
			9'd115 : rdata = 43'b0000111011110001111111101000000000000000000;
			// PEs: 24 -> 25
			// srcs: (358, 86)(1148) 273 --> (1148) 273:PENB, pass, NI21
			9'd116 : rdata = 43'b1100011011110000000001101010000000000000000;
			// PEs: 25 -> 25
			// srcs: (359, 205)(1479) 1412 --> (1479) 1412:NI17, pass, NI17
			9'd117 : rdata = 43'b1100010110001000000001100010000000000000000;
			// PEs: 25, 25 -> 25
			// srcs: (359, 155)(1479) 1412, (1480) 768 --> (1485) 2180:ALU, NI20, +, NI22
			9'd118 : rdata = 43'b0000100111111101101001101100000000000000000;
			// PEs: 24, 25 -> 25
			// srcs: (364, 87)(1118) 391, (1148) 273 --> (1498) 664:PENB, NI21, +, NI17
			9'd119 : rdata = 43'b0000111011110101101011100010000000000000000;
			// PEs: 24 -> 
			// srcs: (366, 88)(1208) -62 --> (1208) -62:PENB, pass, 
			9'd120 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 24, 25 -> 25
			// srcs: (372, 89)(1178) 81, (1208) -62 --> (1499) 19:PENB, ALU, +, NI20
			9'd121 : rdata = 43'b0000111011110001111111101000000000000000000;
			// PEs: 24 -> 25
			// srcs: (374, 90)(669) 187 --> (669) 187:PENB, pass, NI21
			9'd122 : rdata = 43'b1100011011110000000001101010000000000000000;
			// PEs: 25 -> 25
			// srcs: (375, 206)(1498) 664 --> (1498) 664:NI17, pass, NI17
			9'd123 : rdata = 43'b1100010110001000000001100010000000000000000;
			// PEs: 25, 25 -> 25
			// srcs: (375, 156)(1498) 664, (1499) 19 --> (1504) 683:ALU, NI20, +, NI23
			9'd124 : rdata = 43'b0000100111111101101001101110000000000000000;
			// PEs: 24, 25 -> 25
			// srcs: (380, 91)(639) 56, (669) 187 --> (1509) 243:PENB, NI21, +, NI17
			9'd125 : rdata = 43'b0000111011110101101011100010000000000000000;
			// PEs: 24 -> 
			// srcs: (382, 92)(729) 1472 --> (729) 1472:PENB, pass, 
			9'd126 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 24, 25 -> 25
			// srcs: (388, 93)(699) 408, (729) 1472 --> (1510) 1880:PENB, ALU, +, NI20
			9'd127 : rdata = 43'b0000111011110001111111101000000000000000000;
			// PEs: 24 -> 25
			// srcs: (390, 94)(789) 532 --> (789) 532:PENB, pass, NI21
			9'd128 : rdata = 43'b1100011011110000000001101010000000000000000;
			// PEs: 25 -> 25
			// srcs: (391, 207)(1509) 243 --> (1509) 243:NI17, pass, NI17
			9'd129 : rdata = 43'b1100010110001000000001100010000000000000000;
			// PEs: 25, 25 -> 25
			// srcs: (391, 142)(1509) 243, (1510) 1880 --> (1519) 2123:ALU, NI20, +, NI24
			9'd130 : rdata = 43'b0000100111111101101001110000000000000000000;
			// PEs: 24, 25 -> 24
			// srcs: (396, 95)(759) 840, (789) 532 --> (1511) 1372:PENB, NI21, +, PEGB0
			9'd131 : rdata = 43'b0000111011110101101010000000000000010000000;
			// PEs: 24 -> 
			// srcs: (398, 96)(1149) 429 --> (1149) 429:PENB, pass, 
			9'd132 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 24, 25 -> 25
			// srcs: (404, 97)(1119) 322, (1149) 429 --> (1517) 751:PENB, ALU, +, NI17
			9'd133 : rdata = 43'b0000111011110001111111100010000000000000000;
			// PEs: 24 -> 
			// srcs: (406, 98)(1209) 806 --> (1209) 806:PENB, pass, 
			9'd134 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 24, 25 -> 25
			// srcs: (412, 99)(1179) 333, (1209) 806 --> (1518) 1139:PENB, ALU, +, NI20
			9'd135 : rdata = 43'b0000111011110001111111101000000000000000000;
			// PEs: 24 -> 25
			// srcs: (414, 100)(1090) 588 --> (1090) 588:PENB, pass, NI21
			9'd136 : rdata = 43'b1100011011110000000001101010000000000000000;
			// PEs: 25 -> 25
			// srcs: (415, 208)(1517) 751 --> (1517) 751:NI17, pass, NI17
			9'd137 : rdata = 43'b1100010110001000000001100010000000000000000;
			// PEs: 25, 25 -> 24
			// srcs: (415, 157)(1517) 751, (1518) 1139 --> (1523) 1890:ALU, NI20, +, PEGB0
			9'd138 : rdata = 43'b0000100111111101101000000000000000010000000;
			// PEs: 24, 25 -> 24
			// srcs: (420, 101)(1060) 720, (1090) 588 --> (1535) 1308:PENB, NI21, +, PEGB0
			9'd139 : rdata = 43'b0000111011110101101010000000000000010000000;
			// PEs: 24 -> 
			// srcs: (422, 102)(1150) 559 --> (1150) 559:PENB, pass, 
			9'd140 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 24, 25 -> 25
			// srcs: (428, 103)(1120) 437, (1150) 559 --> (1536) 996:PENB, ALU, +, NI17
			9'd141 : rdata = 43'b0000111011110001111111100010000000000000000;
			// PEs: 24 -> 
			// srcs: (430, 104)(1210) 1209 --> (1210) 1209:PENB, pass, 
			9'd142 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 24, 25 -> 25
			// srcs: (436, 105)(1180) 261, (1210) 1209 --> (1537) 1470:PENB, ALU, +, NI20
			9'd143 : rdata = 43'b0000111011110001111111101000000000000000000;
			// PEs: 24 -> 25
			// srcs: (438, 106)(1092) 672 --> (1092) 672:PENB, pass, NI21
			9'd144 : rdata = 43'b1100011011110000000001101010000000000000000;
			// PEs: 25 -> 25
			// srcs: (439, 209)(1536) 996 --> (1536) 996:NI17, pass, NI17
			9'd145 : rdata = 43'b1100010110001000000001100010000000000000000;
			// PEs: 25, 25 -> 24
			// srcs: (439, 158)(1536) 996, (1537) 1470 --> (1542) 2466:ALU, NI20, +, PEGB0
			9'd146 : rdata = 43'b0000100111111101101000000000000000010000000;
			// PEs: 24, 25 -> 24
			// srcs: (444, 107)(1062) 612, (1092) 672 --> (1573) 1284:PENB, NI21, +, PEGB0
			9'd147 : rdata = 43'b0000111011110101101010000000000000010000000;
			// PEs: 24 -> 
			// srcs: (446, 108)(1152) 312 --> (1152) 312:PENB, pass, 
			9'd148 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 24, 25 -> 25
			// srcs: (452, 109)(1122) 920, (1152) 312 --> (1574) 1232:PENB, ALU, +, NI17
			9'd149 : rdata = 43'b0000111011110001111111100010000000000000000;
			// PEs: 24 -> 
			// srcs: (454, 110)(1212) 1085 --> (1212) 1085:PENB, pass, 
			9'd150 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 24, 25 -> 25
			// srcs: (460, 111)(1182) 297, (1212) 1085 --> (1575) 1382:PENB, ALU, +, NI20
			9'd151 : rdata = 43'b0000111011110001111111101000000000000000000;
			// PEs: 24 -> 25
			// srcs: (462, 112)(1154) 273 --> (1154) 273:PENB, pass, NI21
			9'd152 : rdata = 43'b1100011011110000000001101010000000000000000;
			// PEs: 25 -> 25
			// srcs: (463, 210)(1574) 1232 --> (1574) 1232:NI17, pass, NI17
			9'd153 : rdata = 43'b1100010110001000000001100010000000000000000;
			// PEs: 25, 25 -> 24
			// srcs: (463, 159)(1574) 1232, (1575) 1382 --> (1580) 2614:ALU, NI20, +, PEGB0
			9'd154 : rdata = 43'b0000100111111101101000000000000000010000000;
			// PEs: 24, 25 -> 25
			// srcs: (468, 113)(1124) 1127, (1154) 273 --> (1612) 1400:PENB, NI21, +, NI17
			9'd155 : rdata = 43'b0000111011110101101011100010000000000000000;
			// PEs: 24 -> 
			// srcs: (470, 114)(1214) -31 --> (1214) -31:PENB, pass, 
			9'd156 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 24, 25 -> 25
			// srcs: (476, 115)(1184) 81, (1214) -31 --> (1613) 50:PENB, ALU, +, NI20
			9'd157 : rdata = 43'b0000111011110001111111101000000000000000000;
			// PEs: 24 -> 25
			// srcs: (478, 116)(1095) 609 --> (1095) 609:PENB, pass, NI21
			9'd158 : rdata = 43'b1100011011110000000001101010000000000000000;
			// PEs: 25 -> 25
			// srcs: (479, 211)(1612) 1400 --> (1612) 1400:NI17, pass, NI17
			9'd159 : rdata = 43'b1100010110001000000001100010000000000000000;
			// PEs: 25, 25 -> 25
			// srcs: (479, 160)(1612) 1400, (1613) 50 --> (1618) 1450:ALU, NI20, +, NI25
			9'd160 : rdata = 43'b0000100111111101101001110010000000000000000;
			// PEs: 24, 25 -> 24
			// srcs: (484, 117)(1065) 864, (1095) 609 --> (1630) 1473:PENB, NI21, +, PEGB0
			9'd161 : rdata = 43'b0000111011110101101010000000000000010000000;
			// PEs: 24 -> 
			// srcs: (486, 118)(1155) 0 --> (1155) 0:PENB, pass, 
			9'd162 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 24, 25 -> 25
			// srcs: (492, 119)(1125) 138, (1155) 0 --> (1631) 138:PENB, ALU, +, NI17
			9'd163 : rdata = 43'b0000111011110001111111100010000000000000000;
			// PEs: 24 -> 25
			// srcs: (494, 120)(1215) -93 --> (1215) -93:PENB, pass, NI20
			9'd164 : rdata = 43'b1100011011110000000001101000000000000000000;
			// PEs: 25 -> 24
			// srcs: (495, 172)(1314) 3020 --> (1314) 3020:NI8, pass, PEGB0
			9'd165 : rdata = 43'b1100010101000000000000000000000000010000000;
			// PEs: 24, 25 -> 25
			// srcs: (500, 121)(1185) 144, (1215) -93 --> (1632) 51:PENB, NI20, +, NI8
			9'd166 : rdata = 43'b0000111011110101101001010000000000000000000;
			// PEs: 24 -> 25
			// srcs: (502, 122)(1156) 39 --> (1156) 39:PENB, pass, NI20
			9'd167 : rdata = 43'b1100011011110000000001101000000000000000000;
			// PEs: 25 -> 25
			// srcs: (503, 212)(1631) 138 --> (1631) 138:NI17, pass, NI17
			9'd168 : rdata = 43'b1100010110001000000001100010000000000000000;
			// PEs: 25, 25 -> 25
			// srcs: (503, 161)(1631) 138, (1632) 51 --> (1637) 189:ALU, NI8, +, NI21
			9'd169 : rdata = 43'b0000100111111101010001101010000000000000000;
			// PEs: 25 -> 24
			// srcs: (504, 175)(1390) 1954 --> (1390) 1954:NI14, pass, PEGB0
			9'd170 : rdata = 43'b1100010101110000000000000000000000010000000;
			// PEs: 24, 25 -> 25
			// srcs: (508, 123)(1126) 897, (1156) 39 --> (1650) 936:PENB, NI20, +, NI8
			9'd171 : rdata = 43'b0000111011110101101001010000000000000000000;
			// PEs: 24 -> 25
			// srcs: (510, 124)(1216) 341 --> (1216) 341:PENB, pass, NI14
			9'd172 : rdata = 43'b1100011011110000000001011100000000000000000;
			// PEs: 25 -> 24
			// srcs: (512, 176)(1428) 1960 --> (1428) 1960:NI16, pass, PEGB0
			9'd173 : rdata = 43'b1100010110000000000000000000000000010000000;
			// PEs: 24, 25 -> 25
			// srcs: (516, 125)(1186) 198, (1216) 341 --> (1651) 539:PENB, NI14, +, NI16
			9'd174 : rdata = 43'b0000111011110101011101100000000000000000000;
			// PEs: 24 -> 25
			// srcs: (518, 126)(1157) 195 --> (1157) 195:PENB, pass, NI14
			9'd175 : rdata = 43'b1100011011110000000001011100000000000000000;
			// PEs: 25 -> 25
			// srcs: (519, 213)(1650) 936 --> (1650) 936:NI8, pass, NI8
			9'd176 : rdata = 43'b1100010101000000000001010000000000000000000;
			// PEs: 25, 25 -> 25
			// srcs: (519, 162)(1650) 936, (1651) 539 --> (1656) 1475:ALU, NI16, +, NI17
			9'd177 : rdata = 43'b0000100111111101100001100010000000000000000;
			// PEs: 24, 25 -> 25
			// srcs: (524, 127)(1127) 989, (1157) 195 --> (1669) 1184:PENB, NI14, +, NI8
			9'd178 : rdata = 43'b0000111011110101011101010000000000000000000;
			// PEs: 24 -> 
			// srcs: (526, 128)(1217) 310 --> (1217) 310:PENB, pass, 
			9'd179 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 24, 25 -> 26
			// srcs: (532, 129)(1187) 441, (1217) 310 --> (1670) 751:PENB, ALU, +, PENB
			9'd180 : rdata = 43'b0000111011110001111110000000000000100000000;
			// PEs: 25, 24 -> 26
			// srcs: (533, 131)(1245) 1559, (1246) 962 --> (1254) 2521:NI1, PENB, +, PENB
			9'd181 : rdata = 43'b0000110100001110111100000000000000100000000;
			// PEs: 25, 24 -> 26
			// srcs: (534, 135)(1359) 666, (1360) 183 --> (1368) 849:NI2, PENB, +, PENB
			9'd182 : rdata = 43'b0000110100010110111100000000000000100000000;
			// PEs: 24, 25 -> 27
			// srcs: (535, 136)(1363) 930, (1364) 339 --> (1370) 1269:PENB, NI5, +, PEGB3
			9'd183 : rdata = 43'b0000111011110101001010000000000000010110000;
			// PEs: 24, 25 -> 24
			// srcs: (536, 137)(1420) 858, (1421) 1713 --> (1427) 2571:PENB, NI7, +, PEGB0
			9'd184 : rdata = 43'b0000111011110101001110000000000000010000000;
			// PEs: 25, 24 -> 24
			// srcs: (537, 138)(1454) 338, (1455) 789 --> (1463) 1127:NI11, PENB, +, PEGB0
			9'd185 : rdata = 43'b0000110101011110111100000000000000010000000;
			// PEs: 25, 24 -> 26
			// srcs: (538, 140)(1473) 1629, (1474) 1940 --> (1482) 3569:NI12, PENB, +, PENB
			9'd186 : rdata = 43'b0000110101100110111100000000000000100000000;
			// PEs: 24, 25 -> 25
			// srcs: (539, 141)(1477) 870, (1478) 1983 --> (1484) 2853:PENB, NI15, +, NI1
			9'd187 : rdata = 43'b0000111011110101011111000010000000000000000;
			// PEs: 25 -> 26
			// srcs: (540, 163)(1669) 1184 --> (1669) 1184:NI8, pass, PENB
			9'd188 : rdata = 43'b1100010101000000000000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (541, 143)(1702) 1312 --> (1702) 1312:PENB, pass, NI2
			9'd189 : rdata = 43'b1100011011110000000001000100000000000000000;
			// PEs: 25 -> 26
			// srcs: (542, 164)(1253) 2704 --> (1253) 2704:NI4, pass, PENB
			9'd190 : rdata = 43'b1100010100100000000000000000000000100000000;
			// PEs: 25 -> 26
			// srcs: (543, 166)(1367) 873 --> (1367) 873:NI10, pass, PENB
			9'd191 : rdata = 43'b1100010101010000000000000000000000100000000;
			// PEs: 25 -> 26
			// srcs: (545, 167)(1481) 1444 --> (1481) 1444:NI19, pass, PENB
			9'd192 : rdata = 43'b1100010110011000000000000000000000100000000;
			// PEs: 25 -> 24
			// srcs: (546, 168)(1519) 2123 --> (1519) 2123:NI24, pass, PEGB0
			9'd193 : rdata = 43'b1100010111000000000000000000000000010000000;
			// PEs: 24, 25 -> 24
			// srcs: (547, 144)(1701) 1049, (1702) 1312 --> (1710) 2361:PENB, NI2, +, PEGB0
			9'd194 : rdata = 43'b0000111011110101000100000000000000010000000;
			// PEs: 24, 25 -> 24
			// srcs: (548, 145)(1232) 613, (1233) 332 --> (1238) 945:PENB, NI0, +, PEGB0
			9'd195 : rdata = 43'b0000111011110101000000000000000000010000000;
			// PEs: 25, 26 -> 25
			// srcs: (550, 170)(1257) 1068, (1258) 5225 --> (1260) 6293:NI6, PEGB2, +, NI0
			9'd196 : rdata = 43'b0000110100110111001001000000000000000000000;
			// PEs: 25 -> 26
			// srcs: (551, 174)(1371) 1083 --> (1371) 1083:NI13, pass, PENB
			9'd197 : rdata = 43'b1100010101101000000000000000000000100000000;
			// PEs: 25 -> 26
			// srcs: (552, 178)(1485) 2180 --> (1485) 2180:NI22, pass, PENB
			9'd198 : rdata = 43'b1100010110110000000000000000000000100000000;
			// PEs: 25 -> 26
			// srcs: (555, 169)(1484) 2853 --> (1484) 2853:NI1, pass, PENB
			9'd199 : rdata = 43'b1100010100001000000000000000000000100000000;
			// PEs: 25 -> 24
			// srcs: (556, 173)(1352) 855 --> (1352) 855:NI9, pass, PEGB0
			9'd200 : rdata = 43'b1100010101001000000000000000000000010000000;
			// PEs: 25 -> 24
			// srcs: (564, 177)(1466) 2331 --> (1466) 2331:NI18, pass, PEGB0
			9'd201 : rdata = 43'b1100010110010000000000000000000000010000000;
			// PEs: 25 -> 24
			// srcs: (572, 179)(1504) 683 --> (1504) 683:NI23, pass, PEGB0
			9'd202 : rdata = 43'b1100010110111000000000000000000000010000000;
			// PEs: 25 -> 24
			// srcs: (580, 180)(1618) 1450 --> (1618) 1450:NI25, pass, PEGB0
			9'd203 : rdata = 43'b1100010111001000000000000000000000010000000;
			// PEs: 25 -> 24
			// srcs: (588, 181)(1637) 189 --> (1637) 189:NI21, pass, PEGB0
			9'd204 : rdata = 43'b1100010110101000000000000000000000010000000;
			// PEs: 25 -> 24
			// srcs: (596, 182)(1656) 1475 --> (1656) 1475:NI17, pass, PEGB0
			9'd205 : rdata = 43'b1100010110001000000000000000000000010000000;
			// PEs: 25 -> 24
			// srcs: (605, 188)(1279) 6449 --> (1279) 6449:NI3, pass, PEGB0
			9'd206 : rdata = 43'b1100010100011000000000000000000000010000000;
			// PEs: 24 -> 
			// srcs: (727, 183)(1695) 8048 --> (1695) 8048:PENB, pass, 
			9'd207 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 24, 25 -> 25
			// srcs: (734, 184)(1694) 840, (1695) 8048 --> (1697) 8888:PENB, ALU, +, NI1
			9'd208 : rdata = 43'b0000111011110001111111000010000000000000000;
			// PEs: 24 -> 
			// srcs: (736, 185)(1714) 3029 --> (1714) 3029:PENB, pass, 
			9'd209 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 24, 25 -> 25
			// srcs: (742, 186)(1713) 2173, (1714) 3029 --> (1716) 5202:PENB, ALU, +, NI2
			9'd210 : rdata = 43'b0000111011110001111111000100000000000000000;
			// PEs: 24, 25 -> 25
			// srcs: (743, 187)(1259) 3298, (1260) 6293 --> (1261) 9591:PENB, NI0, +, NW0
			9'd211 : rdata = 43'b0000111011110101000000000001000000000000000;
			// PEs: 24, 25 -> 25
			// srcs: (744, 189)(1696) 2251, (1697) 8888 --> (1698) 11139:PENB, NI1, +, NW1
			9'd212 : rdata = 43'b0000111011110101000010000001000010000000000;
			// PEs: 24, 25 -> 25
			// srcs: (752, 190)(1715) 3592, (1716) 5202 --> (1717) 8794:PENB, NI2, +, NW2
			9'd213 : rdata = 43'b0000111011110101000100000001000100000000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 26) begin
	always @(*) begin
		case(address)
			// PEs: 25 -> 26
			// srcs: (534, 0)(1670) 751 --> (1670) 751:PENB, pass, NI0
			9'd0 : rdata = 43'b1100011011110000000001000000000000000000000;
			// PEs: 25 -> 26
			// srcs: (535, 2)(1254) 2521 --> (1254) 2521:PENB, pass, NI1
			9'd1 : rdata = 43'b1100011011110000000001000010000000000000000;
			// PEs: 25 -> 26
			// srcs: (536, 4)(1368) 849 --> (1368) 849:PENB, pass, NI2
			9'd2 : rdata = 43'b1100011011110000000001000100000000000000000;
			// PEs: 25 -> 26
			// srcs: (540, 6)(1482) 3569 --> (1482) 3569:PENB, pass, NI3
			9'd3 : rdata = 43'b1100011011110000000001000110000000000000000;
			// PEs: 25, 26 -> 24
			// srcs: (542, 1)(1669) 1184, (1670) 751 --> (1675) 1935:PENB, NI0, +, PEGB0
			9'd4 : rdata = 43'b0000111011110101000000000000000000010000000;
			// PEs: 25, 26 -> 25
			// srcs: (544, 3)(1253) 2704, (1254) 2521 --> (1258) 5225:PENB, NI1, +, PEGB1
			9'd5 : rdata = 43'b0000111011110101000010000000000000010010000;
			// PEs: 25, 26 -> 26
			// srcs: (545, 5)(1367) 873, (1368) 849 --> (1372) 1722:PENB, NI2, +, NI0
			9'd6 : rdata = 43'b0000111011110101000101000000000000000000000;
			// PEs: 25, 26 -> 26
			// srcs: (547, 7)(1481) 1444, (1482) 3569 --> (1486) 5013:PENB, NI3, +, NI1
			9'd7 : rdata = 43'b0000111011110101000111000010000000000000000;
			// PEs: 25, 26 -> 27
			// srcs: (553, 9)(1371) 1083, (1372) 1722 --> (1374) 2805:PENB, NI0, +, PENB
			9'd8 : rdata = 43'b0000111011110101000000000000000000100000000;
			// PEs: 25, 26 -> 26
			// srcs: (554, 10)(1485) 2180, (1486) 5013 --> (1488) 7193:PENB, NI1, +, NI0
			9'd9 : rdata = 43'b0000111011110101000011000000000000000000000;
			// PEs: 24, 25 -> 
			// srcs: (557, 8)(1483) 3047, (1484) 2853 --> (1487) 5900:PEGB0, PENB, +, 
			9'd10 : rdata = 43'b0000111100000110111100000000000000000000000;
			// PEs: 26, 26 -> 26
			// srcs: (560, 11)(1487) 5900, (1488) 7193 --> (1489) 13093:ALU, NI0, +, NW0
			9'd11 : rdata = 43'b0000100111111101000000000001000000000000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 27) begin
	always @(*) begin
		case(address)
			// PEs: 24 -> 
			// srcs: (552, 0)(1369) 1708 --> (1369) 1708:PEGB0, pass, 
			9'd0 : rdata = 43'b1100011100000000000000000000000000000000000;
			// PEs: 27, 25 -> 
			// srcs: (554, 1)(1369) 1708, (1370) 1269 --> (1373) 2977:ALU, PEGB1, +, 
			9'd1 : rdata = 43'b0000100111111111000100000000000000000000000;
			// PEs: 27, 26 -> 27
			// srcs: (557, 2)(1373) 2977, (1374) 2805 --> (1375) 5782:ALU, PENB, +, NW0
			9'd2 : rdata = 43'b0000100111111110111100000001000000000000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 28) begin
	always @(*) begin
		case(address)
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 29) begin
	always @(*) begin
		case(address)
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 30) begin
	always @(*) begin
		case(address)
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 31) begin
	always @(*) begin
		case(address)
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 32) begin
	always @(*) begin
		case(address)
			// PEs: 0 -> 32
			// srcs: (13, 0)(684) 1032 --> (684) 1032:PUGB0, pass, NI0
			9'd0 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 0 -> 33
			// srcs: (14, 1)(714) 2116 --> (714) 2116:PUGB0, pass, PENB
			9'd1 : rdata = 43'b1100011100001000000000000000000000100000000;
			// PEs: 32 -> 33
			// srcs: (20, 2)(684) 1032 --> (684) 1032:NI0, pass, PENB
			9'd2 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 32
			// srcs: (21, 3)(744) 120 --> (744) 120:PUGB0, pass, NI0
			9'd3 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 0 -> 33
			// srcs: (22, 4)(774) 722 --> (774) 722:PUGB0, pass, PENB
			9'd4 : rdata = 43'b1100011100001000000000000000000000100000000;
			// PEs: 33 -> 48
			// srcs: (27, 99)(1225) 3148 --> (1225) 3148:PEGB1, pass, PUGB6
			9'd5 : rdata = 43'b1100011100010000000000000000000000000001110;
			// PEs: 32 -> 33
			// srcs: (28, 5)(744) 120 --> (744) 120:NI0, pass, PENB
			9'd6 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 8 -> 32
			// srcs: (29, 6)(864) 1216 --> (864) 1216:PUGB1, pass, NI0
			9'd7 : rdata = 43'b1100011100011000000001000000000000000000000;
			// PEs: 8 -> 33
			// srcs: (30, 7)(894) -22 --> (894) -22:PUGB1, pass, PENB
			9'd8 : rdata = 43'b1100011100011000000000000000000000100000000;
			// PEs: 33 -> 40
			// srcs: (35, 100)(1226) 842 --> (1226) 842:PEGB1, pass, PUNB
			9'd9 : rdata = 43'b1100011100010000000000000000000001000000000;
			// PEs: 32 -> 33
			// srcs: (36, 8)(864) 1216 --> (864) 1216:NI0, pass, PENB
			9'd10 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 8 -> 32
			// srcs: (37, 9)(924) 667 --> (924) 667:PUGB1, pass, NI0
			9'd11 : rdata = 43'b1100011100011000000001000000000000000000000;
			// PEs: 8 -> 33
			// srcs: (38, 10)(954) 1551 --> (954) 1551:PUGB1, pass, PENB
			9'd12 : rdata = 43'b1100011100011000000000000000000000100000000;
			// PEs: 32 -> 33
			// srcs: (44, 11)(924) 667 --> (924) 667:NI0, pass, PENB
			9'd13 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 8 -> 32
			// srcs: (45, 12)(984) 92 --> (984) 92:PUGB1, pass, NI0
			9'd14 : rdata = 43'b1100011100011000000001000000000000000000000;
			// PEs: 8 -> 33
			// srcs: (46, 13)(1014) 462 --> (1014) 462:PUGB1, pass, PENB
			9'd15 : rdata = 43'b1100011100011000000000000000000000100000000;
			// PEs: 32 -> 33
			// srcs: (52, 14)(984) 92 --> (984) 92:NI0, pass, PENB
			9'd16 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 32
			// srcs: (53, 15)(627) 238 --> (627) 238:PUGB0, pass, NI0
			9'd17 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 0 -> 33
			// srcs: (54, 16)(657) 66 --> (657) 66:PUGB0, pass, PENB
			9'd18 : rdata = 43'b1100011100001000000000000000000000100000000;
			// PEs: 33 -> 40
			// srcs: (59, 101)(1230) 554 --> (1230) 554:PEGB1, pass, PUNB
			9'd19 : rdata = 43'b1100011100010000000000000000000001000000000;
			// PEs: 32 -> 33
			// srcs: (60, 17)(627) 238 --> (627) 238:NI0, pass, PENB
			9'd20 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 32
			// srcs: (61, 18)(687) 168 --> (687) 168:PUGB0, pass, NI0
			9'd21 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 0 -> 33
			// srcs: (62, 19)(717) 598 --> (717) 598:PUGB0, pass, PENB
			9'd22 : rdata = 43'b1100011100001000000000000000000000100000000;
			// PEs: 32 -> 33
			// srcs: (68, 20)(687) 168 --> (687) 168:NI0, pass, PENB
			9'd23 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 32
			// srcs: (69, 21)(747) 864 --> (747) 864:PUGB0, pass, NI0
			9'd24 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 0 -> 33
			// srcs: (70, 22)(777) 703 --> (777) 703:PUGB0, pass, PENB
			9'd25 : rdata = 43'b1100011100001000000000000000000000100000000;
			// PEs: 32 -> 33
			// srcs: (76, 23)(747) 864 --> (747) 864:NI0, pass, PENB
			9'd26 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 32
			// srcs: (77, 24)(630) 252 --> (630) 252:PUGB0, pass, NI0
			9'd27 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 0 -> 33
			// srcs: (78, 25)(660) -22 --> (660) -22:PUGB0, pass, PENB
			9'd28 : rdata = 43'b1100011100001000000000000000000000100000000;
			// PEs: 33 -> 40
			// srcs: (83, 102)(1283) 1567 --> (1283) 1567:PEGB1, pass, PUNB
			9'd29 : rdata = 43'b1100011100010000000000000000000001000000000;
			// PEs: 32 -> 33
			// srcs: (84, 26)(630) 252 --> (630) 252:NI0, pass, PENB
			9'd30 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 32
			// srcs: (85, 27)(690) 192 --> (690) 192:PUGB0, pass, NI0
			9'd31 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 0 -> 33
			// srcs: (86, 28)(720) 1288 --> (720) 1288:PUGB0, pass, PENB
			9'd32 : rdata = 43'b1100011100001000000000000000000000100000000;
			// PEs: 32 -> 33
			// srcs: (92, 29)(690) 192 --> (690) 192:NI0, pass, PENB
			9'd33 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 32
			// srcs: (93, 30)(750) 816 --> (750) 816:PUGB0, pass, NI0
			9'd34 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 0 -> 33
			// srcs: (94, 31)(780) 855 --> (780) 855:PUGB0, pass, PENB
			9'd35 : rdata = 43'b1100011100001000000000000000000000100000000;
			// PEs: 32 -> 33
			// srcs: (100, 32)(750) 816 --> (750) 816:NI0, pass, PENB
			9'd36 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 32
			// srcs: (101, 33)(810) 1178 --> (810) 1178:PUGB0, pass, NI0
			9'd37 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 8 -> 33
			// srcs: (102, 34)(840) 64 --> (840) 64:PUGB1, pass, PENB
			9'd38 : rdata = 43'b1100011100011000000000000000000000100000000;
			// PEs: 32 -> 33
			// srcs: (108, 35)(810) 1178 --> (810) 1178:NI0, pass, PENB
			9'd39 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 8 -> 32
			// srcs: (109, 36)(870) 1024 --> (870) 1024:PUGB1, pass, NI0
			9'd40 : rdata = 43'b1100011100011000000001000000000000000000000;
			// PEs: 8 -> 33
			// srcs: (110, 37)(900) 2 --> (900) 2:PUGB1, pass, PENB
			9'd41 : rdata = 43'b1100011100011000000000000000000000100000000;
			// PEs: 32 -> 33
			// srcs: (116, 38)(870) 1024 --> (870) 1024:NI0, pass, PENB
			9'd42 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 8 -> 32
			// srcs: (117, 39)(930) 1305 --> (930) 1305:PUGB1, pass, NI0
			9'd43 : rdata = 43'b1100011100011000000001000000000000000000000;
			// PEs: 8 -> 33
			// srcs: (118, 40)(960) -33 --> (960) -33:PUGB1, pass, PENB
			9'd44 : rdata = 43'b1100011100011000000000000000000000100000000;
			// PEs: 32 -> 33
			// srcs: (124, 41)(930) 1305 --> (930) 1305:NI0, pass, PENB
			9'd45 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 8 -> 32
			// srcs: (125, 42)(990) 82 --> (990) 82:PUGB1, pass, NI0
			9'd46 : rdata = 43'b1100011100011000000001000000000000000000000;
			// PEs: 8 -> 33
			// srcs: (126, 43)(1020) -22 --> (1020) -22:PUGB1, pass, PENB
			9'd47 : rdata = 43'b1100011100011000000000000000000000100000000;
			// PEs: 32 -> 33
			// srcs: (132, 44)(990) 82 --> (990) 82:NI0, pass, PENB
			9'd48 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 32
			// srcs: (133, 45)(633) 672 --> (633) 672:PUGB0, pass, NI0
			9'd49 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 0 -> 33
			// srcs: (134, 46)(663) 165 --> (663) 165:PUGB0, pass, PENB
			9'd50 : rdata = 43'b1100011100001000000000000000000000100000000;
			// PEs: 33 -> 8
			// srcs: (139, 103)(1344) 60 --> (1344) 60:PEGB1, pass, PUGB1
			9'd51 : rdata = 43'b1100011100010000000000000000000000000001001;
			// PEs: 32 -> 33
			// srcs: (140, 47)(633) 672 --> (633) 672:NI0, pass, PENB
			9'd52 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 32
			// srcs: (141, 48)(693) 864 --> (693) 864:PUGB0, pass, NI0
			9'd53 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 0 -> 33
			// srcs: (142, 49)(723) 184 --> (723) 184:PUGB0, pass, PENB
			9'd54 : rdata = 43'b1100011100001000000000000000000000100000000;
			// PEs: 32 -> 33
			// srcs: (148, 50)(693) 864 --> (693) 864:NI0, pass, PENB
			9'd55 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 32
			// srcs: (149, 51)(753) 816 --> (753) 816:PUGB0, pass, NI0
			9'd56 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 0 -> 33
			// srcs: (150, 52)(783) 836 --> (783) 836:PUGB0, pass, PENB
			9'd57 : rdata = 43'b1100011100001000000000000000000000100000000;
			// PEs: 33 -> 8
			// srcs: (151, 117)(1291) 1070 --> (1291) 1070:PEGB1, pass, PUGB1
			9'd58 : rdata = 43'b1100011100010000000000000000000000000001001;
			// PEs: 32 -> 33
			// srcs: (156, 53)(753) 816 --> (753) 816:NI0, pass, PENB
			9'd59 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 32
			// srcs: (157, 54)(813) 62 --> (813) 62:PUGB0, pass, NI0
			9'd60 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 8 -> 33
			// srcs: (158, 55)(843) 1344 --> (843) 1344:PUGB1, pass, PENB
			9'd61 : rdata = 43'b1100011100011000000000000000000000100000000;
			// PEs: 32 -> 33
			// srcs: (164, 56)(813) 62 --> (813) 62:NI0, pass, PENB
			9'd62 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 8 -> 32
			// srcs: (165, 57)(873) 352 --> (873) 352:PUGB1, pass, NI0
			9'd63 : rdata = 43'b1100011100011000000001000000000000000000000;
			// PEs: 8 -> 33
			// srcs: (166, 58)(903) -37 --> (903) -37:PUGB1, pass, PENB
			9'd64 : rdata = 43'b1100011100011000000000000000000000100000000;
			// PEs: 32 -> 33
			// srcs: (172, 59)(873) 352 --> (873) 352:NI0, pass, PENB
			9'd65 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 8 -> 32
			// srcs: (173, 60)(933) 406 --> (933) 406:PUGB1, pass, NI0
			9'd66 : rdata = 43'b1100011100011000000001000000000000000000000;
			// PEs: 8 -> 33
			// srcs: (174, 61)(963) 33 --> (963) 33:PUGB1, pass, PENB
			9'd67 : rdata = 43'b1100011100011000000000000000000000100000000;
			// PEs: 32 -> 33
			// srcs: (180, 62)(933) 406 --> (933) 406:NI0, pass, PENB
			9'd68 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 8 -> 32
			// srcs: (181, 63)(993) 74 --> (993) 74:PUGB1, pass, NI0
			9'd69 : rdata = 43'b1100011100011000000001000000000000000000000;
			// PEs: 8 -> 33
			// srcs: (182, 64)(1023) 616 --> (1023) 616:PUGB1, pass, PENB
			9'd70 : rdata = 43'b1100011100011000000000000000000000100000000;
			// PEs: 32 -> 33
			// srcs: (188, 65)(993) 74 --> (993) 74:NI0, pass, PENB
			9'd71 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 32
			// srcs: (189, 66)(638) 28 --> (638) 28:PUGB0, pass, NI0
			9'd72 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 0 -> 33
			// srcs: (190, 67)(668) 264 --> (668) 264:PUGB0, pass, PENB
			9'd73 : rdata = 43'b1100011100001000000000000000000000100000000;
			// PEs: 33 -> 40
			// srcs: (195, 104)(1401) 690 --> (1401) 690:PEGB1, pass, PUNB
			9'd74 : rdata = 43'b1100011100010000000000000000000001000000000;
			// PEs: 32 -> 33
			// srcs: (196, 68)(638) 28 --> (638) 28:NI0, pass, PENB
			9'd75 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 32
			// srcs: (197, 69)(698) 432 --> (698) 432:PUGB0, pass, NI0
			9'd76 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 0 -> 33
			// srcs: (198, 70)(728) 966 --> (728) 966:PUGB0, pass, PENB
			9'd77 : rdata = 43'b1100011100001000000000000000000000100000000;
			// PEs: 32 -> 33
			// srcs: (204, 71)(698) 432 --> (698) 432:NI0, pass, PENB
			9'd78 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 32
			// srcs: (205, 72)(758) 936 --> (758) 936:PUGB0, pass, NI0
			9'd79 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 0 -> 33
			// srcs: (206, 73)(788) 399 --> (788) 399:PUGB0, pass, PENB
			9'd80 : rdata = 43'b1100011100001000000000000000000000100000000;
			// PEs: 32 -> 33
			// srcs: (212, 74)(758) 936 --> (758) 936:NI0, pass, PENB
			9'd81 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 32
			// srcs: (213, 75)(818) 837 --> (818) 837:PUGB0, pass, NI0
			9'd82 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 8 -> 33
			// srcs: (214, 76)(848) 864 --> (848) 864:PUGB1, pass, PENB
			9'd83 : rdata = 43'b1100011100011000000000000000000000100000000;
			// PEs: 32 -> 33
			// srcs: (220, 77)(818) 837 --> (818) 837:NI0, pass, PENB
			9'd84 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 8 -> 32
			// srcs: (221, 78)(878) 608 --> (878) 608:PUGB1, pass, NI0
			9'd85 : rdata = 43'b1100011100011000000001000000000000000000000;
			// PEs: 8 -> 33
			// srcs: (222, 79)(908) -20 --> (908) -20:PUGB1, pass, PENB
			9'd86 : rdata = 43'b1100011100011000000000000000000000100000000;
			// PEs: 32 -> 33
			// srcs: (228, 80)(878) 608 --> (878) 608:NI0, pass, PENB
			9'd87 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 8 -> 32
			// srcs: (229, 81)(938) -87 --> (938) -87:PUGB1, pass, NI0
			9'd88 : rdata = 43'b1100011100011000000001000000000000000000000;
			// PEs: 8 -> 33
			// srcs: (230, 82)(968) 231 --> (968) 231:PUGB1, pass, PENB
			9'd89 : rdata = 43'b1100011100011000000000000000000000100000000;
			// PEs: 32 -> 33
			// srcs: (236, 83)(938) -87 --> (938) -87:NI0, pass, PENB
			9'd90 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 8 -> 32
			// srcs: (237, 84)(998) 0 --> (998) 0:PUGB1, pass, NI0
			9'd91 : rdata = 43'b1100011100011000000001000000000000000000000;
			// PEs: 8 -> 33
			// srcs: (238, 85)(1028) 990 --> (1028) 990:PUGB1, pass, PENB
			9'd92 : rdata = 43'b1100011100011000000000000000000000100000000;
			// PEs: 32 -> 33
			// srcs: (244, 86)(998) 0 --> (998) 0:NI0, pass, PENB
			9'd93 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 32
			// srcs: (245, 87)(819) 868 --> (819) 868:PUGB0, pass, NI0
			9'd94 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 8 -> 33
			// srcs: (246, 88)(849) 320 --> (849) 320:PUGB1, pass, PENB
			9'd95 : rdata = 43'b1100011100011000000000000000000000100000000;
			// PEs: 33 -> 40
			// srcs: (251, 111)(1496) 990 --> (1496) 990:PEGB1, pass, PUNB
			9'd96 : rdata = 43'b1100011100010000000000000000000001000000000;
			// PEs: 32 -> 33
			// srcs: (252, 89)(819) 868 --> (819) 868:NI0, pass, PENB
			9'd97 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 8 -> 32
			// srcs: (253, 90)(879) 128 --> (879) 128:PUGB1, pass, NI0
			9'd98 : rdata = 43'b1100011100011000000001000000000000000000000;
			// PEs: 8 -> 33
			// srcs: (254, 91)(909) -37 --> (909) -37:PUGB1, pass, PENB
			9'd99 : rdata = 43'b1100011100011000000000000000000000100000000;
			// PEs: 32 -> 33
			// srcs: (260, 92)(879) 128 --> (879) 128:NI0, pass, PENB
			9'd100 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 8 -> 32
			// srcs: (261, 93)(939) 783 --> (939) 783:PUGB1, pass, NI0
			9'd101 : rdata = 43'b1100011100011000000001000000000000000000000;
			// PEs: 8 -> 33
			// srcs: (262, 94)(969) 858 --> (969) 858:PUGB1, pass, PENB
			9'd102 : rdata = 43'b1100011100011000000000000000000000100000000;
			// PEs: 33 -> 40
			// srcs: (263, 130)(1236) 3412 --> (1236) 3412:PEGB1, pass, PUNB
			9'd103 : rdata = 43'b1100011100010000000000000000000001000000000;
			// PEs: 32 -> 33
			// srcs: (268, 95)(939) 783 --> (939) 783:NI0, pass, PENB
			9'd104 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 8 -> 32
			// srcs: (269, 96)(999) 44 --> (999) 44:PUGB1, pass, NI0
			9'd105 : rdata = 43'b1100011100011000000001000000000000000000000;
			// PEs: 8 -> 33
			// srcs: (270, 97)(1029) -22 --> (1029) -22:PUGB1, pass, PENB
			9'd106 : rdata = 43'b1100011100011000000000000000000000100000000;
			// PEs: 33 -> 40
			// srcs: (271, 131)(1350) 2298 --> (1350) 2298:PEGB1, pass, PUNB
			9'd107 : rdata = 43'b1100011100010000000000000000000001000000000;
			// PEs: 32 -> 33
			// srcs: (276, 98)(999) 44 --> (999) 44:NI0, pass, PENB
			9'd108 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 56 -> 32
			// srcs: (277, 105)(1439) 368 --> (1439) 368:PUGB7, pass, NI0
			9'd109 : rdata = 43'b1100011101111000000001000000000000000000000;
			// PEs: 33 -> 40
			// srcs: (279, 132)(1407) 754 --> (1407) 754:PEGB1, pass, PUNB
			9'd110 : rdata = 43'b1100011100010000000000000000000001000000000;
			// PEs: 33 -> 40
			// srcs: (287, 134)(1502) 732 --> (1502) 732:PEGB1, pass, PUNB
			9'd111 : rdata = 43'b1100011100010000000000000000000001000000000;
			// PEs: 33 -> 40
			// srcs: (295, 136)(1410) 4943 --> (1410) 4943:PEGB1, pass, PUNB
			9'd112 : rdata = 43'b1100011100010000000000000000000001000000000;
			// PEs: 16 -> 33
			// srcs: (327, 106)(1440) 1572 --> (1440) 1572:PUGB2, pass, PENB
			9'd113 : rdata = 43'b1100011100101000000000000000000000100000000;
			// PEs: 32 -> 33
			// srcs: (333, 107)(1439) 368 --> (1439) 368:NI0, pass, PENB
			9'd114 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 56 -> 32
			// srcs: (334, 108)(1452) 118 --> (1452) 118:PUGB7, pass, NI0
			9'd115 : rdata = 43'b1100011101111000000001000000000000000000000;
			// PEs: 24 -> 33
			// srcs: (335, 109)(1453) 2034 --> (1453) 2034:PUNB, pass, PENB
			9'd116 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 33 -> 48
			// srcs: (340, 133)(1446) 1940 --> (1446) 1940:PEGB1, pass, PUGB6
			9'd117 : rdata = 43'b1100011100010000000000000000000000000001110;
			// PEs: 32 -> 33
			// srcs: (341, 110)(1452) 118 --> (1452) 118:NI0, pass, PENB
			9'd118 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 24 -> 33
			// srcs: (403, 112)(1511) 1372 --> (1511) 1372:PUNB, pass, PENB
			9'd119 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 16 -> 33
			// srcs: (404, 113)(1516) 474 --> (1516) 474:PUGB2, pass, PENB
			9'd120 : rdata = 43'b1100011100101000000000000000000000100000000;
			// PEs: 0 -> 32
			// srcs: (405, 114)(1739) 863 --> (1739) 863:PUGB0, pass, NI0
			9'd121 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 8 -> 33
			// srcs: (406, 115)(1740) 2120 --> (1740) 2120:PUGB1, pass, PENB
			9'd122 : rdata = 43'b1100011100011000000000000000000000100000000;
			// PEs: 32 -> 33
			// srcs: (412, 116)(1739) 863 --> (1739) 863:NI0, pass, PENB
			9'd123 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 33 -> 48
			// srcs: (415, 171)(1525) 2228 --> (1525) 2228:PEGB1, pass, PUGB6
			9'd124 : rdata = 43'b1100011100010000000000000000000000000001110;
			// PEs: 24 -> 33
			// srcs: (544, 118)(1463) 1127 --> (1463) 1127:PUNB, pass, PENB
			9'd125 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 24 -> 33
			// srcs: (705, 119)(1519) 2123 --> (1519) 2123:PUNB, pass, PENB
			9'd126 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 0 -> 32
			// srcs: (706, 120)(1690) 3957 --> (1690) 3957:PUGB0, pass, NI0
			9'd127 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 8 -> 33
			// srcs: (707, 121)(1691) 4091 --> (1691) 4091:PUGB1, pass, PENB
			9'd128 : rdata = 43'b1100011100011000000000000000000000100000000;
			// PEs: 33 -> 16
			// srcs: (712, 139)(1524) 4683 --> (1524) 4683:PEGB1, pass, PUGB2
			9'd129 : rdata = 43'b1100011100010000000000000000000000000001010;
			// PEs: 32 -> 33
			// srcs: (713, 122)(1690) 3957 --> (1690) 3957:NI0, pass, PENB
			9'd130 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 32
			// srcs: (714, 123)(1709) 668 --> (1709) 668:PUGB0, pass, NI0
			9'd131 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 24 -> 33
			// srcs: (715, 124)(1710) 2361 --> (1710) 2361:PUNB, pass, PENB
			9'd132 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 33 -> 24
			// srcs: (720, 152)(1695) 8048 --> (1695) 8048:PEGB1, pass, PUGB3
			9'd133 : rdata = 43'b1100011100010000000000000000000000000001011;
			// PEs: 32 -> 33
			// srcs: (721, 125)(1709) 668 --> (1709) 668:NI0, pass, PENB
			9'd134 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 33
			// srcs: (722, 126)(1747) 1080 --> (1747) 1080:PUGB0, pass, PENB
			9'd135 : rdata = 43'b1100011100001000000000000000000000100000000;
			// PEs: 0 -> 32
			// srcs: (723, 127)(1785) 3847 --> (1785) 3847:PUGB0, pass, NI0
			9'd136 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 40 -> 33
			// srcs: (724, 128)(1786) 3047 --> (1786) 3047:PUGB5, pass, PENB
			9'd137 : rdata = 43'b1100011101011000000000000000000000100000000;
			// PEs: 33 -> 24
			// srcs: (728, 153)(1714) 3029 --> (1714) 3029:PEGB1, pass, PUGB3
			9'd138 : rdata = 43'b1100011100010000000000000000000000000001011;
			// PEs: 32 -> 33
			// srcs: (730, 129)(1785) 3847 --> (1785) 3847:NI0, pass, PENB
			9'd139 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 24 -> 33
			// srcs: (926, 135)(1352) 855 --> (1352) 855:PUNB, pass, PENB
			9'd140 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 24 -> 33
			// srcs: (927, 137)(1466) 2331 --> (1466) 2331:PUNB, pass, PENB
			9'd141 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 24 -> 33
			// srcs: (928, 138)(1504) 683 --> (1504) 683:PUNB, pass, PENB
			9'd142 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 24 -> 32
			// srcs: (929, 140)(1618) 1450 --> (1618) 1450:PUNB, pass, NI0
			9'd143 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 8 -> 33
			// srcs: (930, 141)(1619) 3843 --> (1619) 3843:PUGB1, pass, PENB
			9'd144 : rdata = 43'b1100011100011000000000000000000000100000000;
			// PEs: 33 -> 40
			// srcs: (933, 168)(1355) 5478 --> (1355) 5478:PEGB1, pass, PUNB
			9'd145 : rdata = 43'b1100011100010000000000000000000001000000000;
			// PEs: 33 -> 40
			// srcs: (934, 169)(1469) 5610 --> (1469) 5610:PEGB1, pass, PUNB
			9'd146 : rdata = 43'b1100011100010000000000000000000001000000000;
			// PEs: 33 -> 40
			// srcs: (935, 170)(1507) 5409 --> (1507) 5409:PEGB1, pass, PUNB
			9'd147 : rdata = 43'b1100011100010000000000000000000001000000000;
			// PEs: 32 -> 33
			// srcs: (936, 142)(1618) 1450 --> (1618) 1450:NI0, pass, PENB
			9'd148 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 24 -> 32
			// srcs: (937, 143)(1637) 189 --> (1637) 189:PUNB, pass, NI0
			9'd149 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 8 -> 33
			// srcs: (938, 144)(1638) 3081 --> (1638) 3081:PUGB1, pass, PENB
			9'd150 : rdata = 43'b1100011100011000000000000000000000100000000;
			// PEs: 33 -> 48
			// srcs: (943, 172)(1621) 5293 --> (1621) 5293:PEGB1, pass, PUGB6
			9'd151 : rdata = 43'b1100011100010000000000000000000000000001110;
			// PEs: 32 -> 33
			// srcs: (944, 145)(1637) 189 --> (1637) 189:NI0, pass, PENB
			9'd152 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 24 -> 32
			// srcs: (945, 146)(1656) 1475 --> (1656) 1475:PUNB, pass, NI0
			9'd153 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 8 -> 33
			// srcs: (946, 147)(1657) 4043 --> (1657) 4043:PUGB1, pass, PENB
			9'd154 : rdata = 43'b1100011100011000000000000000000000100000000;
			// PEs: 33 -> 56
			// srcs: (951, 173)(1640) 3270 --> (1640) 3270:PEGB1, pass, PUGB7
			9'd155 : rdata = 43'b1100011100010000000000000000000000000001111;
			// PEs: 32 -> 33
			// srcs: (952, 148)(1656) 1475 --> (1656) 1475:NI0, pass, PENB
			9'd156 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 24 -> 32
			// srcs: (953, 149)(1675) 1935 --> (1675) 1935:PUNB, pass, NI0
			9'd157 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 8 -> 33
			// srcs: (954, 150)(1676) 3447 --> (1676) 3447:PUGB1, pass, PENB
			9'd158 : rdata = 43'b1100011100011000000000000000000000100000000;
			// PEs: 33 -> 56
			// srcs: (959, 174)(1659) 5518 --> (1659) 5518:PEGB1, pass, PUGB7
			9'd159 : rdata = 43'b1100011100010000000000000000000000000001111;
			// PEs: 32 -> 33
			// srcs: (960, 151)(1675) 1935 --> (1675) 1935:NI0, pass, PENB
			9'd160 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 16 -> 33
			// srcs: (961, 154)(1751) 2005 --> (1751) 2005:PUGB2, pass, PENB
			9'd161 : rdata = 43'b1100011100101000000000000000000000100000000;
			// PEs: 16 -> 33
			// srcs: (962, 155)(1789) 2117 --> (1789) 2117:PUGB2, pass, PENB
			9'd162 : rdata = 43'b1100011100101000000000000000000000100000000;
			// PEs: 40 -> 32
			// srcs: (963, 156)(1240) 4722 --> (1240) 4722:PUGB5, pass, NI0
			9'd163 : rdata = 43'b1100011101011000000001000000000000000000000;
			// PEs: 0 -> 33
			// srcs: (964, 157)(1241) 7417 --> (1241) 7417:PUGB0, pass, PENB
			9'd164 : rdata = 43'b1100011100001000000000000000000000100000000;
			// PEs: 33 -> 56
			// srcs: (967, 175)(1678) 5382 --> (1678) 5382:PEGB1, pass, PUGB7
			9'd165 : rdata = 43'b1100011100010000000000000000000000000001111;
			// PEs: 33 -> 56
			// srcs: (968, 176)(1754) 6068 --> (1754) 6068:PEGB1, pass, PUGB7
			9'd166 : rdata = 43'b1100011100010000000000000000000000000001111;
			// PEs: 33 -> 0
			// srcs: (969, 177)(1792) 9011 --> (1792) 9011:PEGB1, pass, PUGB0
			9'd167 : rdata = 43'b1100011100010000000000000000000000000001000;
			// PEs: 32 -> 33
			// srcs: (970, 158)(1240) 4722 --> (1240) 4722:NI0, pass, PENB
			9'd168 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 56 -> 32
			// srcs: (971, 159)(1278) 2151 --> (1278) 2151:PUGB7, pass, NI0
			9'd169 : rdata = 43'b1100011101111000000001000000000000000000000;
			// PEs: 24 -> 33
			// srcs: (1077, 160)(1279) 6449 --> (1279) 6449:PUNB, pass, PENB
			9'd170 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 32 -> 33
			// srcs: (1083, 161)(1278) 2151 --> (1278) 2151:NI0, pass, PENB
			9'd171 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 40 -> 32
			// srcs: (1084, 162)(1297) 5224 --> (1297) 5224:PUGB5, pass, NI0
			9'd172 : rdata = 43'b1100011101011000000001000000000000000000000;
			// PEs: 8 -> 33
			// srcs: (1085, 163)(1298) 6944 --> (1298) 6944:PUGB1, pass, PENB
			9'd173 : rdata = 43'b1100011100011000000000000000000000100000000;
			// PEs: 32 -> 33
			// srcs: (1091, 164)(1297) 5224 --> (1297) 5224:NI0, pass, PENB
			9'd174 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 56 -> 32
			// srcs: (1092, 165)(1316) 2571 --> (1316) 2571:PUGB7, pass, NI0
			9'd175 : rdata = 43'b1100011101111000000001000000000000000000000;
			// PEs: 8 -> 33
			// srcs: (1093, 166)(1317) 7939 --> (1317) 7939:PUGB1, pass, PENB
			9'd176 : rdata = 43'b1100011100011000000000000000000000100000000;
			// PEs: 32 -> 33
			// srcs: (1099, 167)(1316) 2571 --> (1316) 2571:NI0, pass, PENB
			9'd177 : rdata = 43'b1100010100000000000000000000000000100000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 33) begin
	always @(*) begin
		case(address)
			// PEs: 32 -> 
			// srcs: (16, 0)(714) 2116 --> (714) 2116:PENB, pass, 
			9'd0 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 32, 33 -> 32
			// srcs: (22, 1)(684) 1032, (714) 2116 --> (1225) 3148:PENB, ALU, +, PEGB0
			9'd1 : rdata = 43'b0000111011110001111110000000000000010000000;
			// PEs: 32 -> 
			// srcs: (24, 2)(774) 722 --> (774) 722:PENB, pass, 
			9'd2 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 32, 33 -> 32
			// srcs: (30, 3)(744) 120, (774) 722 --> (1226) 842:PENB, ALU, +, PEGB0
			9'd3 : rdata = 43'b0000111011110001111110000000000000010000000;
			// PEs: 32 -> 
			// srcs: (32, 4)(894) -22 --> (894) -22:PENB, pass, 
			9'd4 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 32, 33 -> 33
			// srcs: (38, 5)(864) 1216, (894) -22 --> (1228) 1194:PENB, ALU, +, NI0
			9'd5 : rdata = 43'b0000111011110001111111000000000000000000000;
			// PEs: 32 -> 
			// srcs: (40, 6)(954) 1551 --> (954) 1551:PENB, pass, 
			9'd6 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 32, 33 -> 33
			// srcs: (46, 7)(924) 667, (954) 1551 --> (1229) 2218:PENB, ALU, +, NI1
			9'd7 : rdata = 43'b0000111011110001111111000010000000000000000;
			// PEs: 32 -> 33
			// srcs: (48, 8)(1014) 462 --> (1014) 462:PENB, pass, NI2
			9'd8 : rdata = 43'b1100011011110000000001000100000000000000000;
			// PEs: 33 -> 33
			// srcs: (49, 126)(1228) 1194 --> (1228) 1194:NI0, pass, NI0
			9'd9 : rdata = 43'b1100010100000000000001000000000000000000000;
			// PEs: 33, 33 -> 33
			// srcs: (49, 66)(1228) 1194, (1229) 2218 --> (1236) 3412:ALU, NI1, +, NI3
			9'd10 : rdata = 43'b0000100111111101000011000110000000000000000;
			// PEs: 32, 33 -> 32
			// srcs: (54, 9)(984) 92, (1014) 462 --> (1230) 554:PENB, NI2, +, PEGB0
			9'd11 : rdata = 43'b0000111011110101000100000000000000010000000;
			// PEs: 32 -> 
			// srcs: (56, 10)(657) 66 --> (657) 66:PENB, pass, 
			9'd12 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 32, 33 -> 33
			// srcs: (62, 11)(627) 238, (657) 66 --> (1281) 304:PENB, ALU, +, NI0
			9'd13 : rdata = 43'b0000111011110001111111000000000000000000000;
			// PEs: 32 -> 
			// srcs: (64, 12)(717) 598 --> (717) 598:PENB, pass, 
			9'd14 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 32, 33 -> 33
			// srcs: (70, 13)(687) 168, (717) 598 --> (1282) 766:PENB, ALU, +, NI1
			9'd15 : rdata = 43'b0000111011110001111111000010000000000000000;
			// PEs: 32 -> 33
			// srcs: (72, 14)(777) 703 --> (777) 703:PENB, pass, NI2
			9'd16 : rdata = 43'b1100011011110000000001000100000000000000000;
			// PEs: 33 -> 33
			// srcs: (73, 127)(1281) 304 --> (1281) 304:NI0, pass, NI0
			9'd17 : rdata = 43'b1100010100000000000001000000000000000000000;
			// PEs: 33, 33 -> 33
			// srcs: (73, 67)(1281) 304, (1282) 766 --> (1291) 1070:ALU, NI1, +, NI4
			9'd18 : rdata = 43'b0000100111111101000011001000000000000000000;
			// PEs: 32, 33 -> 32
			// srcs: (78, 15)(747) 864, (777) 703 --> (1283) 1567:PENB, NI2, +, PEGB0
			9'd19 : rdata = 43'b0000111011110101000100000000000000010000000;
			// PEs: 32 -> 
			// srcs: (80, 16)(660) -22 --> (660) -22:PENB, pass, 
			9'd20 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 32, 33 -> 33
			// srcs: (86, 17)(630) 252, (660) -22 --> (1338) 230:PENB, ALU, +, NI0
			9'd21 : rdata = 43'b0000111011110001111111000000000000000000000;
			// PEs: 32 -> 
			// srcs: (88, 18)(720) 1288 --> (720) 1288:PENB, pass, 
			9'd22 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 32, 33 -> 33
			// srcs: (94, 19)(690) 192, (720) 1288 --> (1339) 1480:PENB, ALU, +, NI1
			9'd23 : rdata = 43'b0000111011110001111111000010000000000000000;
			// PEs: 32 -> 33
			// srcs: (96, 20)(780) 855 --> (780) 855:PENB, pass, NI2
			9'd24 : rdata = 43'b1100011011110000000001000100000000000000000;
			// PEs: 33 -> 33
			// srcs: (97, 128)(1338) 230 --> (1338) 230:NI0, pass, NI0
			9'd25 : rdata = 43'b1100010100000000000001000000000000000000000;
			// PEs: 33, 33 -> 33
			// srcs: (97, 68)(1338) 230, (1339) 1480 --> (1348) 1710:ALU, NI1, +, NI5
			9'd26 : rdata = 43'b0000100111111101000011001010000000000000000;
			// PEs: 32, 33 -> 33
			// srcs: (102, 21)(750) 816, (780) 855 --> (1340) 1671:PENB, NI2, +, NI0
			9'd27 : rdata = 43'b0000111011110101000101000000000000000000000;
			// PEs: 32 -> 
			// srcs: (104, 22)(840) 64 --> (840) 64:PENB, pass, 
			9'd28 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 32, 33 -> 33
			// srcs: (110, 23)(810) 1178, (840) 64 --> (1341) 1242:PENB, ALU, +, NI1
			9'd29 : rdata = 43'b0000111011110001111111000010000000000000000;
			// PEs: 32 -> 33
			// srcs: (112, 24)(900) 2 --> (900) 2:PENB, pass, NI2
			9'd30 : rdata = 43'b1100011011110000000001000100000000000000000;
			// PEs: 33 -> 33
			// srcs: (113, 129)(1340) 1671 --> (1340) 1671:NI0, pass, NI0
			9'd31 : rdata = 43'b1100010100000000000001000000000000000000000;
			// PEs: 33, 33 -> 
			// srcs: (113, 69)(1340) 1671, (1341) 1242 --> (1349) 2913:ALU, NI1, +, 
			9'd32 : rdata = 43'b0000100111111101000010000000000000000000000;
			// PEs: 33, 33 -> 33
			// srcs: (116, 87)(1348) 1710, (1349) 2913 --> (1353) 4623:NI5, ALU, +, NI0
			9'd33 : rdata = 43'b0000110100101001111111000000000000000000000;
			// PEs: 32, 33 -> 33
			// srcs: (118, 25)(870) 1024, (900) 2 --> (1342) 1026:PENB, NI2, +, NI1
			9'd34 : rdata = 43'b0000111011110101000101000010000000000000000;
			// PEs: 32 -> 
			// srcs: (120, 26)(960) -33 --> (960) -33:PENB, pass, 
			9'd35 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 32, 33 -> 33
			// srcs: (126, 27)(930) 1305, (960) -33 --> (1343) 1272:PENB, ALU, +, NI2
			9'd36 : rdata = 43'b0000111011110001111111000100000000000000000;
			// PEs: 32 -> 33
			// srcs: (128, 28)(1020) -22 --> (1020) -22:PENB, pass, NI5
			9'd37 : rdata = 43'b1100011011110000000001001010000000000000000;
			// PEs: 33 -> 33
			// srcs: (129, 130)(1342) 1026 --> (1342) 1026:NI1, pass, NI1
			9'd38 : rdata = 43'b1100010100001000000001000010000000000000000;
			// PEs: 33, 33 -> 33
			// srcs: (129, 70)(1342) 1026, (1343) 1272 --> (1350) 2298:ALU, NI2, +, NI6
			9'd39 : rdata = 43'b0000100111111101000101001100000000000000000;
			// PEs: 32, 33 -> 32
			// srcs: (134, 29)(990) 82, (1020) -22 --> (1344) 60:PENB, NI5, +, PEGB0
			9'd40 : rdata = 43'b0000111011110101001010000000000000010000000;
			// PEs: 32 -> 
			// srcs: (136, 30)(663) 165 --> (663) 165:PENB, pass, 
			9'd41 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 32, 33 -> 33
			// srcs: (142, 31)(633) 672, (663) 165 --> (1395) 837:PENB, ALU, +, NI1
			9'd42 : rdata = 43'b0000111011110001111111000010000000000000000;
			// PEs: 32 -> 33
			// srcs: (144, 32)(723) 184 --> (723) 184:PENB, pass, NI2
			9'd43 : rdata = 43'b1100011011110000000001000100000000000000000;
			// PEs: 33 -> 32
			// srcs: (145, 86)(1291) 1070 --> (1291) 1070:NI4, pass, PEGB0
			9'd44 : rdata = 43'b1100010100100000000000000000000000010000000;
			// PEs: 32, 33 -> 33
			// srcs: (150, 33)(693) 864, (723) 184 --> (1396) 1048:PENB, NI2, +, NI4
			9'd45 : rdata = 43'b0000111011110101000101001000000000000000000;
			// PEs: 32 -> 33
			// srcs: (152, 34)(783) 836 --> (783) 836:PENB, pass, NI2
			9'd46 : rdata = 43'b1100011011110000000001000100000000000000000;
			// PEs: 33 -> 33
			// srcs: (153, 131)(1395) 837 --> (1395) 837:NI1, pass, NI1
			9'd47 : rdata = 43'b1100010100001000000001000010000000000000000;
			// PEs: 33, 33 -> 33
			// srcs: (153, 71)(1395) 837, (1396) 1048 --> (1405) 1885:ALU, NI4, +, NI5
			9'd48 : rdata = 43'b0000100111111101001001001010000000000000000;
			// PEs: 32, 33 -> 33
			// srcs: (158, 35)(753) 816, (783) 836 --> (1397) 1652:PENB, NI2, +, NI1
			9'd49 : rdata = 43'b0000111011110101000101000010000000000000000;
			// PEs: 32 -> 
			// srcs: (160, 36)(843) 1344 --> (843) 1344:PENB, pass, 
			9'd50 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 32, 33 -> 33
			// srcs: (166, 37)(813) 62, (843) 1344 --> (1398) 1406:PENB, ALU, +, NI2
			9'd51 : rdata = 43'b0000111011110001111111000100000000000000000;
			// PEs: 32 -> 33
			// srcs: (168, 38)(903) -37 --> (903) -37:PENB, pass, NI4
			9'd52 : rdata = 43'b1100011011110000000001001000000000000000000;
			// PEs: 33 -> 33
			// srcs: (169, 132)(1397) 1652 --> (1397) 1652:NI1, pass, NI1
			9'd53 : rdata = 43'b1100010100001000000001000010000000000000000;
			// PEs: 33, 33 -> 
			// srcs: (169, 72)(1397) 1652, (1398) 1406 --> (1406) 3058:ALU, NI2, +, 
			9'd54 : rdata = 43'b0000100111111101000100000000000000000000000;
			// PEs: 33, 33 -> 33
			// srcs: (172, 88)(1405) 1885, (1406) 3058 --> (1410) 4943:NI5, ALU, +, NI1
			9'd55 : rdata = 43'b0000110100101001111111000010000000000000000;
			// PEs: 32, 33 -> 33
			// srcs: (174, 39)(873) 352, (903) -37 --> (1399) 315:PENB, NI4, +, NI2
			9'd56 : rdata = 43'b0000111011110101001001000100000000000000000;
			// PEs: 32 -> 
			// srcs: (176, 40)(963) 33 --> (963) 33:PENB, pass, 
			9'd57 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 32, 33 -> 33
			// srcs: (182, 41)(933) 406, (963) 33 --> (1400) 439:PENB, ALU, +, NI4
			9'd58 : rdata = 43'b0000111011110001111111001000000000000000000;
			// PEs: 32 -> 33
			// srcs: (184, 42)(1023) 616 --> (1023) 616:PENB, pass, NI5
			9'd59 : rdata = 43'b1100011011110000000001001010000000000000000;
			// PEs: 33 -> 33
			// srcs: (185, 133)(1399) 315 --> (1399) 315:NI2, pass, NI2
			9'd60 : rdata = 43'b1100010100010000000001000100000000000000000;
			// PEs: 33, 33 -> 33
			// srcs: (185, 73)(1399) 315, (1400) 439 --> (1407) 754:ALU, NI4, +, NI7
			9'd61 : rdata = 43'b0000100111111101001001001110000000000000000;
			// PEs: 32, 33 -> 32
			// srcs: (190, 43)(993) 74, (1023) 616 --> (1401) 690:PENB, NI5, +, PEGB0
			9'd62 : rdata = 43'b0000111011110101001010000000000000010000000;
			// PEs: 32 -> 
			// srcs: (192, 44)(668) 264 --> (668) 264:PENB, pass, 
			9'd63 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 32, 33 -> 33
			// srcs: (198, 45)(638) 28, (668) 264 --> (1490) 292:PENB, ALU, +, NI2
			9'd64 : rdata = 43'b0000111011110001111111000100000000000000000;
			// PEs: 32 -> 
			// srcs: (200, 46)(728) 966 --> (728) 966:PENB, pass, 
			9'd65 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 32, 33 -> 33
			// srcs: (206, 47)(698) 432, (728) 966 --> (1491) 1398:PENB, ALU, +, NI4
			9'd66 : rdata = 43'b0000111011110001111111001000000000000000000;
			// PEs: 32 -> 33
			// srcs: (208, 48)(788) 399 --> (788) 399:PENB, pass, NI5
			9'd67 : rdata = 43'b1100011011110000000001001010000000000000000;
			// PEs: 33 -> 33
			// srcs: (209, 134)(1490) 292 --> (1490) 292:NI2, pass, NI2
			9'd68 : rdata = 43'b1100010100010000000001000100000000000000000;
			// PEs: 33, 33 -> 33
			// srcs: (209, 78)(1490) 292, (1491) 1398 --> (1500) 1690:ALU, NI4, +, NI8
			9'd69 : rdata = 43'b0000100111111101001001010000000000000000000;
			// PEs: 32, 33 -> 33
			// srcs: (214, 49)(758) 936, (788) 399 --> (1492) 1335:PENB, NI5, +, NI2
			9'd70 : rdata = 43'b0000111011110101001011000100000000000000000;
			// PEs: 32 -> 
			// srcs: (216, 50)(848) 864 --> (848) 864:PENB, pass, 
			9'd71 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 32, 33 -> 33
			// srcs: (222, 51)(818) 837, (848) 864 --> (1493) 1701:PENB, ALU, +, NI4
			9'd72 : rdata = 43'b0000111011110001111111001000000000000000000;
			// PEs: 32 -> 33
			// srcs: (224, 52)(908) -20 --> (908) -20:PENB, pass, NI5
			9'd73 : rdata = 43'b1100011011110000000001001010000000000000000;
			// PEs: 33 -> 33
			// srcs: (225, 135)(1492) 1335 --> (1492) 1335:NI2, pass, NI2
			9'd74 : rdata = 43'b1100010100010000000001000100000000000000000;
			// PEs: 33, 33 -> 
			// srcs: (225, 79)(1492) 1335, (1493) 1701 --> (1501) 3036:ALU, NI4, +, 
			9'd75 : rdata = 43'b0000100111111101001000000000000000000000000;
			// PEs: 33, 33 -> 33
			// srcs: (228, 90)(1500) 1690, (1501) 3036 --> (1505) 4726:NI8, ALU, +, NI2
			9'd76 : rdata = 43'b0000110101000001111111000100000000000000000;
			// PEs: 32, 33 -> 33
			// srcs: (230, 53)(878) 608, (908) -20 --> (1494) 588:PENB, NI5, +, NI4
			9'd77 : rdata = 43'b0000111011110101001011001000000000000000000;
			// PEs: 32 -> 
			// srcs: (232, 54)(968) 231 --> (968) 231:PENB, pass, 
			9'd78 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 32, 33 -> 33
			// srcs: (238, 55)(938) -87, (968) 231 --> (1495) 144:PENB, ALU, +, NI5
			9'd79 : rdata = 43'b0000111011110001111111001010000000000000000;
			// PEs: 32 -> 33
			// srcs: (240, 56)(1028) 990 --> (1028) 990:PENB, pass, NI8
			9'd80 : rdata = 43'b1100011011110000000001010000000000000000000;
			// PEs: 33 -> 33
			// srcs: (241, 136)(1494) 588 --> (1494) 588:NI4, pass, NI4
			9'd81 : rdata = 43'b1100010100100000000001001000000000000000000;
			// PEs: 33, 33 -> 33
			// srcs: (241, 80)(1494) 588, (1495) 144 --> (1502) 732:ALU, NI5, +, NI9
			9'd82 : rdata = 43'b0000100111111101001011010010000000000000000;
			// PEs: 32, 33 -> 32
			// srcs: (246, 57)(998) 0, (1028) 990 --> (1496) 990:PENB, NI8, +, PEGB0
			9'd83 : rdata = 43'b0000111011110101010000000000000000010000000;
			// PEs: 32 -> 
			// srcs: (248, 58)(849) 320 --> (849) 320:PENB, pass, 
			9'd84 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 32, 33 -> 33
			// srcs: (254, 59)(819) 868, (849) 320 --> (1512) 1188:PENB, ALU, +, NI4
			9'd85 : rdata = 43'b0000111011110001111111001000000000000000000;
			// PEs: 32 -> 33
			// srcs: (256, 60)(909) -37 --> (909) -37:PENB, pass, NI5
			9'd86 : rdata = 43'b1100011011110000000001001010000000000000000;
			// PEs: 33 -> 32
			// srcs: (257, 99)(1236) 3412 --> (1236) 3412:NI3, pass, PEGB0
			9'd87 : rdata = 43'b1100010100011000000000000000000000010000000;
			// PEs: 32, 33 -> 33
			// srcs: (262, 61)(879) 128, (909) -37 --> (1513) 91:PENB, NI5, +, NI3
			9'd88 : rdata = 43'b0000111011110101001011000110000000000000000;
			// PEs: 32 -> 33
			// srcs: (264, 62)(969) 858 --> (969) 858:PENB, pass, NI5
			9'd89 : rdata = 43'b1100011011110000000001001010000000000000000;
			// PEs: 33 -> 32
			// srcs: (266, 100)(1350) 2298 --> (1350) 2298:NI6, pass, PEGB0
			9'd90 : rdata = 43'b1100010100110000000000000000000000010000000;
			// PEs: 32, 33 -> 33
			// srcs: (270, 63)(939) 783, (969) 858 --> (1514) 1641:PENB, NI5, +, NI6
			9'd91 : rdata = 43'b0000111011110101001011001100000000000000000;
			// PEs: 32 -> 33
			// srcs: (272, 64)(1029) -22 --> (1029) -22:PENB, pass, NI5
			9'd92 : rdata = 43'b1100011011110000000001001010000000000000000;
			// PEs: 33 -> 33
			// srcs: (273, 137)(1513) 91 --> (1513) 91:NI3, pass, NI3
			9'd93 : rdata = 43'b1100010100011000000001000110000000000000000;
			// PEs: 33, 33 -> 33
			// srcs: (273, 82)(1513) 91, (1514) 1641 --> (1521) 1732:ALU, NI6, +, NI8
			9'd94 : rdata = 43'b0000100111111101001101010000000000000000000;
			// PEs: 33 -> 32
			// srcs: (274, 101)(1407) 754 --> (1407) 754:NI7, pass, PEGB0
			9'd95 : rdata = 43'b1100010100111000000000000000000000010000000;
			// PEs: 32, 33 -> 33
			// srcs: (278, 65)(999) 44, (1029) -22 --> (1515) 22:PENB, NI5, +, NI3
			9'd96 : rdata = 43'b0000111011110101001011000110000000000000000;
			// PEs: 33 -> 32
			// srcs: (282, 102)(1502) 732 --> (1502) 732:NI9, pass, PEGB0
			9'd97 : rdata = 43'b1100010101001000000000000000000000010000000;
			// PEs: 33 -> 32
			// srcs: (290, 105)(1410) 4943 --> (1410) 4943:NI1, pass, PEGB0
			9'd98 : rdata = 43'b1100010100001000000000000000000000010000000;
			// PEs: 32 -> 
			// srcs: (329, 74)(1440) 1572 --> (1440) 1572:PENB, pass, 
			9'd99 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 32, 33 -> 32
			// srcs: (335, 75)(1439) 368, (1440) 1572 --> (1446) 1940:PENB, ALU, +, PEGB0
			9'd100 : rdata = 43'b0000111011110001111110000000000000010000000;
			// PEs: 32 -> 
			// srcs: (337, 76)(1453) 2034 --> (1453) 2034:PENB, pass, 
			9'd101 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 32, 33 -> 33
			// srcs: (343, 77)(1452) 118, (1453) 2034 --> (1462) 2152:PENB, ALU, +, NI1
			9'd102 : rdata = 43'b0000111011110001111111000010000000000000000;
			// PEs: 32, 33 -> 33
			// srcs: (406, 81)(1511) 1372, (1512) 1188 --> (1520) 2560:PENB, NI4, +, NI5
			9'd103 : rdata = 43'b0000111011110101001001001010000000000000000;
			// PEs: 33, 32 -> 33
			// srcs: (407, 83)(1515) 22, (1516) 474 --> (1522) 496:NI3, PENB, +, NI4
			9'd104 : rdata = 43'b0000110100011110111101001000000000000000000;
			// PEs: 32 -> 33
			// srcs: (408, 84)(1740) 2120 --> (1740) 2120:PENB, pass, NI3
			9'd105 : rdata = 43'b1100011011110000000001000110000000000000000;
			// PEs: 33 -> 33
			// srcs: (410, 138)(1521) 1732 --> (1521) 1732:NI8, pass, NI8
			9'd106 : rdata = 43'b1100010101000000000001010000000000000000000;
			// PEs: 33, 33 -> 32
			// srcs: (410, 103)(1521) 1732, (1522) 496 --> (1525) 2228:ALU, NI4, +, PEGB0
			9'd107 : rdata = 43'b0000100111111101001000000000000000010000000;
			// PEs: 32, 33 -> 33
			// srcs: (414, 85)(1739) 863, (1740) 2120 --> (1748) 2983:PENB, NI3, +, NI4
			9'd108 : rdata = 43'b0000111011110101000111001000000000000000000;
			// PEs: 33, 32 -> 33
			// srcs: (547, 89)(1462) 2152, (1463) 1127 --> (1467) 3279:NI1, PENB, +, NI3
			9'd109 : rdata = 43'b0000110100001110111101000110000000000000000;
			// PEs: 32, 33 -> 32
			// srcs: (707, 91)(1519) 2123, (1520) 2560 --> (1524) 4683:PENB, NI5, +, PEGB0
			9'd110 : rdata = 43'b0000111011110101001010000000000000010000000;
			// PEs: 32 -> 
			// srcs: (709, 92)(1691) 4091 --> (1691) 4091:PENB, pass, 
			9'd111 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 32, 33 -> 32
			// srcs: (715, 93)(1690) 3957, (1691) 4091 --> (1695) 8048:PENB, ALU, +, PEGB0
			9'd112 : rdata = 43'b0000111011110001111110000000000000010000000;
			// PEs: 32 -> 
			// srcs: (717, 94)(1710) 2361 --> (1710) 2361:PENB, pass, 
			9'd113 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 32, 33 -> 32
			// srcs: (723, 95)(1709) 668, (1710) 2361 --> (1714) 3029:PENB, ALU, +, PEGB0
			9'd114 : rdata = 43'b0000111011110001111110000000000000010000000;
			// PEs: 32, 33 -> 33
			// srcs: (724, 96)(1747) 1080, (1748) 2983 --> (1752) 4063:PENB, NI4, +, NI1
			9'd115 : rdata = 43'b0000111011110101001001000010000000000000000;
			// PEs: 32 -> 
			// srcs: (726, 97)(1786) 3047 --> (1786) 3047:PENB, pass, 
			9'd116 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 32, 33 -> 33
			// srcs: (732, 98)(1785) 3847, (1786) 3047 --> (1790) 6894:PENB, ALU, +, NI4
			9'd117 : rdata = 43'b0000111011110001111111001000000000000000000;
			// PEs: 32, 33 -> 32
			// srcs: (928, 104)(1352) 855, (1353) 4623 --> (1355) 5478:PENB, NI0, +, PEGB0
			9'd118 : rdata = 43'b0000111011110101000000000000000000010000000;
			// PEs: 32, 33 -> 32
			// srcs: (929, 106)(1466) 2331, (1467) 3279 --> (1469) 5610:PENB, NI3, +, PEGB0
			9'd119 : rdata = 43'b0000111011110101000110000000000000010000000;
			// PEs: 32, 33 -> 32
			// srcs: (930, 107)(1504) 683, (1505) 4726 --> (1507) 5409:PENB, NI2, +, PEGB0
			9'd120 : rdata = 43'b0000111011110101000100000000000000010000000;
			// PEs: 32 -> 
			// srcs: (932, 108)(1619) 3843 --> (1619) 3843:PENB, pass, 
			9'd121 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 32, 33 -> 32
			// srcs: (938, 109)(1618) 1450, (1619) 3843 --> (1621) 5293:PENB, ALU, +, PEGB0
			9'd122 : rdata = 43'b0000111011110001111110000000000000010000000;
			// PEs: 32 -> 
			// srcs: (940, 110)(1638) 3081 --> (1638) 3081:PENB, pass, 
			9'd123 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 32, 33 -> 32
			// srcs: (946, 111)(1637) 189, (1638) 3081 --> (1640) 3270:PENB, ALU, +, PEGB0
			9'd124 : rdata = 43'b0000111011110001111110000000000000010000000;
			// PEs: 32 -> 
			// srcs: (948, 112)(1657) 4043 --> (1657) 4043:PENB, pass, 
			9'd125 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 32, 33 -> 32
			// srcs: (954, 113)(1656) 1475, (1657) 4043 --> (1659) 5518:PENB, ALU, +, PEGB0
			9'd126 : rdata = 43'b0000111011110001111110000000000000010000000;
			// PEs: 32 -> 
			// srcs: (956, 114)(1676) 3447 --> (1676) 3447:PENB, pass, 
			9'd127 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 32, 33 -> 32
			// srcs: (962, 115)(1675) 1935, (1676) 3447 --> (1678) 5382:PENB, ALU, +, PEGB0
			9'd128 : rdata = 43'b0000111011110001111110000000000000010000000;
			// PEs: 32, 33 -> 32
			// srcs: (963, 116)(1751) 2005, (1752) 4063 --> (1754) 6068:PENB, NI1, +, PEGB0
			9'd129 : rdata = 43'b0000111011110101000010000000000000010000000;
			// PEs: 32, 33 -> 32
			// srcs: (964, 117)(1789) 2117, (1790) 6894 --> (1792) 9011:PENB, NI4, +, PEGB0
			9'd130 : rdata = 43'b0000111011110101001000000000000000010000000;
			// PEs: 32 -> 
			// srcs: (966, 118)(1241) 7417 --> (1241) 7417:PENB, pass, 
			9'd131 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 32, 33 -> 33
			// srcs: (972, 119)(1240) 4722, (1241) 7417 --> (1242) 12139:PENB, ALU, +, NW0
			9'd132 : rdata = 43'b0000111011110001111110000001000000000000000;
			// PEs: 32 -> 
			// srcs: (1079, 120)(1279) 6449 --> (1279) 6449:PENB, pass, 
			9'd133 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 32, 33 -> 33
			// srcs: (1085, 121)(1278) 2151, (1279) 6449 --> (1280) 8600:PENB, ALU, +, NW1
			9'd134 : rdata = 43'b0000111011110001111110000001000010000000000;
			// PEs: 32 -> 
			// srcs: (1087, 122)(1298) 6944 --> (1298) 6944:PENB, pass, 
			9'd135 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 32, 33 -> 33
			// srcs: (1093, 123)(1297) 5224, (1298) 6944 --> (1299) 12168:PENB, ALU, +, NW2
			9'd136 : rdata = 43'b0000111011110001111110000001000100000000000;
			// PEs: 32 -> 
			// srcs: (1095, 124)(1317) 7939 --> (1317) 7939:PENB, pass, 
			9'd137 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 32, 33 -> 33
			// srcs: (1101, 125)(1316) 2571, (1317) 7939 --> (1318) 10510:PENB, ALU, +, NW3
			9'd138 : rdata = 43'b0000111011110001111110000001000110000000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 34) begin
	always @(*) begin
		case(address)
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 35) begin
	always @(*) begin
		case(address)
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 36) begin
	always @(*) begin
		case(address)
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 37) begin
	always @(*) begin
		case(address)
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 38) begin
	always @(*) begin
		case(address)
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 39) begin
	always @(*) begin
		case(address)
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 40) begin
	always @(*) begin
		case(address)
			// PEs: 8 -> 40
			// srcs: (28, 0)(926) 116 --> (926) 116:PUGB1, pass, NI0
			9'd0 : rdata = 43'b1100011100011000000001000000000000000000000;
			// PEs: 8 -> 41
			// srcs: (29, 1)(956) 165 --> (956) 165:PUGB1, pass, PENB
			9'd1 : rdata = 43'b1100011100011000000000000000000000100000000;
			// PEs: 40 -> 41
			// srcs: (35, 2)(926) 116 --> (926) 116:NI0, pass, PENB
			9'd2 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 8 -> 40
			// srcs: (36, 3)(986) 56 --> (986) 56:PUGB1, pass, NI0
			9'd3 : rdata = 43'b1100011100011000000001000000000000000000000;
			// PEs: 8 -> 41
			// srcs: (37, 4)(1016) -22 --> (1016) -22:PUGB1, pass, PENB
			9'd4 : rdata = 43'b1100011100011000000000000000000000100000000;
			// PEs: 41 -> 56
			// srcs: (42, 87)(1267) 281 --> (1267) 281:PEGB1, pass, PUGB7
			9'd5 : rdata = 43'b1100011100010000000000000000000000000001111;
			// PEs: 40 -> 41
			// srcs: (43, 5)(986) 56 --> (986) 56:NI0, pass, PENB
			9'd6 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 40
			// srcs: (44, 6)(807) 310 --> (807) 310:PUGB0, pass, NI0
			9'd7 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 8 -> 41
			// srcs: (45, 7)(837) 1440 --> (837) 1440:PUGB1, pass, PENB
			9'd8 : rdata = 43'b1100011100011000000000000000000000100000000;
			// PEs: 41 -> 56
			// srcs: (50, 88)(1268) 34 --> (1268) 34:PEGB1, pass, PUGB7
			9'd9 : rdata = 43'b1100011100010000000000000000000000000001111;
			// PEs: 40 -> 41
			// srcs: (51, 8)(807) 310 --> (807) 310:NI0, pass, PENB
			9'd10 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 8 -> 40
			// srcs: (52, 9)(867) 896 --> (867) 896:PUGB1, pass, NI0
			9'd11 : rdata = 43'b1100011100011000000001000000000000000000000;
			// PEs: 8 -> 41
			// srcs: (53, 10)(897) -9 --> (897) -9:PUGB1, pass, PENB
			9'd12 : rdata = 43'b1100011100011000000000000000000000100000000;
			// PEs: 40 -> 41
			// srcs: (59, 11)(867) 896 --> (867) 896:NI0, pass, PENB
			9'd13 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 8 -> 40
			// srcs: (60, 12)(927) 29 --> (927) 29:PUGB1, pass, NI0
			9'd14 : rdata = 43'b1100011100011000000001000000000000000000000;
			// PEs: 8 -> 41
			// srcs: (61, 13)(957) 1320 --> (957) 1320:PUGB1, pass, PENB
			9'd15 : rdata = 43'b1100011100011000000000000000000000100000000;
			// PEs: 40 -> 41
			// srcs: (67, 14)(927) 29 --> (927) 29:NI0, pass, PENB
			9'd16 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 8 -> 40
			// srcs: (68, 15)(987) 94 --> (987) 94:PUGB1, pass, NI0
			9'd17 : rdata = 43'b1100011100011000000001000000000000000000000;
			// PEs: 8 -> 41
			// srcs: (69, 16)(1017) 968 --> (1017) 968:PUGB1, pass, PENB
			9'd18 : rdata = 43'b1100011100011000000000000000000000100000000;
			// PEs: 40 -> 41
			// srcs: (75, 17)(987) 94 --> (987) 94:NI0, pass, PENB
			9'd19 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 16 -> 40
			// srcs: (76, 18)(1047) 1044 --> (1047) 1044:PUGB2, pass, NI0
			9'd20 : rdata = 43'b1100011100101000000001000000000000000000000;
			// PEs: 16 -> 41
			// srcs: (77, 19)(1077) 882 --> (1077) 882:PUGB2, pass, PENB
			9'd21 : rdata = 43'b1100011100101000000000000000000000100000000;
			// PEs: 40 -> 41
			// srcs: (83, 20)(1047) 1044 --> (1047) 1044:NI0, pass, PENB
			9'd22 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 16 -> 40
			// srcs: (84, 21)(1107) 805 --> (1107) 805:PUGB2, pass, NI0
			9'd23 : rdata = 43'b1100011100101000000001000000000000000000000;
			// PEs: 16 -> 41
			// srcs: (85, 22)(1137) 598 --> (1137) 598:PUGB2, pass, PENB
			9'd24 : rdata = 43'b1100011100101000000000000000000000100000000;
			// PEs: 40 -> 41
			// srcs: (91, 23)(1107) 805 --> (1107) 805:NI0, pass, PENB
			9'd25 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 16 -> 40
			// srcs: (92, 24)(1167) 162 --> (1167) 162:PUGB2, pass, NI0
			9'd26 : rdata = 43'b1100011100101000000001000000000000000000000;
			// PEs: 16 -> 41
			// srcs: (93, 25)(1197) 992 --> (1197) 992:PUGB2, pass, PENB
			9'd27 : rdata = 43'b1100011100101000000000000000000000100000000;
			// PEs: 40 -> 41
			// srcs: (99, 26)(1167) 162 --> (1167) 162:NI0, pass, PENB
			9'd28 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 40
			// srcs: (100, 27)(628) 336 --> (628) 336:PUGB0, pass, NI0
			9'd29 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 0 -> 41
			// srcs: (101, 28)(658) 308 --> (658) 308:PUGB0, pass, PENB
			9'd30 : rdata = 43'b1100011100001000000000000000000000100000000;
			// PEs: 40 -> 41
			// srcs: (107, 29)(628) 336 --> (628) 336:NI0, pass, PENB
			9'd31 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 40
			// srcs: (108, 30)(632) 112 --> (632) 112:PUGB0, pass, NI0
			9'd32 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 0 -> 41
			// srcs: (109, 31)(662) 264 --> (662) 264:PUGB0, pass, PENB
			9'd33 : rdata = 43'b1100011100001000000000000000000000100000000;
			// PEs: 41 -> 48
			// srcs: (114, 90)(1300) 644 --> (1300) 644:PEGB1, pass, PUNB
			9'd34 : rdata = 43'b1100011100010000000000000000000001000000000;
			// PEs: 40 -> 41
			// srcs: (115, 32)(632) 112 --> (632) 112:NI0, pass, PENB
			9'd35 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 40
			// srcs: (116, 33)(692) 456 --> (692) 456:PUGB0, pass, NI0
			9'd36 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 0 -> 41
			// srcs: (117, 34)(722) 1564 --> (722) 1564:PUGB0, pass, PENB
			9'd37 : rdata = 43'b1100011100001000000000000000000000100000000;
			// PEs: 40 -> 41
			// srcs: (123, 35)(692) 456 --> (692) 456:NI0, pass, PENB
			9'd38 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 40
			// srcs: (124, 36)(752) 312 --> (752) 312:PUGB0, pass, NI0
			9'd39 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 0 -> 41
			// srcs: (125, 37)(782) 589 --> (782) 589:PUGB0, pass, PENB
			9'd40 : rdata = 43'b1100011100001000000000000000000000100000000;
			// PEs: 40 -> 41
			// srcs: (131, 38)(752) 312 --> (752) 312:NI0, pass, PENB
			9'd41 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 16 -> 40
			// srcs: (132, 39)(1113) 299 --> (1113) 299:PUGB2, pass, NI0
			9'd42 : rdata = 43'b1100011100101000000001000000000000000000000;
			// PEs: 16 -> 41
			// srcs: (133, 40)(1143) 390 --> (1143) 390:PUGB2, pass, PENB
			9'd43 : rdata = 43'b1100011100101000000000000000000000100000000;
			// PEs: 41 -> 48
			// srcs: (138, 91)(1378) 901 --> (1378) 901:PEGB1, pass, PUNB
			9'd44 : rdata = 43'b1100011100010000000000000000000001000000000;
			// PEs: 40 -> 41
			// srcs: (139, 41)(1113) 299 --> (1113) 299:NI0, pass, PENB
			9'd45 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 16 -> 40
			// srcs: (140, 42)(1173) 36 --> (1173) 36:PUGB2, pass, NI0
			9'd46 : rdata = 43'b1100011100101000000001000000000000000000000;
			// PEs: 16 -> 41
			// srcs: (141, 43)(1203) 527 --> (1203) 527:PUGB2, pass, PENB
			9'd47 : rdata = 43'b1100011100101000000000000000000000100000000;
			// PEs: 40 -> 41
			// srcs: (147, 44)(1173) 36 --> (1173) 36:NI0, pass, PENB
			9'd48 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 40
			// srcs: (148, 45)(634) 448 --> (634) 448:PUGB0, pass, NI0
			9'd49 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 0 -> 41
			// srcs: (149, 46)(664) 528 --> (664) 528:PUGB0, pass, PENB
			9'd50 : rdata = 43'b1100011100001000000000000000000000100000000;
			// PEs: 40 -> 41
			// srcs: (155, 47)(634) 448 --> (634) 448:NI0, pass, PENB
			9'd51 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 40
			// srcs: (156, 48)(694) 960 --> (694) 960:PUGB0, pass, NI0
			9'd52 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 0 -> 41
			// srcs: (157, 49)(724) 874 --> (724) 874:PUGB0, pass, PENB
			9'd53 : rdata = 43'b1100011100001000000000000000000000100000000;
			// PEs: 40 -> 41
			// srcs: (163, 50)(694) 960 --> (694) 960:NI0, pass, PENB
			9'd54 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 40
			// srcs: (164, 51)(754) 1176 --> (754) 1176:PUGB0, pass, NI0
			9'd55 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 0 -> 41
			// srcs: (165, 52)(784) -38 --> (784) -38:PUGB0, pass, PENB
			9'd56 : rdata = 43'b1100011100001000000000000000000000100000000;
			// PEs: 40 -> 41
			// srcs: (171, 53)(754) 1176 --> (754) 1176:NI0, pass, PENB
			9'd57 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 40
			// srcs: (172, 54)(814) 744 --> (814) 744:PUGB0, pass, NI0
			9'd58 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 8 -> 41
			// srcs: (173, 55)(844) 160 --> (844) 160:PUGB1, pass, PENB
			9'd59 : rdata = 43'b1100011100011000000000000000000000100000000;
			// PEs: 40 -> 41
			// srcs: (179, 56)(814) 744 --> (814) 744:NI0, pass, PENB
			9'd60 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 8 -> 40
			// srcs: (180, 57)(874) 1568 --> (874) 1568:PUGB1, pass, NI0
			9'd61 : rdata = 43'b1100011100011000000001000000000000000000000;
			// PEs: 8 -> 41
			// srcs: (181, 58)(904) -4 --> (904) -4:PUGB1, pass, PENB
			9'd62 : rdata = 43'b1100011100011000000000000000000000100000000;
			// PEs: 40 -> 41
			// srcs: (187, 59)(874) 1568 --> (874) 1568:NI0, pass, PENB
			9'd63 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 40
			// srcs: (188, 60)(640) -28 --> (640) -28:PUGB0, pass, NI0
			9'd64 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 0 -> 41
			// srcs: (189, 61)(670) 44 --> (670) 44:PUGB0, pass, PENB
			9'd65 : rdata = 43'b1100011100001000000000000000000000100000000;
			// PEs: 41 -> 48
			// srcs: (194, 95)(1418) 1564 --> (1418) 1564:PEGB1, pass, PUNB
			9'd66 : rdata = 43'b1100011100010000000000000000000001000000000;
			// PEs: 40 -> 41
			// srcs: (195, 62)(640) -28 --> (640) -28:NI0, pass, PENB
			9'd67 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 40
			// srcs: (196, 63)(700) 624 --> (700) 624:PUGB0, pass, NI0
			9'd68 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 0 -> 41
			// srcs: (197, 64)(730) 828 --> (730) 828:PUGB0, pass, PENB
			9'd69 : rdata = 43'b1100011100001000000000000000000000100000000;
			// PEs: 40 -> 41
			// srcs: (203, 65)(700) 624 --> (700) 624:NI0, pass, PENB
			9'd70 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 40
			// srcs: (204, 66)(760) 600 --> (760) 600:PUGB0, pass, NI0
			9'd71 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 0 -> 41
			// srcs: (205, 67)(790) 779 --> (790) 779:PUGB0, pass, PENB
			9'd72 : rdata = 43'b1100011100001000000000000000000000100000000;
			// PEs: 40 -> 41
			// srcs: (211, 68)(760) 600 --> (760) 600:NI0, pass, PENB
			9'd73 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 40
			// srcs: (212, 69)(820) 837 --> (820) 837:PUGB0, pass, NI0
			9'd74 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 8 -> 41
			// srcs: (213, 70)(850) 480 --> (850) 480:PUGB1, pass, PENB
			9'd75 : rdata = 43'b1100011100011000000000000000000000100000000;
			// PEs: 40 -> 41
			// srcs: (219, 71)(820) 837 --> (820) 837:NI0, pass, PENB
			9'd76 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 8 -> 40
			// srcs: (220, 72)(880) 704 --> (880) 704:PUGB1, pass, NI0
			9'd77 : rdata = 43'b1100011100011000000001000000000000000000000;
			// PEs: 8 -> 41
			// srcs: (221, 73)(910) -2 --> (910) -2:PUGB1, pass, PENB
			9'd78 : rdata = 43'b1100011100011000000000000000000000100000000;
			// PEs: 40 -> 41
			// srcs: (227, 74)(880) 704 --> (880) 704:NI0, pass, PENB
			9'd79 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 8 -> 40
			// srcs: (228, 75)(940) 348 --> (940) 348:PUGB1, pass, NI0
			9'd80 : rdata = 43'b1100011100011000000001000000000000000000000;
			// PEs: 8 -> 41
			// srcs: (229, 76)(970) 891 --> (970) 891:PUGB1, pass, PENB
			9'd81 : rdata = 43'b1100011100011000000000000000000000100000000;
			// PEs: 41 -> 16
			// srcs: (232, 117)(1543) 4164 --> (1543) 4164:PEGB1, pass, PUGB2
			9'd82 : rdata = 43'b1100011100010000000000000000000000000001010;
			// PEs: 40 -> 41
			// srcs: (235, 77)(940) 348 --> (940) 348:NI0, pass, PENB
			9'd83 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 8 -> 40
			// srcs: (236, 78)(1000) 52 --> (1000) 52:PUGB1, pass, NI0
			9'd84 : rdata = 43'b1100011100011000000001000000000000000000000;
			// PEs: 8 -> 41
			// srcs: (237, 79)(1030) 462 --> (1030) 462:PUGB1, pass, PENB
			9'd85 : rdata = 43'b1100011100011000000000000000000000100000000;
			// PEs: 40 -> 41
			// srcs: (243, 80)(1000) 52 --> (1000) 52:NI0, pass, PENB
			9'd86 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 32 -> 40
			// srcs: (244, 81)(1226) 842 --> (1226) 842:PUNB, pass, NI0
			9'd87 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 16 -> 41
			// srcs: (245, 82)(1227) 2387 --> (1227) 2387:PUGB2, pass, PENB
			9'd88 : rdata = 43'b1100011100101000000000000000000000100000000;
			// PEs: 41 -> 48
			// srcs: (250, 99)(1534) 514 --> (1534) 514:PEGB1, pass, PUNB
			9'd89 : rdata = 43'b1100011100010000000000000000000001000000000;
			// PEs: 40 -> 41
			// srcs: (251, 83)(1226) 842 --> (1226) 842:NI0, pass, PENB
			9'd90 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 32 -> 40
			// srcs: (252, 84)(1230) 554 --> (1230) 554:PUNB, pass, NI0
			9'd91 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 41 -> 48
			// srcs: (258, 103)(1235) 3229 --> (1235) 3229:PEGB1, pass, PUNB
			9'd92 : rdata = 43'b1100011100010000000000000000000001000000000;
			// PEs: 41 -> 48
			// srcs: (266, 105)(1386) 2396 --> (1386) 2396:PEGB1, pass, PUNB
			9'd93 : rdata = 43'b1100011100010000000000000000000001000000000;
			// PEs: 41 -> 48
			// srcs: (274, 113)(1540) 1941 --> (1540) 1941:PEGB1, pass, PUNB
			9'd94 : rdata = 43'b1100011100010000000000000000000001000000000;
			// PEs: 16 -> 41
			// srcs: (331, 85)(1231) 756 --> (1231) 756:PUGB2, pass, PENB
			9'd95 : rdata = 43'b1100011100101000000000000000000000100000000;
			// PEs: 40 -> 41
			// srcs: (337, 86)(1230) 554 --> (1230) 554:NI0, pass, PENB
			9'd96 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 32 -> 41
			// srcs: (338, 89)(1283) 1567 --> (1283) 1567:PUNB, pass, PENB
			9'd97 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 32 -> 40
			// srcs: (339, 92)(1401) 690 --> (1401) 690:PUNB, pass, NI0
			9'd98 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 16 -> 41
			// srcs: (340, 93)(1402) 1053 --> (1402) 1053:PUGB2, pass, PENB
			9'd99 : rdata = 43'b1100011100101000000000000000000000100000000;
			// PEs: 41 -> 8
			// srcs: (345, 104)(1292) 3317 --> (1292) 3317:PEGB1, pass, PUGB1
			9'd100 : rdata = 43'b1100011100010000000000000000000000000001001;
			// PEs: 40 -> 41
			// srcs: (346, 94)(1401) 690 --> (1401) 690:NI0, pass, PENB
			9'd101 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 32 -> 40
			// srcs: (347, 96)(1496) 990 --> (1496) 990:PUNB, pass, NI0
			9'd102 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 16 -> 41
			// srcs: (348, 97)(1497) 1764 --> (1497) 1764:PUGB2, pass, PENB
			9'd103 : rdata = 43'b1100011100101000000000000000000000100000000;
			// PEs: 40 -> 41
			// srcs: (354, 98)(1496) 990 --> (1496) 990:NI0, pass, PENB
			9'd104 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 40
			// srcs: (355, 100)(1777) 1462 --> (1777) 1462:PUGB0, pass, NI0
			9'd105 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 8 -> 41
			// srcs: (356, 101)(1778) 1585 --> (1778) 1585:PUGB1, pass, PENB
			9'd106 : rdata = 43'b1100011100011000000000000000000000100000000;
			// PEs: 41 -> 8
			// srcs: (357, 114)(1295) 2557 --> (1295) 2557:PEGB1, pass, PUGB1
			9'd107 : rdata = 43'b1100011100010000000000000000000000000001001;
			// PEs: 40 -> 41
			// srcs: (362, 102)(1777) 1462 --> (1777) 1462:NI0, pass, PENB
			9'd108 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 41 -> 8
			// srcs: (365, 116)(1429) 4852 --> (1429) 4852:PEGB1, pass, PUGB1
			9'd109 : rdata = 43'b1100011100010000000000000000000000000001001;
			// PEs: 41 -> 32
			// srcs: (369, 106)(1786) 3047 --> (1786) 3047:PEGB1, pass, PUGB4
			9'd110 : rdata = 43'b1100011100010000000000000000000000000001100;
			// PEs: 32 -> 41
			// srcs: (471, 107)(1236) 3412 --> (1236) 3412:PUNB, pass, PENB
			9'd111 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 32 -> 40
			// srcs: (472, 108)(1350) 2298 --> (1350) 2298:PUNB, pass, NI0
			9'd112 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 8 -> 41
			// srcs: (473, 109)(1351) 1875 --> (1351) 1875:PUGB1, pass, PENB
			9'd113 : rdata = 43'b1100011100011000000000000000000000100000000;
			// PEs: 32 -> 42
			// srcs: (474, 111)(1407) 754 --> (1407) 754:PUNB, pass, PEGB2
			9'd114 : rdata = 43'b1100011011111000000000000000000000010100000;
			// PEs: 41 -> 32
			// srcs: (478, 118)(1240) 4722 --> (1240) 4722:PEGB1, pass, PUGB4
			9'd115 : rdata = 43'b1100011100010000000000000000000000000001100;
			// PEs: 40 -> 41
			// srcs: (479, 110)(1350) 2298 --> (1350) 2298:NI0, pass, PENB
			9'd116 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 32 -> 41
			// srcs: (480, 112)(1502) 732 --> (1502) 732:PUNB, pass, PENB
			9'd117 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 32 -> 41
			// srcs: (481, 115)(1410) 4943 --> (1410) 4943:PUNB, pass, PENB
			9'd118 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 0 -> 40
			// srcs: (482, 120)(1335) 4432 --> (1335) 4432:PUGB0, pass, NI0
			9'd119 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 41 -> 32
			// srcs: (489, 119)(1297) 5224 --> (1297) 5224:PEGB1, pass, PUGB4
			9'd120 : rdata = 43'b1100011100010000000000000000000000000001100;
			// PEs: 16 -> 41
			// srcs: (1020, 121)(1336) 4389 --> (1336) 4389:PUGB2, pass, PENB
			9'd121 : rdata = 43'b1100011100101000000000000000000000100000000;
			// PEs: 40 -> 41
			// srcs: (1027, 122)(1335) 4432 --> (1335) 4432:NI0, pass, PENB
			9'd122 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 32 -> 41
			// srcs: (1028, 123)(1355) 5478 --> (1355) 5478:PUNB, pass, PENB
			9'd123 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 48 -> 40
			// srcs: (1029, 124)(1430) 5992 --> (1430) 5992:PUGB6, pass, NI0
			9'd124 : rdata = 43'b1100011101101000000001000000000000000000000;
			// PEs: 8 -> 41
			// srcs: (1030, 125)(1431) 6812 --> (1431) 6812:PUGB1, pass, PENB
			9'd125 : rdata = 43'b1100011100011000000000000000000000100000000;
			// PEs: 40 -> 41
			// srcs: (1036, 126)(1430) 5992 --> (1430) 5992:NI0, pass, PENB
			9'd126 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 16 -> 40
			// srcs: (1841, 127)(1468) 3219 --> (1468) 3219:PUGB2, pass, NI0
			9'd127 : rdata = 43'b1100011100101000000001000000000000000000000;
			// PEs: 32 -> 41
			// srcs: (1842, 128)(1469) 5610 --> (1469) 5610:PUNB, pass, PENB
			9'd128 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 40 -> 41
			// srcs: (1848, 129)(1468) 3219 --> (1468) 3219:NI0, pass, PENB
			9'd129 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 32 -> 41
			// srcs: (1849, 130)(1507) 5409 --> (1507) 5409:PUNB, pass, PENB
			9'd130 : rdata = 43'b1100011011111000000000000000000000100000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 41) begin
	always @(*) begin
		case(address)
			// PEs: 40 -> 
			// srcs: (31, 0)(956) 165 --> (956) 165:PENB, pass, 
			9'd0 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 40, 41 -> 40
			// srcs: (37, 1)(926) 116, (956) 165 --> (1267) 281:PENB, ALU, +, PEGB0
			9'd1 : rdata = 43'b0000111011110001111110000000000000010000000;
			// PEs: 40 -> 
			// srcs: (39, 2)(1016) -22 --> (1016) -22:PENB, pass, 
			9'd2 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 40, 41 -> 40
			// srcs: (45, 3)(986) 56, (1016) -22 --> (1268) 34:PENB, ALU, +, PEGB0
			9'd3 : rdata = 43'b0000111011110001111110000000000000010000000;
			// PEs: 40 -> 
			// srcs: (47, 4)(837) 1440 --> (837) 1440:PENB, pass, 
			9'd4 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 40, 41 -> 41
			// srcs: (53, 5)(807) 310, (837) 1440 --> (1284) 1750:PENB, ALU, +, NI0
			9'd5 : rdata = 43'b0000111011110001111111000000000000000000000;
			// PEs: 40 -> 
			// srcs: (55, 6)(897) -9 --> (897) -9:PENB, pass, 
			9'd6 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 40, 41 -> 41
			// srcs: (61, 7)(867) 896, (897) -9 --> (1285) 887:PENB, ALU, +, NI1
			9'd7 : rdata = 43'b0000111011110001111111000010000000000000000;
			// PEs: 40 -> 
			// srcs: (63, 8)(957) 1320 --> (957) 1320:PENB, pass, 
			9'd8 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 40, 41 -> 41
			// srcs: (69, 9)(927) 29, (957) 1320 --> (1286) 1349:PENB, ALU, +, NI2
			9'd9 : rdata = 43'b0000111011110001111111000100000000000000000;
			// PEs: 40 -> 41
			// srcs: (71, 10)(1017) 968 --> (1017) 968:PENB, pass, NI3
			9'd10 : rdata = 43'b1100011011110000000001000110000000000000000;
			// PEs: 41 -> 41
			// srcs: (72, 96)(1285) 887 --> (1285) 887:NI1, pass, NI1
			9'd11 : rdata = 43'b1100010100001000000001000010000000000000000;
			// PEs: 41, 41 -> 41
			// srcs: (72, 59)(1285) 887, (1286) 1349 --> (1293) 2236:ALU, NI2, +, NI4
			9'd12 : rdata = 43'b0000100111111101000101001000000000000000000;
			// PEs: 40, 41 -> 41
			// srcs: (77, 11)(987) 94, (1017) 968 --> (1287) 1062:PENB, NI3, +, NI1
			9'd13 : rdata = 43'b0000111011110101000111000010000000000000000;
			// PEs: 40 -> 
			// srcs: (79, 12)(1077) 882 --> (1077) 882:PENB, pass, 
			9'd14 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 40, 41 -> 41
			// srcs: (85, 13)(1047) 1044, (1077) 882 --> (1288) 1926:PENB, ALU, +, NI2
			9'd15 : rdata = 43'b0000111011110001111111000100000000000000000;
			// PEs: 40 -> 41
			// srcs: (87, 14)(1137) 598 --> (1137) 598:PENB, pass, NI3
			9'd16 : rdata = 43'b1100011011110000000001000110000000000000000;
			// PEs: 41 -> 41
			// srcs: (88, 97)(1287) 1062 --> (1287) 1062:NI1, pass, NI1
			9'd17 : rdata = 43'b1100010100001000000001000010000000000000000;
			// PEs: 41, 41 -> 
			// srcs: (88, 60)(1287) 1062, (1288) 1926 --> (1294) 2988:ALU, NI2, +, 
			9'd18 : rdata = 43'b0000100111111101000100000000000000000000000;
			// PEs: 41, 41 -> 41
			// srcs: (91, 79)(1293) 2236, (1294) 2988 --> (1297) 5224:NI4, ALU, +, NI1
			9'd19 : rdata = 43'b0000110100100001111111000010000000000000000;
			// PEs: 40, 41 -> 41
			// srcs: (93, 15)(1107) 805, (1137) 598 --> (1289) 1403:PENB, NI3, +, NI2
			9'd20 : rdata = 43'b0000111011110101000111000100000000000000000;
			// PEs: 40 -> 
			// srcs: (95, 16)(1197) 992 --> (1197) 992:PENB, pass, 
			9'd21 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 40, 41 -> 41
			// srcs: (101, 17)(1167) 162, (1197) 992 --> (1290) 1154:PENB, ALU, +, NI3
			9'd22 : rdata = 43'b0000111011110001111111000110000000000000000;
			// PEs: 40 -> 41
			// srcs: (103, 18)(658) 308 --> (658) 308:PENB, pass, NI4
			9'd23 : rdata = 43'b1100011011110000000001001000000000000000000;
			// PEs: 41 -> 41
			// srcs: (104, 98)(1289) 1403 --> (1289) 1403:NI2, pass, NI2
			9'd24 : rdata = 43'b1100010100010000000001000100000000000000000;
			// PEs: 41, 41 -> 41
			// srcs: (104, 73)(1289) 1403, (1290) 1154 --> (1295) 2557:ALU, NI3, +, NI5
			9'd25 : rdata = 43'b0000100111111101000111001010000000000000000;
			// PEs: 40, 41 -> 40
			// srcs: (109, 19)(628) 336, (658) 308 --> (1300) 644:PENB, NI4, +, PEGB0
			9'd26 : rdata = 43'b0000111011110101001000000000000000010000000;
			// PEs: 40 -> 
			// srcs: (111, 20)(662) 264 --> (662) 264:PENB, pass, 
			9'd27 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 40, 41 -> 41
			// srcs: (117, 21)(632) 112, (662) 264 --> (1376) 376:PENB, ALU, +, NI2
			9'd28 : rdata = 43'b0000111011110001111111000100000000000000000;
			// PEs: 40 -> 
			// srcs: (119, 22)(722) 1564 --> (722) 1564:PENB, pass, 
			9'd29 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 40, 41 -> 41
			// srcs: (125, 23)(692) 456, (722) 1564 --> (1377) 2020:PENB, ALU, +, NI3
			9'd30 : rdata = 43'b0000111011110001111111000110000000000000000;
			// PEs: 40 -> 41
			// srcs: (127, 24)(782) 589 --> (782) 589:PENB, pass, NI4
			9'd31 : rdata = 43'b1100011011110000000001001000000000000000000;
			// PEs: 41 -> 41
			// srcs: (128, 99)(1376) 376 --> (1376) 376:NI2, pass, NI2
			9'd32 : rdata = 43'b1100010100010000000001000100000000000000000;
			// PEs: 41, 41 -> 41
			// srcs: (128, 61)(1376) 376, (1377) 2020 --> (1386) 2396:ALU, NI3, +, NI6
			9'd33 : rdata = 43'b0000100111111101000111001100000000000000000;
			// PEs: 40, 41 -> 40
			// srcs: (133, 25)(752) 312, (782) 589 --> (1378) 901:PENB, NI4, +, PEGB0
			9'd34 : rdata = 43'b0000111011110101001000000000000000010000000;
			// PEs: 40 -> 
			// srcs: (135, 26)(1143) 390 --> (1143) 390:PENB, pass, 
			9'd35 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 40, 41 -> 41
			// srcs: (141, 27)(1113) 299, (1143) 390 --> (1403) 689:PENB, ALU, +, NI2
			9'd36 : rdata = 43'b0000111011110001111111000100000000000000000;
			// PEs: 40 -> 
			// srcs: (143, 28)(1203) 527 --> (1203) 527:PENB, pass, 
			9'd37 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 40, 41 -> 41
			// srcs: (149, 29)(1173) 36, (1203) 527 --> (1404) 563:PENB, ALU, +, NI3
			9'd38 : rdata = 43'b0000111011110001111111000110000000000000000;
			// PEs: 40 -> 41
			// srcs: (151, 30)(664) 528 --> (664) 528:PENB, pass, NI4
			9'd39 : rdata = 43'b1100011011110000000001001000000000000000000;
			// PEs: 41 -> 41
			// srcs: (152, 100)(1403) 689 --> (1403) 689:NI2, pass, NI2
			9'd40 : rdata = 43'b1100010100010000000001000100000000000000000;
			// PEs: 41, 41 -> 41
			// srcs: (152, 74)(1403) 689, (1404) 563 --> (1409) 1252:ALU, NI3, +, NI7
			9'd41 : rdata = 43'b0000100111111101000111001110000000000000000;
			// PEs: 40, 41 -> 41
			// srcs: (157, 31)(634) 448, (664) 528 --> (1414) 976:PENB, NI4, +, NI2
			9'd42 : rdata = 43'b0000111011110101001001000100000000000000000;
			// PEs: 40 -> 
			// srcs: (159, 32)(724) 874 --> (724) 874:PENB, pass, 
			9'd43 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 40, 41 -> 41
			// srcs: (165, 33)(694) 960, (724) 874 --> (1415) 1834:PENB, ALU, +, NI3
			9'd44 : rdata = 43'b0000111011110001111111000110000000000000000;
			// PEs: 40 -> 41
			// srcs: (167, 34)(784) -38 --> (784) -38:PENB, pass, NI4
			9'd45 : rdata = 43'b1100011011110000000001001000000000000000000;
			// PEs: 41 -> 41
			// srcs: (168, 101)(1414) 976 --> (1414) 976:NI2, pass, NI2
			9'd46 : rdata = 43'b1100010100010000000001000100000000000000000;
			// PEs: 41, 41 -> 41
			// srcs: (168, 64)(1414) 976, (1415) 1834 --> (1424) 2810:ALU, NI3, +, NI8
			9'd47 : rdata = 43'b0000100111111101000111010000000000000000000;
			// PEs: 40, 41 -> 41
			// srcs: (173, 35)(754) 1176, (784) -38 --> (1416) 1138:PENB, NI4, +, NI2
			9'd48 : rdata = 43'b0000111011110101001001000100000000000000000;
			// PEs: 40 -> 
			// srcs: (175, 36)(844) 160 --> (844) 160:PENB, pass, 
			9'd49 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 40, 41 -> 41
			// srcs: (181, 37)(814) 744, (844) 160 --> (1417) 904:PENB, ALU, +, NI3
			9'd50 : rdata = 43'b0000111011110001111111000110000000000000000;
			// PEs: 40 -> 41
			// srcs: (183, 38)(904) -4 --> (904) -4:PENB, pass, NI4
			9'd51 : rdata = 43'b1100011011110000000001001000000000000000000;
			// PEs: 41 -> 41
			// srcs: (184, 102)(1416) 1138 --> (1416) 1138:NI2, pass, NI2
			9'd52 : rdata = 43'b1100010100010000000001000100000000000000000;
			// PEs: 41, 41 -> 
			// srcs: (184, 65)(1416) 1138, (1417) 904 --> (1425) 2042:ALU, NI3, +, 
			9'd53 : rdata = 43'b0000100111111101000110000000000000000000000;
			// PEs: 41, 41 -> 41
			// srcs: (187, 76)(1424) 2810, (1425) 2042 --> (1429) 4852:NI8, ALU, +, NI2
			9'd54 : rdata = 43'b0000110101000001111111000100000000000000000;
			// PEs: 40, 41 -> 40
			// srcs: (189, 39)(874) 1568, (904) -4 --> (1418) 1564:PENB, NI4, +, PEGB0
			9'd55 : rdata = 43'b0000111011110101001000000000000000010000000;
			// PEs: 40 -> 
			// srcs: (191, 40)(670) 44 --> (670) 44:PENB, pass, 
			9'd56 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 40, 41 -> 41
			// srcs: (197, 41)(640) -28, (670) 44 --> (1528) 16:PENB, ALU, +, NI3
			9'd57 : rdata = 43'b0000111011110001111111000110000000000000000;
			// PEs: 40 -> 
			// srcs: (199, 42)(730) 828 --> (730) 828:PENB, pass, 
			9'd58 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 40, 41 -> 41
			// srcs: (205, 43)(700) 624, (730) 828 --> (1529) 1452:PENB, ALU, +, NI4
			9'd59 : rdata = 43'b0000111011110001111111001000000000000000000;
			// PEs: 40 -> 41
			// srcs: (207, 44)(790) 779 --> (790) 779:PENB, pass, NI8
			9'd60 : rdata = 43'b1100011011110000000001010000000000000000000;
			// PEs: 41 -> 41
			// srcs: (208, 103)(1528) 16 --> (1528) 16:NI3, pass, NI3
			9'd61 : rdata = 43'b1100010100011000000001000110000000000000000;
			// PEs: 41, 41 -> 41
			// srcs: (208, 68)(1528) 16, (1529) 1452 --> (1538) 1468:ALU, NI4, +, NI9
			9'd62 : rdata = 43'b0000100111111101001001010010000000000000000;
			// PEs: 40, 41 -> 41
			// srcs: (213, 45)(760) 600, (790) 779 --> (1530) 1379:PENB, NI8, +, NI3
			9'd63 : rdata = 43'b0000111011110101010001000110000000000000000;
			// PEs: 40 -> 
			// srcs: (215, 46)(850) 480 --> (850) 480:PENB, pass, 
			9'd64 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 40, 41 -> 41
			// srcs: (221, 47)(820) 837, (850) 480 --> (1531) 1317:PENB, ALU, +, NI4
			9'd65 : rdata = 43'b0000111011110001111111001000000000000000000;
			// PEs: 40 -> 41
			// srcs: (223, 48)(910) -2 --> (910) -2:PENB, pass, NI8
			9'd66 : rdata = 43'b1100011011110000000001010000000000000000000;
			// PEs: 41 -> 41
			// srcs: (224, 104)(1530) 1379 --> (1530) 1379:NI3, pass, NI3
			9'd67 : rdata = 43'b1100010100011000000001000110000000000000000;
			// PEs: 41, 41 -> 
			// srcs: (224, 69)(1530) 1379, (1531) 1317 --> (1539) 2696:ALU, NI4, +, 
			9'd68 : rdata = 43'b0000100111111101001000000000000000000000000;
			// PEs: 41, 41 -> 40
			// srcs: (227, 77)(1538) 1468, (1539) 2696 --> (1543) 4164:NI9, ALU, +, PEGB0
			9'd69 : rdata = 43'b0000110101001001111110000000000000010000000;
			// PEs: 40, 41 -> 41
			// srcs: (229, 49)(880) 704, (910) -2 --> (1532) 702:PENB, NI8, +, NI3
			9'd70 : rdata = 43'b0000111011110101010001000110000000000000000;
			// PEs: 40 -> 
			// srcs: (231, 50)(970) 891 --> (970) 891:PENB, pass, 
			9'd71 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 40, 41 -> 41
			// srcs: (237, 51)(940) 348, (970) 891 --> (1533) 1239:PENB, ALU, +, NI4
			9'd72 : rdata = 43'b0000111011110001111111001000000000000000000;
			// PEs: 40 -> 41
			// srcs: (239, 52)(1030) 462 --> (1030) 462:PENB, pass, NI8
			9'd73 : rdata = 43'b1100011011110000000001010000000000000000000;
			// PEs: 41 -> 41
			// srcs: (240, 105)(1532) 702 --> (1532) 702:NI3, pass, NI3
			9'd74 : rdata = 43'b1100010100011000000001000110000000000000000;
			// PEs: 41, 41 -> 41
			// srcs: (240, 70)(1532) 702, (1533) 1239 --> (1540) 1941:ALU, NI4, +, NI9
			9'd75 : rdata = 43'b0000100111111101001001010010000000000000000;
			// PEs: 40, 41 -> 40
			// srcs: (245, 53)(1000) 52, (1030) 462 --> (1534) 514:PENB, NI8, +, PEGB0
			9'd76 : rdata = 43'b0000111011110101010000000000000000010000000;
			// PEs: 40 -> 
			// srcs: (247, 54)(1227) 2387 --> (1227) 2387:PENB, pass, 
			9'd77 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 40, 41 -> 40
			// srcs: (253, 55)(1226) 842, (1227) 2387 --> (1235) 3229:PENB, ALU, +, PEGB0
			9'd78 : rdata = 43'b0000111011110001111110000000000000010000000;
			// PEs: 41 -> 40
			// srcs: (261, 75)(1386) 2396 --> (1386) 2396:NI6, pass, PEGB0
			9'd79 : rdata = 43'b1100010100110000000000000000000000010000000;
			// PEs: 41 -> 40
			// srcs: (269, 83)(1540) 1941 --> (1540) 1941:NI9, pass, PEGB0
			9'd80 : rdata = 43'b1100010101001000000000000000000000010000000;
			// PEs: 40 -> 
			// srcs: (333, 56)(1231) 756 --> (1231) 756:PENB, pass, 
			9'd81 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 40, 41 -> 41
			// srcs: (339, 57)(1230) 554, (1231) 756 --> (1237) 1310:PENB, ALU, +, NI3
			9'd82 : rdata = 43'b0000111011110001111111000110000000000000000;
			// PEs: 40, 41 -> 40
			// srcs: (340, 58)(1283) 1567, (1284) 1750 --> (1292) 3317:PENB, NI0, +, PEGB0
			9'd83 : rdata = 43'b0000111011110101000000000000000000010000000;
			// PEs: 40 -> 
			// srcs: (342, 62)(1402) 1053 --> (1402) 1053:PENB, pass, 
			9'd84 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 40, 41 -> 42
			// srcs: (348, 63)(1401) 690, (1402) 1053 --> (1408) 1743:PENB, ALU, +, PENB
			9'd85 : rdata = 43'b0000111011110001111110000000000000100000000;
			// PEs: 40 -> 41
			// srcs: (350, 66)(1497) 1764 --> (1497) 1764:PENB, pass, NI0
			9'd86 : rdata = 43'b1100011011110000000001000000000000000000000;
			// PEs: 41 -> 40
			// srcs: (351, 84)(1295) 2557 --> (1295) 2557:NI5, pass, PEGB0
			9'd87 : rdata = 43'b1100010100101000000000000000000000010000000;
			// PEs: 40, 41 -> 41
			// srcs: (356, 67)(1496) 990, (1497) 1764 --> (1503) 2754:PENB, NI0, +, NI4
			9'd88 : rdata = 43'b0000111011110101000001001000000000000000000;
			// PEs: 40 -> 41
			// srcs: (358, 71)(1778) 1585 --> (1778) 1585:PENB, pass, NI0
			9'd89 : rdata = 43'b1100011011110000000001000000000000000000000;
			// PEs: 41 -> 40
			// srcs: (360, 86)(1429) 4852 --> (1429) 4852:NI2, pass, PEGB0
			9'd90 : rdata = 43'b1100010100010000000000000000000000010000000;
			// PEs: 40, 41 -> 40
			// srcs: (364, 72)(1777) 1462, (1778) 1585 --> (1786) 3047:PENB, NI0, +, PEGB0
			9'd91 : rdata = 43'b0000111011110101000000000000000000010000000;
			// PEs: 40, 41 -> 40
			// srcs: (473, 78)(1236) 3412, (1237) 1310 --> (1240) 4722:PENB, NI3, +, PEGB0
			9'd92 : rdata = 43'b0000111011110101000110000000000000010000000;
			// PEs: 40 -> 
			// srcs: (475, 80)(1351) 1875 --> (1351) 1875:PENB, pass, 
			9'd93 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 40, 41 -> 41
			// srcs: (481, 81)(1350) 2298, (1351) 1875 --> (1354) 4173:PENB, ALU, +, NI0
			9'd94 : rdata = 43'b0000111011110001111111000000000000000000000;
			// PEs: 40, 41 -> 41
			// srcs: (482, 82)(1502) 732, (1503) 2754 --> (1506) 3486:PENB, NI4, +, NI2
			9'd95 : rdata = 43'b0000111011110101001001000100000000000000000;
			// PEs: 41, 40 -> 42
			// srcs: (483, 85)(1409) 1252, (1410) 4943 --> (1412) 6195:NI7, PENB, +, PENB
			9'd96 : rdata = 43'b0000110100111110111100000000000000100000000;
			// PEs: 41 -> 40
			// srcs: (484, 87)(1297) 5224 --> (1297) 5224:NI1, pass, PEGB0
			9'd97 : rdata = 43'b1100010100001000000000000000000000010000000;
			// PEs: 40 -> 
			// srcs: (1022, 88)(1336) 4389 --> (1336) 4389:PENB, pass, 
			9'd98 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 40, 41 -> 41
			// srcs: (1029, 89)(1335) 4432, (1336) 4389 --> (1337) 8821:PENB, ALU, +, NW0
			9'd99 : rdata = 43'b0000111011110001111110000001000000000000000;
			// PEs: 41, 40 -> 41
			// srcs: (1030, 90)(1354) 4173, (1355) 5478 --> (1356) 9651:NI0, PENB, +, NW1
			9'd100 : rdata = 43'b0000110100000110111100000001000010000000000;
			// PEs: 40 -> 
			// srcs: (1032, 91)(1431) 6812 --> (1431) 6812:PENB, pass, 
			9'd101 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 40, 41 -> 41
			// srcs: (1038, 92)(1430) 5992, (1431) 6812 --> (1432) 12804:PENB, ALU, +, NW2
			9'd102 : rdata = 43'b0000111011110001111110000001000100000000000;
			// PEs: 40 -> 
			// srcs: (1844, 93)(1469) 5610 --> (1469) 5610:PENB, pass, 
			9'd103 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 40, 41 -> 41
			// srcs: (1850, 94)(1468) 3219, (1469) 5610 --> (1470) 8829:PENB, ALU, +, NW3
			9'd104 : rdata = 43'b0000111011110001111110000001000110000000000;
			// PEs: 41, 40 -> 41
			// srcs: (1851, 95)(1506) 3486, (1507) 5409 --> (1508) 8895:NI2, PENB, +, NW4
			9'd105 : rdata = 43'b0000110100010110111100000001001000000000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 42) begin
	always @(*) begin
		case(address)
			// PEs: 40, 41 -> 
			// srcs: (479, 0)(1407) 754, (1408) 1743 --> (1411) 2497:PEGB0, PENB, +, 
			9'd0 : rdata = 43'b0000111100000110111100000000000000000000000;
			// PEs: 42, 41 -> 42
			// srcs: (486, 1)(1411) 2497, (1412) 6195 --> (1413) 8692:ALU, PENB, +, NW0
			9'd1 : rdata = 43'b0000100111111110111100000001000000000000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 43) begin
	always @(*) begin
		case(address)
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 44) begin
	always @(*) begin
		case(address)
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 45) begin
	always @(*) begin
		case(address)
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 46) begin
	always @(*) begin
		case(address)
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 47) begin
	always @(*) begin
		case(address)
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 48) begin
	always @(*) begin
		case(address)
			// PEs: 0 -> 48
			// srcs: (39, 0)(688) 1032 --> (688) 1032:PUGB0, pass, NI0
			9'd0 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 0 -> 49
			// srcs: (40, 1)(718) 1564 --> (718) 1564:PUGB0, pass, PENB
			9'd1 : rdata = 43'b1100011100001000000000000000000000100000000;
			// PEs: 48 -> 49
			// srcs: (46, 2)(688) 1032 --> (688) 1032:NI0, pass, PENB
			9'd2 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 48
			// srcs: (47, 3)(748) 984 --> (748) 984:PUGB0, pass, NI0
			9'd3 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 0 -> 49
			// srcs: (48, 4)(778) 532 --> (778) 532:PUGB0, pass, PENB
			9'd4 : rdata = 43'b1100011100001000000000000000000000100000000;
			// PEs: 48 -> 49
			// srcs: (54, 5)(748) 984 --> (748) 984:NI0, pass, PENB
			9'd5 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 48
			// srcs: (55, 6)(808) -93 --> (808) -93:PUGB0, pass, NI0
			9'd6 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 8 -> 49
			// srcs: (56, 7)(838) 256 --> (838) 256:PUGB1, pass, PENB
			9'd7 : rdata = 43'b1100011100011000000000000000000000100000000;
			// PEs: 48 -> 49
			// srcs: (62, 8)(808) -93 --> (808) -93:NI0, pass, PENB
			9'd8 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 8 -> 48
			// srcs: (63, 9)(868) 32 --> (868) 32:PUGB1, pass, NI0
			9'd9 : rdata = 43'b1100011100011000000001000000000000000000000;
			// PEs: 8 -> 49
			// srcs: (64, 10)(898) -9 --> (898) -9:PUGB1, pass, PENB
			9'd10 : rdata = 43'b1100011100011000000000000000000000100000000;
			// PEs: 48 -> 49
			// srcs: (70, 11)(868) 32 --> (868) 32:NI0, pass, PENB
			9'd11 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 8 -> 48
			// srcs: (71, 12)(928) 29 --> (928) 29:PUGB1, pass, NI0
			9'd12 : rdata = 43'b1100011100011000000001000000000000000000000;
			// PEs: 8 -> 49
			// srcs: (72, 13)(958) 759 --> (958) 759:PUGB1, pass, PENB
			9'd13 : rdata = 43'b1100011100011000000000000000000000100000000;
			// PEs: 48 -> 49
			// srcs: (78, 14)(928) 29 --> (928) 29:NI0, pass, PENB
			9'd14 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 8 -> 48
			// srcs: (79, 15)(988) 18 --> (988) 18:PUGB1, pass, NI0
			9'd15 : rdata = 43'b1100011100011000000001000000000000000000000;
			// PEs: 8 -> 49
			// srcs: (80, 16)(1018) 440 --> (1018) 440:PUGB1, pass, PENB
			9'd16 : rdata = 43'b1100011100011000000000000000000000100000000;
			// PEs: 48 -> 49
			// srcs: (86, 17)(988) 18 --> (988) 18:NI0, pass, PENB
			9'd17 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 8 -> 48
			// srcs: (87, 18)(934) 1131 --> (934) 1131:PUGB1, pass, NI0
			9'd18 : rdata = 43'b1100011100011000000001000000000000000000000;
			// PEs: 8 -> 49
			// srcs: (88, 19)(964) 726 --> (964) 726:PUGB1, pass, PENB
			9'd19 : rdata = 43'b1100011100011000000000000000000000100000000;
			// PEs: 49 -> 56
			// srcs: (93, 58)(1306) 458 --> (1306) 458:PEGB1, pass, PUNB
			9'd20 : rdata = 43'b1100011100010000000000000000000001000000000;
			// PEs: 48 -> 49
			// srcs: (94, 20)(934) 1131 --> (934) 1131:NI0, pass, PENB
			9'd21 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 8 -> 48
			// srcs: (95, 21)(994) 22 --> (994) 22:PUGB1, pass, NI0
			9'd22 : rdata = 43'b1100011100011000000001000000000000000000000;
			// PEs: 8 -> 49
			// srcs: (96, 22)(1024) 836 --> (1024) 836:PUGB1, pass, PENB
			9'd23 : rdata = 43'b1100011100011000000000000000000000100000000;
			// PEs: 48 -> 49
			// srcs: (102, 23)(994) 22 --> (994) 22:NI0, pass, PENB
			9'd24 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 48
			// srcs: (103, 24)(635) 434 --> (635) 434:PUGB0, pass, NI0
			9'd25 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 0 -> 49
			// srcs: (104, 25)(665) 429 --> (665) 429:PUGB0, pass, PENB
			9'd26 : rdata = 43'b1100011100001000000000000000000000100000000;
			// PEs: 49 -> 24
			// srcs: (109, 63)(1420) 858 --> (1420) 858:PEGB1, pass, PUGB3
			9'd27 : rdata = 43'b1100011100010000000000000000000000000001011;
			// PEs: 48 -> 49
			// srcs: (110, 26)(635) 434 --> (635) 434:NI0, pass, PENB
			9'd28 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 48
			// srcs: (111, 27)(695) 336 --> (695) 336:PUGB0, pass, NI0
			9'd29 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 0 -> 49
			// srcs: (112, 28)(725) 184 --> (725) 184:PUGB0, pass, PENB
			9'd30 : rdata = 43'b1100011100001000000000000000000000100000000;
			// PEs: 48 -> 49
			// srcs: (118, 29)(695) 336 --> (695) 336:NI0, pass, PENB
			9'd31 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 48
			// srcs: (119, 30)(755) -24 --> (755) -24:PUGB0, pass, NI0
			9'd32 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 0 -> 49
			// srcs: (120, 31)(785) 304 --> (785) 304:PUGB0, pass, PENB
			9'd33 : rdata = 43'b1100011100001000000000000000000000100000000;
			// PEs: 48 -> 49
			// srcs: (126, 32)(755) -24 --> (755) -24:NI0, pass, PENB
			9'd34 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 48
			// srcs: (128, 33)(641) 112 --> (641) 112:PUGB0, pass, NI0
			9'd35 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 0 -> 49
			// srcs: (129, 34)(671) 242 --> (671) 242:PUGB0, pass, PENB
			9'd36 : rdata = 43'b1100011100001000000000000000000000100000000;
			// PEs: 49 -> 56
			// srcs: (133, 64)(1435) 280 --> (1435) 280:PEGB1, pass, PUNB
			9'd37 : rdata = 43'b1100011100010000000000000000000001000000000;
			// PEs: 48 -> 49
			// srcs: (135, 35)(641) 112 --> (641) 112:NI0, pass, PENB
			9'd38 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 48
			// srcs: (136, 36)(701) -72 --> (701) -72:PUGB0, pass, NI0
			9'd39 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 0 -> 49
			// srcs: (137, 37)(731) -92 --> (731) -92:PUGB0, pass, PENB
			9'd40 : rdata = 43'b1100011100001000000000000000000000100000000;
			// PEs: 48 -> 49
			// srcs: (143, 38)(701) -72 --> (701) -72:NI0, pass, PENB
			9'd41 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 48
			// srcs: (144, 39)(761) 672 --> (761) 672:PUGB0, pass, NI0
			9'd42 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 0 -> 49
			// srcs: (145, 40)(791) 722 --> (791) 722:PUGB0, pass, PENB
			9'd43 : rdata = 43'b1100011100001000000000000000000000100000000;
			// PEs: 48 -> 49
			// srcs: (151, 41)(761) 672 --> (761) 672:NI0, pass, PENB
			9'd44 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 48
			// srcs: (152, 42)(821) 837 --> (821) 837:PUGB0, pass, NI0
			9'd45 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 8 -> 49
			// srcs: (153, 43)(851) 320 --> (851) 320:PUGB1, pass, PENB
			9'd46 : rdata = 43'b1100011100011000000000000000000000100000000;
			// PEs: 48 -> 49
			// srcs: (159, 44)(821) 837 --> (821) 837:NI0, pass, PENB
			9'd47 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 8 -> 48
			// srcs: (160, 45)(881) 224 --> (881) 224:PUGB1, pass, NI0
			9'd48 : rdata = 43'b1100011100011000000001000000000000000000000;
			// PEs: 8 -> 49
			// srcs: (161, 46)(911) -14 --> (911) -14:PUGB1, pass, PENB
			9'd49 : rdata = 43'b1100011100011000000000000000000000100000000;
			// PEs: 48 -> 49
			// srcs: (167, 47)(881) 224 --> (881) 224:NI0, pass, PENB
			9'd50 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 8 -> 48
			// srcs: (168, 48)(941) 1334 --> (941) 1334:PUGB1, pass, NI0
			9'd51 : rdata = 43'b1100011100011000000001000000000000000000000;
			// PEs: 8 -> 49
			// srcs: (169, 49)(971) 1584 --> (971) 1584:PUGB1, pass, PENB
			9'd52 : rdata = 43'b1100011100011000000000000000000000100000000;
			// PEs: 48 -> 49
			// srcs: (175, 50)(941) 1334 --> (941) 1334:NI0, pass, PENB
			9'd53 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 8 -> 48
			// srcs: (176, 51)(1001) 30 --> (1001) 30:PUGB1, pass, NI0
			9'd54 : rdata = 43'b1100011100011000000001000000000000000000000;
			// PEs: 8 -> 49
			// srcs: (177, 52)(1031) -44 --> (1031) -44:PUGB1, pass, PENB
			9'd55 : rdata = 43'b1100011100011000000000000000000000100000000;
			// PEs: 48 -> 49
			// srcs: (183, 53)(1001) 30 --> (1001) 30:NI0, pass, PENB
			9'd56 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 24 -> 48
			// srcs: (184, 54)(1224) 95 --> (1224) 95:PUGB3, pass, NI0
			9'd57 : rdata = 43'b1100011100111000000001000000000000000000000;
			// PEs: 32 -> 49
			// srcs: (185, 55)(1225) 3148 --> (1225) 3148:PUGB4, pass, PENB
			9'd58 : rdata = 43'b1100011101001000000000000000000000100000000;
			// PEs: 49 -> 56
			// srcs: (190, 68)(1553) -14 --> (1553) -14:PEGB1, pass, PUNB
			9'd59 : rdata = 43'b1100011100010000000000000000000001000000000;
			// PEs: 48 -> 49
			// srcs: (191, 56)(1224) 95 --> (1224) 95:NI0, pass, PENB
			9'd60 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 40 -> 49
			// srcs: (192, 57)(1300) 644 --> (1300) 644:PUNB, pass, PENB
			9'd61 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 40 -> 48
			// srcs: (193, 59)(1378) 901 --> (1378) 901:PUNB, pass, NI0
			9'd62 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 16 -> 49
			// srcs: (194, 60)(1379) 1873 --> (1379) 1873:PUGB2, pass, PENB
			9'd63 : rdata = 43'b1100011100101000000000000000000000100000000;
			// PEs: 48 -> 49
			// srcs: (200, 61)(1378) 901 --> (1378) 901:NI0, pass, PENB
			9'd64 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 40 -> 49
			// srcs: (201, 62)(1418) 1564 --> (1418) 1564:PUNB, pass, PENB
			9'd65 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 49 -> 8
			// srcs: (202, 80)(1315) 4919 --> (1315) 4919:PEGB1, pass, PUGB1
			9'd66 : rdata = 43'b1100011100010000000000000000000000000001001;
			// PEs: 49 -> 56
			// srcs: (203, 71)(1443) 1383 --> (1443) 1383:PEGB1, pass, PUNB
			9'd67 : rdata = 43'b1100011100010000000000000000000001000000000;
			// PEs: 49 -> 56
			// srcs: (211, 72)(1312) 811 --> (1312) 811:PEGB1, pass, PUNB
			9'd68 : rdata = 43'b1100011100010000000000000000000001000000000;
			// PEs: 49 -> 56
			// srcs: (219, 78)(1559) 3128 --> (1559) 3128:PEGB1, pass, PUNB
			9'd69 : rdata = 43'b1100011100010000000000000000000001000000000;
			// PEs: 50 -> 56
			// srcs: (220, 82)(1562) 2741 --> (1562) 2741:PEGB2, pass, PUNB
			9'd70 : rdata = 43'b1100011100100000000000000000000001000000000;
			// PEs: 40 -> 48
			// srcs: (252, 65)(1534) 514 --> (1534) 514:PUNB, pass, NI0
			9'd71 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 24 -> 49
			// srcs: (430, 66)(1535) 1308 --> (1535) 1308:PUGB3, pass, PENB
			9'd72 : rdata = 43'b1100011100111000000000000000000000100000000;
			// PEs: 48 -> 49
			// srcs: (437, 67)(1534) 514 --> (1534) 514:NI0, pass, PENB
			9'd73 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 40 -> 49
			// srcs: (438, 69)(1235) 3229 --> (1235) 3229:PUNB, pass, PENB
			9'd74 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 40 -> 49
			// srcs: (439, 70)(1386) 2396 --> (1386) 2396:PUNB, pass, PENB
			9'd75 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 49 -> 0
			// srcs: (445, 79)(1239) 6472 --> (1239) 6472:PEGB1, pass, PUGB0
			9'd76 : rdata = 43'b1100011100010000000000000000000000000001000;
			// PEs: 49 -> 8
			// srcs: (446, 81)(1391) 5170 --> (1391) 5170:PEGB1, pass, PUGB1
			9'd77 : rdata = 43'b1100011100010000000000000000000000000001001;
			// PEs: 24 -> 49
			// srcs: (546, 73)(1427) 2571 --> (1427) 2571:PUGB3, pass, PENB
			9'd78 : rdata = 43'b1100011100111000000000000000000000100000000;
			// PEs: 56 -> 48
			// srcs: (547, 74)(1445) 2446 --> (1445) 2446:PUGB7, pass, NI0
			9'd79 : rdata = 43'b1100011101111000000001000000000000000000000;
			// PEs: 32 -> 49
			// srcs: (548, 75)(1446) 1940 --> (1446) 1940:PUGB4, pass, PENB
			9'd80 : rdata = 43'b1100011101001000000000000000000000100000000;
			// PEs: 48 -> 49
			// srcs: (554, 76)(1445) 2446 --> (1445) 2446:NI0, pass, PENB
			9'd81 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 40 -> 49
			// srcs: (555, 77)(1540) 1941 --> (1540) 1941:PUNB, pass, PENB
			9'd82 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 49 -> 40
			// srcs: (556, 83)(1430) 5992 --> (1430) 5992:PEGB1, pass, PUGB5
			9'd83 : rdata = 43'b1100011100010000000000000000000000000001101;
			// PEs: 32 -> 48
			// srcs: (557, 85)(1525) 2228 --> (1525) 2228:PUGB4, pass, NI0
			9'd84 : rdata = 43'b1100011101001000000001000000000000000000000;
			// PEs: 49 -> 56
			// srcs: (561, 84)(1449) 4386 --> (1449) 4386:PEGB1, pass, PUNB
			9'd85 : rdata = 43'b1100011100010000000000000000000001000000000;
			// PEs: 16 -> 49
			// srcs: (1032, 86)(1526) 6573 --> (1526) 6573:PUGB2, pass, PENB
			9'd86 : rdata = 43'b1100011100101000000000000000000000100000000;
			// PEs: 48 -> 49
			// srcs: (1038, 87)(1525) 2228 --> (1525) 2228:NI0, pass, PENB
			9'd87 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 16 -> 49
			// srcs: (1039, 88)(1545) 6630 --> (1545) 6630:PUGB2, pass, PENB
			9'd88 : rdata = 43'b1100011100101000000000000000000000100000000;
			// PEs: 0 -> 48
			// srcs: (1040, 89)(1582) 4313 --> (1582) 4313:PUGB0, pass, NI0
			9'd89 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 16 -> 49
			// srcs: (1044, 90)(1583) 8760 --> (1583) 8760:PUGB2, pass, PENB
			9'd90 : rdata = 43'b1100011100101000000000000000000000100000000;
			// PEs: 48 -> 49
			// srcs: (1051, 91)(1582) 4313 --> (1582) 4313:NI0, pass, PENB
			9'd91 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 16 -> 48
			// srcs: (1052, 92)(1620) 2914 --> (1620) 2914:PUGB2, pass, NI0
			9'd92 : rdata = 43'b1100011100101000000001000000000000000000000;
			// PEs: 32 -> 49
			// srcs: (1053, 93)(1621) 5293 --> (1621) 5293:PUGB4, pass, PENB
			9'd93 : rdata = 43'b1100011101001000000000000000000000100000000;
			// PEs: 48 -> 49
			// srcs: (1059, 94)(1620) 2914 --> (1620) 2914:NI0, pass, PENB
			9'd94 : rdata = 43'b1100010100000000000000000000000000100000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 49) begin
	always @(*) begin
		case(address)
			// PEs: 48 -> 
			// srcs: (42, 0)(718) 1564 --> (718) 1564:PENB, pass, 
			9'd0 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 48, 49 -> 49
			// srcs: (48, 1)(688) 1032, (718) 1564 --> (1301) 2596:PENB, ALU, +, NI0
			9'd1 : rdata = 43'b0000111011110001111111000000000000000000000;
			// PEs: 48 -> 
			// srcs: (50, 2)(778) 532 --> (778) 532:PENB, pass, 
			9'd2 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 48, 49 -> 49
			// srcs: (56, 3)(748) 984, (778) 532 --> (1302) 1516:PENB, ALU, +, NI1
			9'd3 : rdata = 43'b0000111011110001111111000010000000000000000;
			// PEs: 48 -> 
			// srcs: (58, 4)(838) 256 --> (838) 256:PENB, pass, 
			9'd4 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 48, 49 -> 49
			// srcs: (64, 5)(808) -93, (838) 256 --> (1303) 163:PENB, ALU, +, NI2
			9'd5 : rdata = 43'b0000111011110001111111000100000000000000000;
			// PEs: 48 -> 49
			// srcs: (66, 6)(898) -9 --> (898) -9:PENB, pass, NI3
			9'd6 : rdata = 43'b1100011011110000000001000110000000000000000;
			// PEs: 49 -> 49
			// srcs: (67, 68)(1302) 1516 --> (1302) 1516:NI1, pass, NI1
			9'd7 : rdata = 43'b1100010100001000000001000010000000000000000;
			// PEs: 49, 49 -> 49
			// srcs: (67, 39)(1302) 1516, (1303) 163 --> (1311) 1679:ALU, NI2, +, NI4
			9'd8 : rdata = 43'b0000100111111101000101001000000000000000000;
			// PEs: 48, 49 -> 49
			// srcs: (72, 7)(868) 32, (898) -9 --> (1304) 23:PENB, NI3, +, NI1
			9'd9 : rdata = 43'b0000111011110101000111000010000000000000000;
			// PEs: 48 -> 
			// srcs: (74, 8)(958) 759 --> (958) 759:PENB, pass, 
			9'd10 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 48, 49 -> 49
			// srcs: (80, 9)(928) 29, (958) 759 --> (1305) 788:PENB, ALU, +, NI2
			9'd11 : rdata = 43'b0000111011110001111111000100000000000000000;
			// PEs: 48 -> 49
			// srcs: (82, 10)(1018) 440 --> (1018) 440:PENB, pass, NI3
			9'd12 : rdata = 43'b1100011011110000000001000110000000000000000;
			// PEs: 49 -> 49
			// srcs: (83, 69)(1304) 23 --> (1304) 23:NI1, pass, NI1
			9'd13 : rdata = 43'b1100010100001000000001000010000000000000000;
			// PEs: 49, 49 -> 49
			// srcs: (83, 40)(1304) 23, (1305) 788 --> (1312) 811:ALU, NI2, +, NI5
			9'd14 : rdata = 43'b0000100111111101000101001010000000000000000;
			// PEs: 48, 49 -> 48
			// srcs: (88, 11)(988) 18, (1018) 440 --> (1306) 458:PENB, NI3, +, PEGB0
			9'd15 : rdata = 43'b0000111011110101000110000000000000010000000;
			// PEs: 48 -> 
			// srcs: (90, 12)(964) 726 --> (964) 726:PENB, pass, 
			9'd16 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 48, 49 -> 49
			// srcs: (96, 13)(934) 1131, (964) 726 --> (1419) 1857:PENB, ALU, +, NI1
			9'd17 : rdata = 43'b0000111011110001111111000010000000000000000;
			// PEs: 48 -> 
			// srcs: (98, 14)(1024) 836 --> (1024) 836:PENB, pass, 
			9'd18 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 48, 49 -> 48
			// srcs: (104, 15)(994) 22, (1024) 836 --> (1420) 858:PENB, ALU, +, PEGB0
			9'd19 : rdata = 43'b0000111011110001111110000000000000010000000;
			// PEs: 48 -> 
			// srcs: (106, 16)(665) 429 --> (665) 429:PENB, pass, 
			9'd20 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 48, 49 -> 49
			// srcs: (112, 17)(635) 434, (665) 429 --> (1433) 863:PENB, ALU, +, NI2
			9'd21 : rdata = 43'b0000111011110001111111000100000000000000000;
			// PEs: 48 -> 
			// srcs: (114, 18)(725) 184 --> (725) 184:PENB, pass, 
			9'd22 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 48, 49 -> 49
			// srcs: (120, 19)(695) 336, (725) 184 --> (1434) 520:PENB, ALU, +, NI3
			9'd23 : rdata = 43'b0000111011110001111111000110000000000000000;
			// PEs: 48 -> 49
			// srcs: (122, 20)(785) 304 --> (785) 304:PENB, pass, NI6
			9'd24 : rdata = 43'b1100011011110000000001001100000000000000000;
			// PEs: 49 -> 49
			// srcs: (123, 70)(1433) 863 --> (1433) 863:NI2, pass, NI2
			9'd25 : rdata = 43'b1100010100010000000001000100000000000000000;
			// PEs: 49, 49 -> 49
			// srcs: (123, 44)(1433) 863, (1434) 520 --> (1443) 1383:ALU, NI3, +, NI7
			9'd26 : rdata = 43'b0000100111111101000111001110000000000000000;
			// PEs: 48, 49 -> 48
			// srcs: (128, 21)(755) -24, (785) 304 --> (1435) 280:PENB, NI6, +, PEGB0
			9'd27 : rdata = 43'b0000111011110101001100000000000000010000000;
			// PEs: 48 -> 
			// srcs: (131, 22)(671) 242 --> (671) 242:PENB, pass, 
			9'd28 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 48, 49 -> 49
			// srcs: (137, 23)(641) 112, (671) 242 --> (1547) 354:PENB, ALU, +, NI2
			9'd29 : rdata = 43'b0000111011110001111111000100000000000000000;
			// PEs: 48 -> 
			// srcs: (139, 24)(731) -92 --> (731) -92:PENB, pass, 
			9'd30 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 48, 49 -> 49
			// srcs: (145, 25)(701) -72, (731) -92 --> (1548) -164:PENB, ALU, +, NI3
			9'd31 : rdata = 43'b0000111011110001111111000110000000000000000;
			// PEs: 48 -> 49
			// srcs: (147, 26)(791) 722 --> (791) 722:PENB, pass, NI6
			9'd32 : rdata = 43'b1100011011110000000001001100000000000000000;
			// PEs: 49 -> 49
			// srcs: (148, 71)(1547) 354 --> (1547) 354:NI2, pass, NI2
			9'd33 : rdata = 43'b1100010100010000000001000100000000000000000;
			// PEs: 49, 49 -> 49
			// srcs: (148, 47)(1547) 354, (1548) -164 --> (1557) 190:ALU, NI3, +, NI8
			9'd34 : rdata = 43'b0000100111111101000111010000000000000000000;
			// PEs: 48, 49 -> 49
			// srcs: (153, 27)(761) 672, (791) 722 --> (1549) 1394:PENB, NI6, +, NI2
			9'd35 : rdata = 43'b0000111011110101001101000100000000000000000;
			// PEs: 48 -> 
			// srcs: (155, 28)(851) 320 --> (851) 320:PENB, pass, 
			9'd36 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 48, 49 -> 50
			// srcs: (161, 29)(821) 837, (851) 320 --> (1550) 1157:PENB, ALU, +, PENB
			9'd37 : rdata = 43'b0000111011110001111110000000000000100000000;
			// PEs: 48 -> 49
			// srcs: (163, 30)(911) -14 --> (911) -14:PENB, pass, NI3
			9'd38 : rdata = 43'b1100011011110000000001000110000000000000000;
			// PEs: 49 -> 50
			// srcs: (168, 48)(1549) 1394 --> (1549) 1394:NI2, pass, PENB
			9'd39 : rdata = 43'b1100010100010000000000000000000000100000000;
			// PEs: 48, 49 -> 49
			// srcs: (169, 31)(881) 224, (911) -14 --> (1551) 210:PENB, NI3, +, NI2
			9'd40 : rdata = 43'b0000111011110101000111000100000000000000000;
			// PEs: 48 -> 49
			// srcs: (171, 32)(971) 1584 --> (971) 1584:PENB, pass, NI3
			9'd41 : rdata = 43'b1100011011110000000001000110000000000000000;
			// PEs: 49 -> 50
			// srcs: (175, 54)(1557) 190 --> (1557) 190:NI8, pass, PENB
			9'd42 : rdata = 43'b1100010101000000000000000000000000100000000;
			// PEs: 48, 49 -> 49
			// srcs: (177, 33)(941) 1334, (971) 1584 --> (1552) 2918:PENB, NI3, +, NI6
			9'd43 : rdata = 43'b0000111011110101000111001100000000000000000;
			// PEs: 48 -> 49
			// srcs: (179, 34)(1031) -44 --> (1031) -44:PENB, pass, NI3
			9'd44 : rdata = 43'b1100011011110000000001000110000000000000000;
			// PEs: 49 -> 49
			// srcs: (180, 72)(1551) 210 --> (1551) 210:NI2, pass, NI2
			9'd45 : rdata = 43'b1100010100010000000001000100000000000000000;
			// PEs: 49, 49 -> 49
			// srcs: (180, 49)(1551) 210, (1552) 2918 --> (1559) 3128:ALU, NI6, +, NI8
			9'd46 : rdata = 43'b0000100111111101001101010000000000000000000;
			// PEs: 48, 49 -> 48
			// srcs: (185, 35)(1001) 30, (1031) -44 --> (1553) -14:PENB, NI3, +, PEGB0
			9'd47 : rdata = 43'b0000111011110101000110000000000000010000000;
			// PEs: 48 -> 
			// srcs: (187, 36)(1225) 3148 --> (1225) 3148:PENB, pass, 
			9'd48 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 48, 49 -> 49
			// srcs: (193, 37)(1224) 95, (1225) 3148 --> (1234) 3243:PENB, ALU, +, NI2
			9'd49 : rdata = 43'b0000111011110001111111000100000000000000000;
			// PEs: 48, 49 -> 49
			// srcs: (194, 38)(1300) 644, (1301) 2596 --> (1310) 3240:PENB, NI0, +, NI3
			9'd50 : rdata = 43'b0000111011110101000001000110000000000000000;
			// PEs: 48 -> 49
			// srcs: (196, 41)(1379) 1873 --> (1379) 1873:PENB, pass, NI0
			9'd51 : rdata = 43'b1100011011110000000001000000000000000000000;
			// PEs: 49 -> 49
			// srcs: (197, 73)(1310) 3240 --> (1310) 3240:NI3, pass, NI3
			9'd52 : rdata = 43'b1100010100011000000001000110000000000000000;
			// PEs: 49, 49 -> 48
			// srcs: (197, 51)(1310) 3240, (1311) 1679 --> (1315) 4919:ALU, NI4, +, PEGB0
			9'd53 : rdata = 43'b0000100111111101001000000000000000010000000;
			// PEs: 49 -> 48
			// srcs: (198, 53)(1443) 1383 --> (1443) 1383:NI7, pass, PEGB0
			9'd54 : rdata = 43'b1100010100111000000000000000000000010000000;
			// PEs: 48, 49 -> 49
			// srcs: (202, 42)(1378) 901, (1379) 1873 --> (1387) 2774:PENB, NI0, +, NI3
			9'd55 : rdata = 43'b0000111011110101000001000110000000000000000;
			// PEs: 48, 49 -> 49
			// srcs: (203, 43)(1418) 1564, (1419) 1857 --> (1426) 3421:PENB, NI1, +, NI0
			9'd56 : rdata = 43'b0000111011110101000011000000000000000000000;
			// PEs: 49 -> 48
			// srcs: (206, 55)(1312) 811 --> (1312) 811:NI5, pass, PEGB0
			9'd57 : rdata = 43'b1100010100101000000000000000000000010000000;
			// PEs: 49 -> 48
			// srcs: (214, 60)(1559) 3128 --> (1559) 3128:NI8, pass, PEGB0
			9'd58 : rdata = 43'b1100010101000000000000000000000000010000000;
			// PEs: 48 -> 
			// srcs: (432, 45)(1535) 1308 --> (1535) 1308:PENB, pass, 
			9'd59 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 48, 49 -> 49
			// srcs: (439, 46)(1534) 514, (1535) 1308 --> (1541) 1822:PENB, ALU, +, NI1
			9'd60 : rdata = 43'b0000111011110001111111000010000000000000000;
			// PEs: 49, 48 -> 48
			// srcs: (440, 50)(1234) 3243, (1235) 3229 --> (1239) 6472:NI2, PENB, +, PEGB0
			9'd61 : rdata = 43'b0000110100010110111100000000000000010000000;
			// PEs: 48, 49 -> 48
			// srcs: (441, 52)(1386) 2396, (1387) 2774 --> (1391) 5170:PENB, NI3, +, PEGB0
			9'd62 : rdata = 43'b0000111011110101000110000000000000010000000;
			// PEs: 49, 48 -> 48
			// srcs: (549, 56)(1426) 3421, (1427) 2571 --> (1430) 5992:NI0, PENB, +, PEGB0
			9'd63 : rdata = 43'b0000110100000110111100000000000000010000000;
			// PEs: 48 -> 
			// srcs: (550, 57)(1446) 1940 --> (1446) 1940:PENB, pass, 
			9'd64 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 48, 49 -> 48
			// srcs: (556, 58)(1445) 2446, (1446) 1940 --> (1449) 4386:PENB, ALU, +, PEGB0
			9'd65 : rdata = 43'b0000111011110001111110000000000000010000000;
			// PEs: 48, 49 -> 49
			// srcs: (557, 59)(1540) 1941, (1541) 1822 --> (1544) 3763:PENB, NI1, +, NI0
			9'd66 : rdata = 43'b0000111011110101000011000000000000000000000;
			// PEs: 48 -> 
			// srcs: (1034, 61)(1526) 6573 --> (1526) 6573:PENB, pass, 
			9'd67 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 48, 49 -> 49
			// srcs: (1040, 62)(1525) 2228, (1526) 6573 --> (1527) 8801:PENB, ALU, +, NW0
			9'd68 : rdata = 43'b0000111011110001111110000001000000000000000;
			// PEs: 49, 48 -> 49
			// srcs: (1041, 63)(1544) 3763, (1545) 6630 --> (1546) 10393:NI0, PENB, +, NW1
			9'd69 : rdata = 43'b0000110100000110111100000001000010000000000;
			// PEs: 48 -> 
			// srcs: (1046, 64)(1583) 8760 --> (1583) 8760:PENB, pass, 
			9'd70 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 48, 49 -> 49
			// srcs: (1053, 65)(1582) 4313, (1583) 8760 --> (1584) 13073:PENB, ALU, +, NW2
			9'd71 : rdata = 43'b0000111011110001111110000001000100000000000;
			// PEs: 48 -> 
			// srcs: (1055, 66)(1621) 5293 --> (1621) 5293:PENB, pass, 
			9'd72 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 48, 49 -> 49
			// srcs: (1061, 67)(1620) 2914, (1621) 5293 --> (1622) 8207:PENB, ALU, +, NW3
			9'd73 : rdata = 43'b0000111011110001111110000001000110000000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 50) begin
	always @(*) begin
		case(address)
			// PEs: 49 -> 
			// srcs: (163, 0)(1550) 1157 --> (1550) 1157:PENB, pass, 
			9'd0 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 49, 50 -> 
			// srcs: (170, 1)(1549) 1394, (1550) 1157 --> (1558) 2551:PENB, ALU, +, 
			9'd1 : rdata = 43'b0000111011110001111110000000000000000000000;
			// PEs: 49, 50 -> 48
			// srcs: (177, 2)(1557) 190, (1558) 2551 --> (1562) 2741:PENB, ALU, +, PEGB0
			9'd2 : rdata = 43'b0000111011110001111110000000000000010000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 51) begin
	always @(*) begin
		case(address)
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 52) begin
	always @(*) begin
		case(address)
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 53) begin
	always @(*) begin
		case(address)
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 54) begin
	always @(*) begin
		case(address)
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 55) begin
	always @(*) begin
		case(address)
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 56) begin
	always @(*) begin
		case(address)
			// PEs: 0 -> 56
			// srcs: (44, 0)(629) 630 --> (629) 630:PUGB0, pass, NI0
			9'd0 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 0 -> 57
			// srcs: (45, 1)(659) 22 --> (659) 22:PUGB0, pass, PENB
			9'd1 : rdata = 43'b1100011100001000000000000000000000100000000;
			// PEs: 56 -> 57
			// srcs: (51, 2)(629) 630 --> (629) 630:NI0, pass, PENB
			9'd2 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 56
			// srcs: (52, 3)(689) 600 --> (689) 600:PUGB0, pass, NI0
			9'd3 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 0 -> 57
			// srcs: (53, 4)(719) 1104 --> (719) 1104:PUGB0, pass, PENB
			9'd4 : rdata = 43'b1100011100001000000000000000000000100000000;
			// PEs: 56 -> 57
			// srcs: (59, 5)(689) 600 --> (689) 600:NI0, pass, PENB
			9'd5 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 56
			// srcs: (60, 6)(749) 360 --> (749) 360:PUGB0, pass, NI0
			9'd6 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 0 -> 57
			// srcs: (61, 7)(779) 95 --> (779) 95:PUGB0, pass, PENB
			9'd7 : rdata = 43'b1100011100001000000000000000000000100000000;
			// PEs: 56 -> 57
			// srcs: (67, 8)(749) 360 --> (749) 360:NI0, pass, PENB
			9'd8 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 56
			// srcs: (68, 9)(809) 310 --> (809) 310:PUGB0, pass, NI0
			9'd9 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 8 -> 57
			// srcs: (69, 10)(839) 736 --> (839) 736:PUGB1, pass, PENB
			9'd10 : rdata = 43'b1100011100011000000000000000000000100000000;
			// PEs: 56 -> 57
			// srcs: (75, 11)(809) 310 --> (809) 310:NI0, pass, PENB
			9'd11 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 8 -> 56
			// srcs: (76, 12)(869) 704 --> (869) 704:PUGB1, pass, NI0
			9'd12 : rdata = 43'b1100011100011000000001000000000000000000000;
			// PEs: 8 -> 57
			// srcs: (77, 13)(899) -4 --> (899) -4:PUGB1, pass, PENB
			9'd13 : rdata = 43'b1100011100011000000000000000000000100000000;
			// PEs: 56 -> 57
			// srcs: (83, 14)(869) 704 --> (869) 704:NI0, pass, PENB
			9'd14 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 8 -> 56
			// srcs: (84, 15)(929) 1015 --> (929) 1015:PUGB1, pass, NI0
			9'd15 : rdata = 43'b1100011100011000000001000000000000000000000;
			// PEs: 8 -> 57
			// srcs: (85, 16)(959) 990 --> (959) 990:PUGB1, pass, PENB
			9'd16 : rdata = 43'b1100011100011000000000000000000000100000000;
			// PEs: 57 -> 16
			// srcs: (88, 90)(1334) 3857 --> (1334) 3857:PEGB1, pass, PUGB2
			9'd17 : rdata = 43'b1100011100010000000000000000000000000001010;
			// PEs: 56 -> 57
			// srcs: (91, 17)(929) 1015 --> (929) 1015:NI0, pass, PENB
			9'd18 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 8 -> 56
			// srcs: (92, 18)(989) 90 --> (989) 90:PUGB1, pass, NI0
			9'd19 : rdata = 43'b1100011100011000000001000000000000000000000;
			// PEs: 8 -> 57
			// srcs: (93, 19)(1019) 506 --> (1019) 506:PUGB1, pass, PENB
			9'd20 : rdata = 43'b1100011100011000000000000000000000100000000;
			// PEs: 56 -> 57
			// srcs: (99, 20)(989) 90 --> (989) 90:NI0, pass, PENB
			9'd21 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 56
			// srcs: (100, 21)(815) 1054 --> (815) 1054:PUGB0, pass, NI0
			9'd22 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 8 -> 57
			// srcs: (101, 22)(845) 672 --> (845) 672:PUGB1, pass, PENB
			9'd23 : rdata = 43'b1100011100011000000000000000000000100000000;
			// PEs: 57 -> 0
			// srcs: (106, 75)(1325) 596 --> (1325) 596:PEGB1, pass, PUNB
			9'd24 : rdata = 43'b1100011100010000000000000000000001000000000;
			// PEs: 56 -> 57
			// srcs: (107, 23)(815) 1054 --> (815) 1054:NI0, pass, PENB
			9'd25 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 8 -> 56
			// srcs: (108, 24)(875) 1536 --> (875) 1536:PUGB1, pass, NI0
			9'd26 : rdata = 43'b1100011100011000000001000000000000000000000;
			// PEs: 8 -> 57
			// srcs: (109, 25)(905) -35 --> (905) -35:PUGB1, pass, PENB
			9'd27 : rdata = 43'b1100011100011000000000000000000000100000000;
			// PEs: 56 -> 57
			// srcs: (115, 26)(875) 1536 --> (875) 1536:NI0, pass, PENB
			9'd28 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 8 -> 56
			// srcs: (116, 27)(935) 1044 --> (935) 1044:PUGB1, pass, NI0
			9'd29 : rdata = 43'b1100011100011000000001000000000000000000000;
			// PEs: 8 -> 57
			// srcs: (117, 28)(965) -99 --> (965) -99:PUGB1, pass, PENB
			9'd30 : rdata = 43'b1100011100011000000000000000000000100000000;
			// PEs: 56 -> 57
			// srcs: (123, 29)(935) 1044 --> (935) 1044:NI0, pass, PENB
			9'd31 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 8 -> 56
			// srcs: (124, 30)(995) 60 --> (995) 60:PUGB1, pass, NI0
			9'd32 : rdata = 43'b1100011100011000000001000000000000000000000;
			// PEs: 8 -> 57
			// srcs: (125, 31)(1025) 308 --> (1025) 308:PUGB1, pass, PENB
			9'd33 : rdata = 43'b1100011100011000000000000000000000100000000;
			// PEs: 56 -> 57
			// srcs: (131, 32)(995) 60 --> (995) 60:NI0, pass, PENB
			9'd34 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 16 -> 56
			// srcs: (132, 33)(1115) 69 --> (1115) 69:PUGB2, pass, NI0
			9'd35 : rdata = 43'b1100011100101000000001000000000000000000000;
			// PEs: 16 -> 57
			// srcs: (133, 34)(1145) 312 --> (1145) 312:PUGB2, pass, PENB
			9'd36 : rdata = 43'b1100011100101000000000000000000000100000000;
			// PEs: 57 -> 48
			// srcs: (134, 87)(1445) 2446 --> (1445) 2446:PEGB1, pass, PUGB6
			9'd37 : rdata = 43'b1100011100010000000000000000000000000001110;
			// PEs: 57 -> 32
			// srcs: (138, 77)(1439) 368 --> (1439) 368:PEGB1, pass, PUGB4
			9'd38 : rdata = 43'b1100011100010000000000000000000000000001100;
			// PEs: 56 -> 57
			// srcs: (139, 35)(1115) 69 --> (1115) 69:NI0, pass, PENB
			9'd39 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 16 -> 56
			// srcs: (140, 36)(1175) 198 --> (1175) 198:PUGB2, pass, NI0
			9'd40 : rdata = 43'b1100011100101000000001000000000000000000000;
			// PEs: 16 -> 57
			// srcs: (141, 37)(1205) 31 --> (1205) 31:PUGB2, pass, PENB
			9'd41 : rdata = 43'b1100011100101000000000000000000000100000000;
			// PEs: 56 -> 57
			// srcs: (147, 38)(1175) 198 --> (1175) 198:NI0, pass, PENB
			9'd42 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 56
			// srcs: (148, 39)(636) 140 --> (636) 140:PUGB0, pass, NI0
			9'd43 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 0 -> 57
			// srcs: (149, 40)(666) -22 --> (666) -22:PUGB0, pass, PENB
			9'd44 : rdata = 43'b1100011100001000000000000000000000100000000;
			// PEs: 56 -> 57
			// srcs: (155, 41)(636) 140 --> (636) 140:NI0, pass, PENB
			9'd45 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 16 -> 56
			// srcs: (156, 42)(1061) 504 --> (1061) 504:PUGB2, pass, NI0
			9'd46 : rdata = 43'b1100011100101000000001000000000000000000000;
			// PEs: 16 -> 57
			// srcs: (157, 43)(1091) 126 --> (1091) 126:PUGB2, pass, PENB
			9'd47 : rdata = 43'b1100011100101000000000000000000000100000000;
			// PEs: 57 -> 32
			// srcs: (162, 78)(1452) 118 --> (1452) 118:PEGB1, pass, PUGB4
			9'd48 : rdata = 43'b1100011100010000000000000000000000000001100;
			// PEs: 56 -> 57
			// srcs: (163, 44)(1061) 504 --> (1061) 504:NI0, pass, PENB
			9'd49 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 16 -> 56
			// srcs: (164, 45)(1121) 966 --> (1121) 966:PUGB2, pass, NI0
			9'd50 : rdata = 43'b1100011100101000000001000000000000000000000;
			// PEs: 16 -> 57
			// srcs: (165, 46)(1151) 533 --> (1151) 533:PUGB2, pass, PENB
			9'd51 : rdata = 43'b1100011100101000000000000000000000100000000;
			// PEs: 56 -> 57
			// srcs: (171, 47)(1121) 966 --> (1121) 966:NI0, pass, PENB
			9'd52 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 16 -> 56
			// srcs: (172, 48)(1181) 378 --> (1181) 378:PUGB2, pass, NI0
			9'd53 : rdata = 43'b1100011100101000000001000000000000000000000;
			// PEs: 16 -> 57
			// srcs: (173, 49)(1211) 1333 --> (1211) 1333:PUGB2, pass, PENB
			9'd54 : rdata = 43'b1100011100101000000000000000000000100000000;
			// PEs: 56 -> 57
			// srcs: (179, 50)(1181) 378 --> (1181) 378:NI0, pass, PENB
			9'd55 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 56
			// srcs: (180, 51)(642) 238 --> (642) 238:PUGB0, pass, NI0
			9'd56 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 0 -> 57
			// srcs: (181, 52)(672) 506 --> (672) 506:PUGB0, pass, PENB
			9'd57 : rdata = 43'b1100011100001000000000000000000000100000000;
			// PEs: 56 -> 57
			// srcs: (187, 53)(642) 238 --> (642) 238:NI0, pass, PENB
			9'd58 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 56
			// srcs: (188, 54)(702) 864 --> (702) 864:PUGB0, pass, NI0
			9'd59 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 0 -> 57
			// srcs: (189, 55)(732) 1748 --> (732) 1748:PUGB0, pass, PENB
			9'd60 : rdata = 43'b1100011100001000000000000000000000100000000;
			// PEs: 56 -> 57
			// srcs: (195, 56)(702) 864 --> (702) 864:NI0, pass, PENB
			9'd61 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 56
			// srcs: (196, 57)(762) 1056 --> (762) 1056:PUGB0, pass, NI0
			9'd62 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 0 -> 57
			// srcs: (197, 58)(792) 114 --> (792) 114:PUGB0, pass, PENB
			9'd63 : rdata = 43'b1100011100001000000000000000000000100000000;
			// PEs: 56 -> 57
			// srcs: (203, 59)(762) 1056 --> (762) 1056:NI0, pass, PENB
			9'd64 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 56
			// srcs: (204, 60)(822) 1364 --> (822) 1364:PUGB0, pass, NI0
			9'd65 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 8 -> 57
			// srcs: (205, 61)(852) 256 --> (852) 256:PUGB1, pass, PENB
			9'd66 : rdata = 43'b1100011100011000000000000000000000100000000;
			// PEs: 56 -> 57
			// srcs: (211, 62)(822) 1364 --> (822) 1364:NI0, pass, PENB
			9'd67 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 8 -> 56
			// srcs: (212, 63)(882) 576 --> (882) 576:PUGB1, pass, NI0
			9'd68 : rdata = 43'b1100011100011000000001000000000000000000000;
			// PEs: 8 -> 57
			// srcs: (213, 64)(912) -20 --> (912) -20:PUGB1, pass, PENB
			9'd69 : rdata = 43'b1100011100011000000000000000000000100000000;
			// PEs: 56 -> 57
			// srcs: (219, 65)(882) 576 --> (882) 576:NI0, pass, PENB
			9'd70 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 24 -> 56
			// srcs: (220, 66)(1266) 411 --> (1266) 411:PUGB3, pass, NI0
			9'd71 : rdata = 43'b1100011100111000000001000000000000000000000;
			// PEs: 40 -> 57
			// srcs: (221, 67)(1267) 281 --> (1267) 281:PUGB5, pass, PENB
			9'd72 : rdata = 43'b1100011101011000000000000000000000100000000;
			// PEs: 57 -> 16
			// srcs: (224, 92)(1581) 6146 --> (1581) 6146:PEGB1, pass, PUGB2
			9'd73 : rdata = 43'b1100011100010000000000000000000000000001010;
			// PEs: 57 -> 0
			// srcs: (226, 80)(1570) 556 --> (1570) 556:PEGB1, pass, PUNB
			9'd74 : rdata = 43'b1100011100010000000000000000000001000000000;
			// PEs: 56 -> 57
			// srcs: (227, 68)(1266) 411 --> (1266) 411:NI0, pass, PENB
			9'd75 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 40 -> 56
			// srcs: (228, 69)(1268) 34 --> (1268) 34:PUGB5, pass, NI0
			9'd76 : rdata = 43'b1100011101011000000001000000000000000000000;
			// PEs: 24 -> 57
			// srcs: (229, 70)(1269) 1425 --> (1269) 1425:PUGB3, pass, PENB
			9'd77 : rdata = 43'b1100011100111000000000000000000000100000000;
			// PEs: 56 -> 57
			// srcs: (235, 71)(1268) 34 --> (1268) 34:NI0, pass, PENB
			9'd78 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 48 -> 56
			// srcs: (236, 72)(1306) 458 --> (1306) 458:PUNB, pass, NI0
			9'd79 : rdata = 43'b1100011011111000000001000000000000000000000;
			// PEs: 57 -> 0
			// srcs: (237, 86)(1331) 2705 --> (1331) 2705:PEGB1, pass, PUNB
			9'd80 : rdata = 43'b1100011100010000000000000000000001000000000;
			// PEs: 57 -> 32
			// srcs: (245, 93)(1278) 2151 --> (1278) 2151:PEGB1, pass, PUGB4
			9'd81 : rdata = 43'b1100011100010000000000000000000000000001100;
			// PEs: 16 -> 57
			// srcs: (326, 73)(1307) 1302 --> (1307) 1302:PUGB2, pass, PENB
			9'd82 : rdata = 43'b1100011100101000000000000000000000100000000;
			// PEs: 56 -> 57
			// srcs: (332, 74)(1306) 458 --> (1306) 458:NI0, pass, PENB
			9'd83 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 48 -> 57
			// srcs: (333, 76)(1435) 280 --> (1435) 280:PUNB, pass, PENB
			9'd84 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 48 -> 57
			// srcs: (334, 79)(1553) -14 --> (1553) -14:PUNB, pass, PENB
			9'd85 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 0 -> 56
			// srcs: (335, 81)(1572) 636 --> (1572) 636:PUGB0, pass, NI0
			9'd86 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 24 -> 57
			// srcs: (454, 82)(1573) 1284 --> (1573) 1284:PUGB3, pass, PENB
			9'd87 : rdata = 43'b1100011100111000000000000000000000100000000;
			// PEs: 56 -> 57
			// srcs: (461, 83)(1572) 636 --> (1572) 636:NI0, pass, PENB
			9'd88 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 48 -> 57
			// srcs: (462, 84)(1443) 1383 --> (1443) 1383:PUNB, pass, PENB
			9'd89 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 48 -> 57
			// srcs: (463, 85)(1312) 811 --> (1312) 811:PUNB, pass, PENB
			9'd90 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 48 -> 57
			// srcs: (464, 88)(1559) 3128 --> (1559) 3128:PUNB, pass, PENB
			9'd91 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 48 -> 57
			// srcs: (465, 91)(1562) 2741 --> (1562) 2741:PUNB, pass, PENB
			9'd92 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 57 -> 0
			// srcs: (468, 89)(1579) 1920 --> (1579) 1920:PEGB1, pass, PUNB
			9'd93 : rdata = 43'b1100011100010000000000000000000001000000000;
			// PEs: 57 -> 32
			// srcs: (470, 94)(1316) 2571 --> (1316) 2571:PEGB1, pass, PUGB4
			9'd94 : rdata = 43'b1100011100010000000000000000000000000001100;
			// PEs: 48 -> 57
			// srcs: (563, 95)(1449) 4386 --> (1449) 4386:PUNB, pass, PENB
			9'd95 : rdata = 43'b1100011011111000000000000000000000100000000;
			// PEs: 16 -> 56
			// srcs: (564, 96)(1639) 3149 --> (1639) 3149:PUGB2, pass, NI0
			9'd96 : rdata = 43'b1100011100101000000001000000000000000000000;
			// PEs: 32 -> 57
			// srcs: (956, 97)(1640) 3270 --> (1640) 3270:PUGB4, pass, PENB
			9'd97 : rdata = 43'b1100011101001000000000000000000000100000000;
			// PEs: 56 -> 57
			// srcs: (963, 98)(1639) 3149 --> (1639) 3149:NI0, pass, PENB
			9'd98 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 16 -> 56
			// srcs: (1046, 99)(1658) 5192 --> (1658) 5192:PUGB2, pass, NI0
			9'd99 : rdata = 43'b1100011100101000000001000000000000000000000;
			// PEs: 32 -> 57
			// srcs: (1047, 100)(1659) 5518 --> (1659) 5518:PUGB4, pass, PENB
			9'd100 : rdata = 43'b1100011101001000000000000000000000100000000;
			// PEs: 56 -> 57
			// srcs: (1053, 101)(1658) 5192 --> (1658) 5192:NI0, pass, PENB
			9'd101 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 16 -> 56
			// srcs: (1717, 102)(1677) 3421 --> (1677) 3421:PUGB2, pass, NI0
			9'd102 : rdata = 43'b1100011100101000000001000000000000000000000;
			// PEs: 32 -> 57
			// srcs: (1718, 103)(1678) 5382 --> (1678) 5382:PUGB4, pass, PENB
			9'd103 : rdata = 43'b1100011101001000000000000000000000100000000;
			// PEs: 56 -> 57
			// srcs: (1724, 104)(1677) 3421 --> (1677) 3421:NI0, pass, PENB
			9'd104 : rdata = 43'b1100010100000000000000000000000000100000000;
			// PEs: 0 -> 56
			// srcs: (1725, 105)(1753) 2905 --> (1753) 2905:PUGB0, pass, NI0
			9'd105 : rdata = 43'b1100011100001000000001000000000000000000000;
			// PEs: 32 -> 57
			// srcs: (1726, 106)(1754) 6068 --> (1754) 6068:PUGB4, pass, PENB
			9'd106 : rdata = 43'b1100011101001000000000000000000000100000000;
			// PEs: 56 -> 57
			// srcs: (1732, 107)(1753) 2905 --> (1753) 2905:NI0, pass, PENB
			9'd107 : rdata = 43'b1100010100000000000000000000000000100000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 57) begin
	always @(*) begin
		case(address)
			// PEs: 56 -> 
			// srcs: (47, 0)(659) 22 --> (659) 22:PENB, pass, 
			9'd0 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 56, 57 -> 57
			// srcs: (53, 1)(629) 630, (659) 22 --> (1319) 652:PENB, ALU, +, NI0
			9'd1 : rdata = 43'b0000111011110001111111000000000000000000000;
			// PEs: 56 -> 
			// srcs: (55, 2)(719) 1104 --> (719) 1104:PENB, pass, 
			9'd2 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 56, 57 -> 57
			// srcs: (61, 3)(689) 600, (719) 1104 --> (1320) 1704:PENB, ALU, +, NI1
			9'd3 : rdata = 43'b0000111011110001111111000010000000000000000;
			// PEs: 56 -> 57
			// srcs: (63, 4)(779) 95 --> (779) 95:PENB, pass, NI2
			9'd4 : rdata = 43'b1100011011110000000001000100000000000000000;
			// PEs: 57 -> 57
			// srcs: (64, 81)(1319) 652 --> (1319) 652:NI0, pass, NI0
			9'd5 : rdata = 43'b1100010100000000000001000000000000000000000;
			// PEs: 57, 57 -> 57
			// srcs: (64, 50)(1319) 652, (1320) 1704 --> (1329) 2356:ALU, NI1, +, NI3
			9'd6 : rdata = 43'b0000100111111101000011000110000000000000000;
			// PEs: 56, 57 -> 57
			// srcs: (69, 5)(749) 360, (779) 95 --> (1321) 455:PENB, NI2, +, NI0
			9'd7 : rdata = 43'b0000111011110101000101000000000000000000000;
			// PEs: 56 -> 
			// srcs: (71, 6)(839) 736 --> (839) 736:PENB, pass, 
			9'd8 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 56, 57 -> 57
			// srcs: (77, 7)(809) 310, (839) 736 --> (1322) 1046:PENB, ALU, +, NI1
			9'd9 : rdata = 43'b0000111011110001111111000010000000000000000;
			// PEs: 56 -> 57
			// srcs: (79, 8)(899) -4 --> (899) -4:PENB, pass, NI2
			9'd10 : rdata = 43'b1100011011110000000001000100000000000000000;
			// PEs: 57 -> 57
			// srcs: (80, 82)(1321) 455 --> (1321) 455:NI0, pass, NI0
			9'd11 : rdata = 43'b1100010100000000000001000000000000000000000;
			// PEs: 57, 57 -> 
			// srcs: (80, 51)(1321) 455, (1322) 1046 --> (1330) 1501:ALU, NI1, +, 
			9'd12 : rdata = 43'b0000100111111101000010000000000000000000000;
			// PEs: 57, 57 -> 56
			// srcs: (83, 62)(1329) 2356, (1330) 1501 --> (1334) 3857:NI3, ALU, +, PEGB0
			9'd13 : rdata = 43'b0000110100011001111110000000000000010000000;
			// PEs: 56, 57 -> 57
			// srcs: (85, 9)(869) 704, (899) -4 --> (1323) 700:PENB, NI2, +, NI0
			9'd14 : rdata = 43'b0000111011110101000101000000000000000000000;
			// PEs: 56 -> 
			// srcs: (87, 10)(959) 990 --> (959) 990:PENB, pass, 
			9'd15 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 56, 57 -> 57
			// srcs: (93, 11)(929) 1015, (959) 990 --> (1324) 2005:PENB, ALU, +, NI1
			9'd16 : rdata = 43'b0000111011110001111111000010000000000000000;
			// PEs: 56 -> 57
			// srcs: (95, 12)(1019) 506 --> (1019) 506:PENB, pass, NI2
			9'd17 : rdata = 43'b1100011011110000000001000100000000000000000;
			// PEs: 57 -> 57
			// srcs: (96, 83)(1323) 700 --> (1323) 700:NI0, pass, NI0
			9'd18 : rdata = 43'b1100010100000000000001000000000000000000000;
			// PEs: 57, 57 -> 57
			// srcs: (96, 52)(1323) 700, (1324) 2005 --> (1331) 2705:ALU, NI1, +, NI3
			9'd19 : rdata = 43'b0000100111111101000011000110000000000000000;
			// PEs: 56, 57 -> 56
			// srcs: (101, 13)(989) 90, (1019) 506 --> (1325) 596:PENB, NI2, +, PEGB0
			9'd20 : rdata = 43'b0000111011110101000100000000000000010000000;
			// PEs: 56 -> 
			// srcs: (103, 14)(845) 672 --> (845) 672:PENB, pass, 
			9'd21 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 56, 57 -> 57
			// srcs: (109, 15)(815) 1054, (845) 672 --> (1436) 1726:PENB, ALU, +, NI0
			9'd22 : rdata = 43'b0000111011110001111111000000000000000000000;
			// PEs: 56 -> 
			// srcs: (111, 16)(905) -35 --> (905) -35:PENB, pass, 
			9'd23 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 56, 57 -> 57
			// srcs: (117, 17)(875) 1536, (905) -35 --> (1437) 1501:PENB, ALU, +, NI1
			9'd24 : rdata = 43'b0000111011110001111111000010000000000000000;
			// PEs: 56 -> 
			// srcs: (119, 18)(965) -99 --> (965) -99:PENB, pass, 
			9'd25 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 56, 57 -> 57
			// srcs: (125, 19)(935) 1044, (965) -99 --> (1438) 945:PENB, ALU, +, NI2
			9'd26 : rdata = 43'b0000111011110001111111000100000000000000000;
			// PEs: 56 -> 57
			// srcs: (127, 20)(1025) 308 --> (1025) 308:PENB, pass, NI4
			9'd27 : rdata = 43'b1100011011110000000001001000000000000000000;
			// PEs: 57 -> 57
			// srcs: (128, 84)(1437) 1501 --> (1437) 1501:NI1, pass, NI1
			9'd28 : rdata = 43'b1100010100001000000001000010000000000000000;
			// PEs: 57, 57 -> 56
			// srcs: (128, 54)(1437) 1501, (1438) 945 --> (1445) 2446:ALU, NI2, +, PEGB0
			9'd29 : rdata = 43'b0000100111111101000100000000000000010000000;
			// PEs: 56, 57 -> 56
			// srcs: (133, 21)(995) 60, (1025) 308 --> (1439) 368:PENB, NI4, +, PEGB0
			9'd30 : rdata = 43'b0000111011110101001000000000000000010000000;
			// PEs: 56 -> 
			// srcs: (135, 22)(1145) 312 --> (1145) 312:PENB, pass, 
			9'd31 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 56, 57 -> 57
			// srcs: (141, 23)(1115) 69, (1145) 312 --> (1441) 381:PENB, ALU, +, NI1
			9'd32 : rdata = 43'b0000111011110001111111000010000000000000000;
			// PEs: 56 -> 
			// srcs: (143, 24)(1205) 31 --> (1205) 31:PENB, pass, 
			9'd33 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 56, 57 -> 57
			// srcs: (149, 25)(1175) 198, (1205) 31 --> (1442) 229:PENB, ALU, +, NI2
			9'd34 : rdata = 43'b0000111011110001111111000100000000000000000;
			// PEs: 56 -> 57
			// srcs: (151, 26)(666) -22 --> (666) -22:PENB, pass, NI4
			9'd35 : rdata = 43'b1100011011110000000001001000000000000000000;
			// PEs: 57 -> 57
			// srcs: (152, 85)(1441) 381 --> (1441) 381:NI1, pass, NI1
			9'd36 : rdata = 43'b1100010100001000000001000010000000000000000;
			// PEs: 57, 57 -> 57
			// srcs: (152, 60)(1441) 381, (1442) 229 --> (1447) 610:ALU, NI2, +, NI5
			9'd37 : rdata = 43'b0000100111111101000101001010000000000000000;
			// PEs: 56, 57 -> 56
			// srcs: (157, 27)(636) 140, (666) -22 --> (1452) 118:PENB, NI4, +, PEGB0
			9'd38 : rdata = 43'b0000111011110101001000000000000000010000000;
			// PEs: 56 -> 
			// srcs: (159, 28)(1091) 126 --> (1091) 126:PENB, pass, 
			9'd39 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 56, 57 -> 57
			// srcs: (165, 29)(1061) 504, (1091) 126 --> (1554) 630:PENB, ALU, +, NI1
			9'd40 : rdata = 43'b0000111011110001111111000010000000000000000;
			// PEs: 56 -> 
			// srcs: (167, 30)(1151) 533 --> (1151) 533:PENB, pass, 
			9'd41 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 56, 57 -> 57
			// srcs: (173, 31)(1121) 966, (1151) 533 --> (1555) 1499:PENB, ALU, +, NI2
			9'd42 : rdata = 43'b0000111011110001111111000100000000000000000;
			// PEs: 56 -> 
			// srcs: (175, 32)(1211) 1333 --> (1211) 1333:PENB, pass, 
			9'd43 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 56, 57 -> 57
			// srcs: (181, 33)(1181) 378, (1211) 1333 --> (1556) 1711:PENB, ALU, +, NI4
			9'd44 : rdata = 43'b0000111011110001111111001000000000000000000;
			// PEs: 56 -> 57
			// srcs: (183, 34)(672) 506 --> (672) 506:PENB, pass, NI6
			9'd45 : rdata = 43'b1100011011110000000001001100000000000000000;
			// PEs: 57 -> 57
			// srcs: (184, 86)(1555) 1499 --> (1555) 1499:NI2, pass, NI2
			9'd46 : rdata = 43'b1100010100010000000001000100000000000000000;
			// PEs: 57, 57 -> 57
			// srcs: (184, 61)(1555) 1499, (1556) 1711 --> (1561) 3210:ALU, NI4, +, NI7
			9'd47 : rdata = 43'b0000100111111101001001001110000000000000000;
			// PEs: 56, 57 -> 57
			// srcs: (189, 35)(642) 238, (672) 506 --> (1566) 744:PENB, NI6, +, NI2
			9'd48 : rdata = 43'b0000111011110101001101000100000000000000000;
			// PEs: 56 -> 
			// srcs: (191, 36)(732) 1748 --> (732) 1748:PENB, pass, 
			9'd49 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 56, 57 -> 57
			// srcs: (197, 37)(702) 864, (732) 1748 --> (1567) 2612:PENB, ALU, +, NI4
			9'd50 : rdata = 43'b0000111011110001111111001000000000000000000;
			// PEs: 56 -> 57
			// srcs: (199, 38)(792) 114 --> (792) 114:PENB, pass, NI6
			9'd51 : rdata = 43'b1100011011110000000001001100000000000000000;
			// PEs: 57 -> 57
			// srcs: (200, 87)(1566) 744 --> (1566) 744:NI2, pass, NI2
			9'd52 : rdata = 43'b1100010100010000000001000100000000000000000;
			// PEs: 57, 57 -> 57
			// srcs: (200, 56)(1566) 744, (1567) 2612 --> (1576) 3356:ALU, NI4, +, NI8
			9'd53 : rdata = 43'b0000100111111101001001010000000000000000000;
			// PEs: 56, 57 -> 57
			// srcs: (205, 39)(762) 1056, (792) 114 --> (1568) 1170:PENB, NI6, +, NI2
			9'd54 : rdata = 43'b0000111011110101001101000100000000000000000;
			// PEs: 56 -> 
			// srcs: (207, 40)(852) 256 --> (852) 256:PENB, pass, 
			9'd55 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 56, 57 -> 57
			// srcs: (213, 41)(822) 1364, (852) 256 --> (1569) 1620:PENB, ALU, +, NI4
			9'd56 : rdata = 43'b0000111011110001111111001000000000000000000;
			// PEs: 56 -> 57
			// srcs: (215, 42)(912) -20 --> (912) -20:PENB, pass, NI6
			9'd57 : rdata = 43'b1100011011110000000001001100000000000000000;
			// PEs: 57 -> 57
			// srcs: (216, 88)(1568) 1170 --> (1568) 1170:NI2, pass, NI2
			9'd58 : rdata = 43'b1100010100010000000001000100000000000000000;
			// PEs: 57, 57 -> 
			// srcs: (216, 57)(1568) 1170, (1569) 1620 --> (1577) 2790:ALU, NI4, +, 
			9'd59 : rdata = 43'b0000100111111101001000000000000000000000000;
			// PEs: 57, 57 -> 56
			// srcs: (219, 64)(1576) 3356, (1577) 2790 --> (1581) 6146:NI8, ALU, +, PEGB0
			9'd60 : rdata = 43'b0000110101000001111110000000000000010000000;
			// PEs: 56, 57 -> 56
			// srcs: (221, 43)(882) 576, (912) -20 --> (1570) 556:PENB, NI6, +, PEGB0
			9'd61 : rdata = 43'b0000111011110101001100000000000000010000000;
			// PEs: 56 -> 
			// srcs: (223, 44)(1267) 281 --> (1267) 281:PENB, pass, 
			9'd62 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 56, 57 -> 57
			// srcs: (229, 45)(1266) 411, (1267) 281 --> (1274) 692:PENB, ALU, +, NI2
			9'd63 : rdata = 43'b0000111011110001111111000100000000000000000;
			// PEs: 56 -> 57
			// srcs: (231, 46)(1269) 1425 --> (1269) 1425:PENB, pass, NI4
			9'd64 : rdata = 43'b1100011011110000000001001000000000000000000;
			// PEs: 57 -> 56
			// srcs: (232, 67)(1331) 2705 --> (1331) 2705:NI3, pass, PEGB0
			9'd65 : rdata = 43'b1100010100011000000000000000000000010000000;
			// PEs: 56, 57 -> 
			// srcs: (237, 47)(1268) 34, (1269) 1425 --> (1275) 1459:PENB, NI4, +, 
			9'd66 : rdata = 43'b0000111011110101001000000000000000000000000;
			// PEs: 57, 57 -> 56
			// srcs: (240, 65)(1274) 692, (1275) 1459 --> (1278) 2151:NI2, ALU, +, PEGB0
			9'd67 : rdata = 43'b0000110100010001111110000000000000010000000;
			// PEs: 56 -> 
			// srcs: (328, 48)(1307) 1302 --> (1307) 1302:PENB, pass, 
			9'd68 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 56, 57 -> 57
			// srcs: (334, 49)(1306) 458, (1307) 1302 --> (1313) 1760:PENB, ALU, +, NI2
			9'd69 : rdata = 43'b0000111011110001111111000100000000000000000;
			// PEs: 56, 57 -> 57
			// srcs: (335, 53)(1435) 280, (1436) 1726 --> (1444) 2006:PENB, NI0, +, NI3
			9'd70 : rdata = 43'b0000111011110101000001000110000000000000000;
			// PEs: 56, 57 -> 57
			// srcs: (336, 55)(1553) -14, (1554) 630 --> (1560) 616:PENB, NI1, +, NI0
			9'd71 : rdata = 43'b0000111011110101000011000000000000000000000;
			// PEs: 56 -> 
			// srcs: (456, 58)(1573) 1284 --> (1573) 1284:PENB, pass, 
			9'd72 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 56, 57 -> 56
			// srcs: (463, 59)(1572) 636, (1573) 1284 --> (1579) 1920:PENB, ALU, +, PEGB0
			9'd73 : rdata = 43'b0000111011110001111110000000000000010000000;
			// PEs: 56, 57 -> 57
			// srcs: (464, 63)(1443) 1383, (1444) 2006 --> (1448) 3389:PENB, NI3, +, NI1
			9'd74 : rdata = 43'b0000111011110101000111000010000000000000000;
			// PEs: 56, 57 -> 56
			// srcs: (465, 66)(1312) 811, (1313) 1760 --> (1316) 2571:PENB, NI2, +, PEGB0
			9'd75 : rdata = 43'b0000111011110101000100000000000000010000000;
			// PEs: 56, 57 -> 57
			// srcs: (466, 68)(1559) 3128, (1560) 616 --> (1563) 3744:PENB, NI0, +, NI2
			9'd76 : rdata = 43'b0000111011110101000001000100000000000000000;
			// PEs: 57 -> 57
			// srcs: (467, 89)(1447) 610 --> (1447) 610:NI5, pass, NI5
			9'd77 : rdata = 43'b1100010100101000000001001010000000000000000;
			// PEs: 57, 57 -> 57
			// srcs: (467, 69)(1447) 610, (1448) 3389 --> (1450) 3999:ALU, NI1, +, NI0
			9'd78 : rdata = 43'b0000100111111101000011000000000000000000000;
			// PEs: 57, 56 -> 
			// srcs: (468, 70)(1561) 3210, (1562) 2741 --> (1564) 5951:NI7, PENB, +, 
			9'd79 : rdata = 43'b0000110100111110111100000000000000000000000;
			// PEs: 57, 57 -> 57
			// srcs: (471, 72)(1563) 3744, (1564) 5951 --> (1565) 9695:NI2, ALU, +, NW1
			9'd80 : rdata = 43'b0000110100010001111110000001000010000000000;
			// PEs: 56, 57 -> 57
			// srcs: (566, 71)(1449) 4386, (1450) 3999 --> (1451) 8385:PENB, NI0, +, NW0
			9'd81 : rdata = 43'b0000111011110101000000000001000000000000000;
			// PEs: 56 -> 
			// srcs: (958, 73)(1640) 3270 --> (1640) 3270:PENB, pass, 
			9'd82 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 56, 57 -> 57
			// srcs: (965, 74)(1639) 3149, (1640) 3270 --> (1641) 6419:PENB, ALU, +, NW2
			9'd83 : rdata = 43'b0000111011110001111110000001000100000000000;
			// PEs: 56 -> 
			// srcs: (1049, 75)(1659) 5518 --> (1659) 5518:PENB, pass, 
			9'd84 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 56, 57 -> 57
			// srcs: (1055, 76)(1658) 5192, (1659) 5518 --> (1660) 10710:PENB, ALU, +, NW3
			9'd85 : rdata = 43'b0000111011110001111110000001000110000000000;
			// PEs: 56 -> 
			// srcs: (1720, 77)(1678) 5382 --> (1678) 5382:PENB, pass, 
			9'd86 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 56, 57 -> 57
			// srcs: (1726, 78)(1677) 3421, (1678) 5382 --> (1679) 8803:PENB, ALU, +, NW4
			9'd87 : rdata = 43'b0000111011110001111110000001001000000000000;
			// PEs: 56 -> 
			// srcs: (1728, 79)(1754) 6068 --> (1754) 6068:PENB, pass, 
			9'd88 : rdata = 43'b1100011011110000000000000000000000000000000;
			// PEs: 56, 57 -> 57
			// srcs: (1734, 80)(1753) 2905, (1754) 6068 --> (1755) 8973:PENB, ALU, +, NW5
			9'd89 : rdata = 43'b0000111011110001111110000001001010000000000;
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 58) begin
	always @(*) begin
		case(address)
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 59) begin
	always @(*) begin
		case(address)
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 60) begin
	always @(*) begin
		case(address)
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 61) begin
	always @(*) begin
		case(address)
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 62) begin
	always @(*) begin
		case(address)
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 63) begin
	always @(*) begin
		case(address)
			default : rdata = 43'b0000000000000000000000000000000000000000000;
		endcase
	end
end

endgenerate
/*****************************************************************************/
endmodule
