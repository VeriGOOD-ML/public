//-----------------------------------------------------------
//Simple Log2 calculation function
//-----------------------------------------------------------
`define C_LOG_2(n) (\
(n) < (1<<0) ? 0 : (n) <= (1<<1) ? 1 :\
(n) <= (1<<2) ? 2 : (n) <= (1<<3) ? 3 :\
(n) <= (1<<4) ? 4 : (n) <= (1<<5) ? 5 :\
(n) <= (1<<6) ? 6 : (n) <= (1<<7) ? 7 :\
(n) <= (1<<8) ? 8 : (n) <= (1<<9) ? 9 :\
(n) <= (1<<10) ? 10 : (n) <= (1<<11) ? 11 :\
(n) <= (1<<12) ? 12 : (n) <= (1<<13) ? 13 :\
(n) <= (1<<14) ? 14 : (n) <= (1<<15) ? 15 :\
(n) <= (1<<16) ? 16 : (n) <= (1<<17) ? 17 :\
(n) <= (1<<18) ? 18 : (n) <= (1<<19) ? 19 :\
(n) <= (1<<20) ? 20 : (n) <= (1<<21) ? 21 :\
(n) <= (1<<22) ? 22 : (n) <= (1<<23) ? 23 :\
(n) <= (1<<24) ? 24 : (n) <= (1<<25) ? 25 :\
(n) <= (1<<26) ? 26 : (n) <= (1<<27) ? 27 :\
(n) <= (1<<28) ? 28 : (n) <= (1<<29) ? 29 :\
(n) <= (1<<30) ? 30 : (n) <= (1<<31) ? 31 : 32)
//-----------------------------------------------------------
//`define WEIGHT_COUNT_MACRO(lanes,pe) (\
//(lanes%8) == 0 ? 0 : (pe == 4)? 56 : 14)

//`define WEIGHT_COUNT_MACRO(lanes,pe) (\
//(lanes == 0 && pe == 0) ? 16'h0 : \
//(lanes == 0 && pe == 1) ? 16'h0 : \
//(lanes == 0 && pe == 2) ? 16'h0 : \
//(lanes == 0 && pe == 3) ? 16'h0 : \
//(lanes == 0 && pe == 4) ? 16'h0 : \
//(lanes == 1 && pe == 0) ? 16'h2 : \
//(lanes == 1 && pe == 1) ? 16'h2 : \
//(lanes == 1 && pe == 2) ? 16'h2 : \
//(lanes == 1 && pe == 3) ? 16'h2 : \
//(lanes == 1 && pe == 4) ? 16'h8 : \
//(lanes == 2 && pe == 0) ? 16'h2 : \
//(lanes == 2 && pe == 1) ? 16'h2 : \
//(lanes == 2 && pe == 2) ? 16'h2 : \
//(lanes == 2 && pe == 3) ? 16'h2 : \
//(lanes == 2 && pe == 4) ? 16'h8 : \
//(lanes == 3 && pe == 0) ? 16'h2 : \
//(lanes == 3 && pe == 1) ? 16'h2 : \
//(lanes == 3 && pe == 2) ? 16'h2 : \
//(lanes == 3 && pe == 3) ? 16'h1 : \
//(lanes == 3 && pe == 4) ? 16'h7 : \
//(lanes == 4 && pe == 0) ? 16'h2 : \
//(lanes == 4 && pe == 1) ? 16'h2 : \
//(lanes == 4 && pe == 2) ? 16'h2 : \
//(lanes == 4 && pe == 3) ? 16'h1 : \
//(lanes == 4 && pe == 4) ? 16'h7 : \
//(lanes == 5 && pe == 0) ? 16'h2 : \
//(lanes == 5 && pe == 1) ? 16'h2 : \
//(lanes == 5 && pe == 2) ? 16'h2 : \
//(lanes == 5 && pe == 3) ? 16'h1 : \
//(lanes == 5 && pe == 4) ? 16'h7 : \
//(lanes == 6 && pe == 0) ? 16'h2 : \
//(lanes == 6 && pe == 1) ? 16'h2 : \
//(lanes == 6 && pe == 2) ? 16'h2 : \
//(lanes == 6 && pe == 3) ? 16'h1 : \
//(lanes == 6 && pe == 4) ? 16'h7 : \
//(lanes == 7 && pe == 0) ? 16'h2 : \
//(lanes == 7 && pe == 1) ? 16'h2 : \
//(lanes == 7 && pe == 2) ? 16'h2 : \
//(lanes == 7 && pe == 3) ? 16'h1 : \
//(lanes == 7 && pe == 4) ? 16'h7 : \
//(lanes == 8 && pe == 0) ? 16'h0 : \
//(lanes == 8 && pe == 1) ? 16'h0 : \
//(lanes == 8 && pe == 2) ? 16'h0 : \
//(lanes == 8 && pe == 3) ? 16'h0 : \
//(lanes == 8 && pe == 4) ? 16'h0 : \
//(lanes == 9 && pe == 0) ? 16'h2 : \
//(lanes == 9 && pe == 1) ? 16'h2 : \
//(lanes == 9 && pe == 2) ? 16'h2 : \
//(lanes == 9 && pe == 3) ? 16'h1 : \
//(lanes == 9 && pe == 4) ? 16'h7 : \
//(lanes == 10 && pe == 0) ? 16'h2 : \
//(lanes == 10 && pe == 1) ? 16'h2 : \
//(lanes == 10 && pe == 2) ? 16'h2 : \
//(lanes == 10 && pe == 3) ? 16'h1 : \
//(lanes == 10 && pe == 4) ? 16'h7 : \
//(lanes == 11 && pe == 0) ? 16'h2 : \
//(lanes == 11 && pe == 1) ? 16'h2 : \
//(lanes == 11 && pe == 2) ? 16'h2 : \
//(lanes == 11 && pe == 3) ? 16'h1 : \
//(lanes == 11 && pe == 4) ? 16'h7 : \
//(lanes == 12 && pe == 0) ? 16'h2 : \
//(lanes == 12 && pe == 1) ? 16'h2 : \
//(lanes == 12 && pe == 2) ? 16'h2 : \
//(lanes == 12 && pe == 3) ? 16'h1 : \
//(lanes == 12 && pe == 4) ? 16'h7 : \
//(lanes == 13 && pe == 0) ? 16'h2 : \
//(lanes == 13 && pe == 1) ? 16'h2 : \
//(lanes == 13 && pe == 2) ? 16'h2 : \
//(lanes == 13 && pe == 3) ? 16'h1 : \
//(lanes == 13 && pe == 4) ? 16'h7 : \
//(lanes == 14 && pe == 0) ? 16'h2 : \
//(lanes == 14 && pe == 1) ? 16'h2 : \
//(lanes == 14 && pe == 2) ? 16'h2 : \
//(lanes == 14 && pe == 3) ? 16'h1 : \
//(lanes == 14 && pe == 4) ? 16'h7 : \
//(lanes == 15 && pe == 0) ? 16'h2 : \
//(lanes == 15 && pe == 1) ? 16'h2 : \
//(lanes == 15 && pe == 2) ? 16'h2 : \
//(lanes == 15 && pe == 3) ? 16'h1 : \
//16'h7)