`timescale 1ns/1ps

module ROM_ASIC #(
// Parameters
    parameter   DATA_WIDTH          = 16,
    parameter   ADDR_WIDTH          = 9,
    parameter   INIT                = "weight.txt",
    parameter   TYPE                = "block",
    parameter   ROM_DEPTH           = 1<<ADDR_WIDTH
) (
// Port Declarations
    input  wire                         CLK,
    input  wire                         RESET,
    input  wire  [ADDR_WIDTH-1:0]       ADDRESS,
    input  wire                         ENABLE,
    output reg   [DATA_WIDTH-1:0]       DATA_OUT,
    output reg                          DATA_OUT_VALID
);

// ******************************************************************
// Internal variables
// ******************************************************************

  localparam DEPTH = ROM_DEPTH;

  reg     [DATA_WIDTH-1:0]        rdata;
  wire     [ADDR_WIDTH-1:0]        address;

  assign address = ADDRESS;


  // `include "instructions.v"   // TODO
  always @(*) begin
	case(address)
/*****************************************************************************************/
//
// read [True, False, False, False]
// ['x2(0,)', 'x2(1,)', 'x2(3,)', 'x2(4,)', 'r2(60,)', 'r2(108,)', 'r2(123,)', 'r2(39,)', 'y2(108,)', 'y2(123,)', 'y2(34,)', 'r1(25,)', 'y1(117,)', 'r1(60,)', 'y1(60,)', 'r1(64,)']
// Data values: [1, 3, 3, 1, 1, 0, 1, 1, 1, 2, 5, 0, 4, 0, 1, 1]
// Dest PEs: [1, 2, 3, 4, 28, 29, 30, 31, 29, 30, 31, 34, 27, 34, 35, 42]
9'd0: rdata =    56'b00000000000000000000000000000000000000000000000000000001;
//
// shift amount: 15, Lanes IDs: [1, 2, 3, 4]
9'd1: rdata =    56'b00000000000000000000000000000000000100100100100001011111;
//
// read [True, False, False, False]
// ['x2(5,)', 'x2(6,)', 'x2(8,)', 'x2(9,)', 'r2(60,)', 'r2(108,)', 'r2(123,)', 'r2(39,)', 'y2(108,)', 'y2(123,)', 'y2(34,)', 'r1(25,)', 'y1(117,)', 'r1(60,)', 'y1(60,)', 'r1(64,)']
// Data values: [1, 5, 1, 2, 1, 0, 1, 1, 1, 2, 5, 0, 4, 0, 1, 1]
// Dest PEs: [5, 6, 7, 9, 28, 29, 30, 31, 29, 30, 31, 34, 27, 34, 35, 42]
9'd2: rdata =    56'b00000000000000000000000000000000000000000000000000000001;
//
// shift amount: 10, Lanes IDs: [9]
9'd3: rdata =    56'b00000000000000000000100000000000000000000000000001011010;
//
// shift amount: 11, Lanes IDs: [5, 6, 7]
9'd4: rdata =    56'b00000000000000000000000000100100100000000000000001011011;
//
// read [True, False, False, False]
// ['x1(0,)', 'x1(1,)', 'x1(3,)', 'x1(4,)', 'r2(60,)', 'r2(108,)', 'r2(123,)', 'r2(39,)', 'y2(108,)', 'y2(123,)', 'y2(34,)', 'r1(25,)', 'y1(117,)', 'r1(60,)', 'y1(60,)', 'r1(64,)']
// Data values: [3, 4, 2, 5, 1, 0, 1, 1, 1, 2, 5, 0, 4, 0, 1, 1]
// Dest PEs: [10, 11, 12, 13, 28, 29, 30, 31, 29, 30, 31, 34, 27, 34, 35, 42]
9'd5: rdata =    56'b00000000000000000000000000000000000000000000000000000001;
//
// shift amount: 6, Lanes IDs: [10, 11, 12, 13]
9'd6: rdata =    56'b00000000100100100100000000000000000000000000000001010110;
//
// read [True, False, False, False]
// ['x1(5,)', 'x1(6,)', 'x1(8,)', 'x1(9,)', 'r2(60,)', 'r2(108,)', 'r2(123,)', 'r2(39,)', 'y2(108,)', 'y2(123,)', 'y2(34,)', 'r1(25,)', 'y1(117,)', 'r1(60,)', 'y1(60,)', 'r1(64,)']
// Data values: [5, 5, 1, 1, 1, 0, 1, 1, 1, 2, 5, 0, 4, 0, 1, 1]
// Dest PEs: [14, 15, 17, 18, 28, 29, 30, 31, 29, 30, 31, 34, 27, 34, 35, 42]
9'd7: rdata =    56'b00000000000000000000000000000000000000000000000000000001;
//
// shift amount: 1, Lanes IDs: [1, 2]
9'd8: rdata =    56'b00000000000000000000000000000000000000001101100001010001;
//
// shift amount: 2, Lanes IDs: [14, 15]
9'd9: rdata =    56'b00100100000000000000000000000000000000000000000001010010;
//
// read [True, False, False, False]
// ['x2(2,)', 'x2(7,)', 'x1(2,)', 'x1(7,)', 'r2(60,)', 'r2(108,)', 'r2(123,)', 'r2(39,)', 'y2(108,)', 'y2(123,)', 'y2(34,)', 'r1(25,)', 'y1(117,)', 'r1(60,)', 'y1(60,)', 'r1(64,)']
// Data values: [3, 3, 5, 4, 1, 0, 1, 1, 1, 2, 5, 0, 4, 0, 1, 1]
// Dest PEs: [19, 20, 21, 22, 28, 29, 30, 31, 29, 30, 31, 34, 27, 34, 35, 42]
9'd10: rdata =   56'b00000000000000000000000000000000000000000000000000000001;
//
// shift amount: 13, Lanes IDs: [3, 4, 5, 6]
9'd11: rdata =   56'b00000000000000000000000000001101101101100000000001011101;
//
// read [True, False, False, False]
// ['r1(22,)', 'r1(54,)', 'r1(82,)', 'r1(112,)', 'r2(60,)', 'r2(108,)', 'r2(123,)', 'r2(39,)', 'y2(108,)', 'y2(123,)', 'y2(34,)', 'r1(25,)', 'y1(117,)', 'r1(60,)', 'y1(60,)', 'r1(64,)']
// Data values: [1, 1, 1, 0, 1, 0, 1, 1, 1, 2, 5, 0, 4, 0, 1, 1]
// Dest PEs: [23, 26, 27, 28, 28, 29, 30, 31, 29, 30, 31, 34, 27, 34, 35, 42]
9'd12: rdata =   56'b00000000000000000000000000000000000000000000000000000001;
//
// shift amount: 9, Lanes IDs: [7]
9'd13: rdata =   56'b00000000000000000000000001100000000000000000000001011001;
//
// shift amount: 7, Lanes IDs: [10, 11, 12]
9'd14: rdata =   56'b00000000001101101100000000000000000000000000000001010111;
//
// read [True, True, False, False]
// ['r2(2,)', 'r2(34,)', 'r1(34,)', 'r1(7,)', 'r2(60,)', 'r2(108,)', 'r2(123,)', 'r2(39,)', 'y2(108,)', 'y2(123,)', 'y2(34,)', 'r1(25,)', 'y1(117,)', 'r1(60,)', 'y1(60,)', 'r1(64,)']
// Data values: [1, 0, 1, 0, 1, 0, 1, 1, 1, 2, 5, 0, 4, 0, 1, 1]
// Dest PEs: [29, 30, 31, 34, 28, 29, 30, 31, 29, 30, 31, 34, 27, 34, 35, 42]
9'd15: rdata =   56'b00000000000000000000000000000000000000000000000000000011;
//
// shift amount: 1, Lanes IDs: [2]
9'd16: rdata =   56'b00000000000000000000000000000000000000010100000001010001;
//
// shift amount: 3, Lanes IDs: [13, 14, 15]
9'd17: rdata =   56'b01101101100000000000000000000000000000000000000001010011;
//
// shift amount: 8, Lanes IDs: [12, 13, 14, 15]
9'd18: rdata =   56'b01101101101100000000000000000000000000000000000001011000;
//
// read [True, False, False, False]
// ['r1(77,)', 'y1(77,)', 'r1(102,)', 'y1(102,)', 'r1(12,)', 'y1(7,)', 'r1(15,)', 'y1(15,)', 'y2(108,)', 'y2(123,)', 'y2(34,)', 'r1(25,)', 'y1(117,)', 'r1(60,)', 'y1(60,)', 'r1(64,)']
// Data values: [1, 5, 1, 0, 0, 4, 1, 0, 1, 2, 5, 0, 4, 0, 1, 1]
// Dest PEs: [35, 36, 37, 38, 34, 35, 42, 43, 29, 30, 31, 34, 27, 34, 35, 42]
9'd19: rdata =   56'b00000000000000000000000000000000000000000000000000000001;
//
// shift amount: 13, Lanes IDs: [3, 4, 5, 6]
9'd20: rdata =   56'b00000000000000000000000000010110110110100000000001011101;
//
// read [True, True, False, False]
// ['r1(4,)', 'y1(4,)', 'r1(0,)', 'y1(0,)', 'r1(12,)', 'y1(7,)', 'r1(15,)', 'y1(15,)', 'y2(108,)', 'y2(123,)', 'y2(34,)', 'r1(25,)', 'y1(117,)', 'r1(60,)', 'y1(60,)', 'r1(64,)']
// Data values: [0, 5, 1, 0, 0, 4, 1, 0, 1, 2, 5, 0, 4, 0, 1, 1]
// Dest PEs: [42, 43, 50, 51, 34, 35, 42, 43, 29, 30, 31, 34, 27, 34, 35, 42]
9'd21: rdata =   56'b00000000000000000000000000000000000000000000000000000011;
//
// shift amount: 0, Lanes IDs: [2, 3]
9'd22: rdata =   56'b00000000000000000000000000000000000011111100000001010000;
//
// shift amount: 2, Lanes IDs: [2, 3]
9'd23: rdata =   56'b00000000000000000000000000000000000010110100000001010010;
//
// shift amount: 6, Lanes IDs: [10, 11]
9'd24: rdata =   56'b00000000000010110100000000000000000000000000000001010110;
//
// shift amount: 12, Lanes IDs: [10, 11]
9'd25: rdata =   56'b00000000000010110100000000000000000000000000000001011100;
//
// read [True, True, False, False]
// ['r1(20,)', 'y1(20,)', 'r2(10,)', 'r1(1,)', 'r1(2,)', 'y1(2,)', 'y2(10,)', 'r1(8,)', 'y2(108,)', 'y2(123,)', 'y2(34,)', 'r1(25,)', 'y1(117,)', 'r1(60,)', 'y1(60,)', 'r1(64,)']
// Data values: [0, 5, 0, 1, 1, 0, 0, 0, 1, 2, 5, 0, 4, 0, 1, 1]
// Dest PEs: [53, 54, 55, 58, 50, 51, 55, 58, 29, 30, 31, 34, 27, 34, 35, 42]
9'd26: rdata =   56'b00000000000000000000000000000000000000000000000000000011;
//
// shift amount: 2, Lanes IDs: [2, 3]
9'd27: rdata =   56'b00000000000000000000000000000000000011111100000001010010;
//
// shift amount: 9, Lanes IDs: [10]
9'd28: rdata =   56'b00000000000000011100000000000000000000000000000001011001;
//
// shift amount: 11, Lanes IDs: [5, 6, 7]
9'd29: rdata =   56'b00000000000000000000000011111111100000000000000001011011;
//
// shift amount: 13, Lanes IDs: [10]
9'd30: rdata =   56'b00000000000000011100000000000000000000000000000001011101;
//
// shift amount: 15, Lanes IDs: [7]
9'd31: rdata =   56'b00000000000000000000000011100000000000000000000001011111;
//
// read [True, True, False, False]
// ['y1(1,)', 'r1(85,)', 'r2(11,)', 'r2(26,)', 'y1(8,)', 'y1(85,)', 'y2(11,)', 'y2(26,)', 'y2(108,)', 'y2(123,)', 'y2(34,)', 'r1(25,)', 'y1(117,)', 'r1(60,)', 'y1(60,)', 'r1(64,)']
// Data values: [0, 1, 0, 0, 2, 1, 1, 2, 1, 2, 5, 0, 4, 0, 1, 1]
// Dest PEs: [59, 61, 62, 63, 59, 61, 62, 63, 29, 30, 31, 34, 27, 34, 35, 42]
9'd32: rdata =   56'b00000000000000000000000000000000000000000000000000000011;
//
// shift amount: 4, Lanes IDs: [13, 14, 15]
9'd33: rdata =   56'b11111111100000000000000000000000000000000000000001010100;
//
// shift amount: 8, Lanes IDs: [13, 14, 15]
9'd34: rdata =   56'b11111111100000000000000000000000000000000000000001011000;
//
// shift amount: 5, Lanes IDs: [11]
9'd35: rdata =   56'b00000000000011100000000000000000000000000000000001010101;
//
// shift amount: 9, Lanes IDs: [11]
9'd36: rdata =   56'b00000000000011100000000000000000000000000000000001011001;
//
// read [True, False, False, False]
// ['r1(6,)', 'r1(3,)', 'r1(21,)', 'y1(21,)', 'r1(9,)', 'y1(3,)', 'r1(30,)', 'y1(105,)', 'y2(108,)', 'y2(123,)', 'y2(34,)', 'r1(25,)', 'y1(117,)', 'r1(60,)', 'y1(60,)', 'r1(64,)']
// Data values: [1, 0, 0, 4, 0, 1, 1, 2, 1, 2, 5, 0, 4, 0, 1, 1]
// Dest PEs: [2, 3, 4, 5, 2, 3, 4, 6, 29, 30, 31, 34, 27, 34, 35, 42]
9'd37: rdata =   56'b00000000000000000000000000000000000000000000000000000001;
//
// shift amount: 14, Lanes IDs: [2, 3, 4, 5]
9'd38: rdata =   56'b00000000000000000000000000000000100100100100000001011110;
//
// read [True, True, False, False]
// ['r1(105,)', 'r1(5,)', 'r1(133,)', 'r2(88,)', 'r1(9,)', 'y1(3,)', 'r1(30,)', 'y1(105,)', 'y2(108,)', 'y2(123,)', 'y2(34,)', 'r1(25,)', 'y1(117,)', 'r1(60,)', 'y1(60,)', 'r1(64,)']
// Data values: [0, 1, 0, 1, 0, 1, 1, 2, 1, 2, 5, 0, 4, 0, 1, 1]
// Dest PEs: [6, 10, 11, 12, 2, 3, 4, 6, 29, 30, 31, 34, 27, 34, 35, 42]
9'd39: rdata =   56'b00000000000000000000000000000000000000000000000000000011;
//
// shift amount: 10, Lanes IDs: [6]
9'd40: rdata =   56'b00000000000000000000000000000100000000000000000001011010;
//
// shift amount: 1, Lanes IDs: [6]
9'd41: rdata =   56'b00000000000000000000000000000100000000000000000001010001;
//
// shift amount: 2, Lanes IDs: [2, 3, 4]
9'd42: rdata =   56'b00000000000000000000000000000000000100100100000001010010;
//
// shift amount: 7, Lanes IDs: [10, 11, 12]
9'd43: rdata =   56'b00000000000100100100000000000000000000000000000001010111;
//
// read [True, True, False, False]
// ['r1(26,)', 'r1(17,)', 'r1(39,)', 'r1(126,)', 'r1(11,)', 'r1(135,)', 'y1(133,)', 'r1(32,)', 'y2(108,)', 'y2(123,)', 'y2(34,)', 'r1(25,)', 'y1(117,)', 'r1(60,)', 'y1(60,)', 'r1(64,)']
// Data values: [0, 1, 1, 1, 0, 0, 2, 1, 1, 2, 5, 0, 4, 0, 1, 1]
// Dest PEs: [13, 14, 15, 17, 10, 11, 12, 13, 29, 30, 31, 34, 27, 34, 35, 42]
9'd44: rdata =   56'b00000000000000000000000000000000000000000000000000000011;
//
// shift amount: 2, Lanes IDs: [1]
9'd45: rdata =   56'b00000000000000000000000000000000000000000001100001010010;
//
// shift amount: 3, Lanes IDs: [13, 14, 15]
9'd46: rdata =   56'b00100100100000000000000000000000000000000000000001010011;
//
// shift amount: 10, Lanes IDs: [10, 11, 12, 13]
9'd47: rdata =   56'b00000000100100100100000000000000000000000000000001011010;
//
// read [True, True, False, False]
// ['r1(33,)', 'r1(27,)', 'r1(119,)', 'r1(61,)', 'y1(17,)', 'r1(56,)', 'y1(126,)', 'r1(38,)', 'y2(108,)', 'y2(123,)', 'y2(34,)', 'r1(25,)', 'y1(117,)', 'r1(60,)', 'y1(60,)', 'r1(64,)']
// Data values: [1, 1, 1, 0, 4, 1, 1, 0, 1, 2, 5, 0, 4, 0, 1, 1]
// Dest PEs: [18, 19, 20, 21, 14, 15, 17, 18, 29, 30, 31, 34, 27, 34, 35, 42]
9'd48: rdata =   56'b00000000000000000000000000000000000000000000000000000011;
//
// shift amount: 14, Lanes IDs: [2, 3, 4, 5]
9'd49: rdata =   56'b00000000000000000000000000000001101101101100000001011110;
//
// shift amount: 5, Lanes IDs: [1, 2]
9'd50: rdata =   56'b00000000000000000000000000000000000000001101100001010101;
//
// shift amount: 6, Lanes IDs: [14, 15]
9'd51: rdata =   56'b00100100000000000000000000000000000000000000000001010110;
//
// read [True, True, False, False]
// ['r1(73,)', 'r1(84,)', 'r1(71,)', 'r2(120,)', 'r1(58,)', 'r1(130,)', 'r1(100,)', 'r1(91,)', 'y2(108,)', 'y2(123,)', 'y2(34,)', 'r1(25,)', 'y1(117,)', 'r1(60,)', 'y1(60,)', 'r1(64,)']
// Data values: [0, 1, 0, 0, 0, 1, 0, 0, 1, 2, 5, 0, 4, 0, 1, 1]
// Dest PEs: [22, 23, 26, 27, 19, 20, 21, 22, 29, 30, 31, 34, 27, 34, 35, 42]
9'd52: rdata =   56'b00000000000000000000000000000000000000000000000000000011;
//
// shift amount: 8, Lanes IDs: [10, 11]
9'd53: rdata =   56'b00000000000001101100000000000000000000000000000001011000;
//
// shift amount: 10, Lanes IDs: [6, 7]
9'd54: rdata =   56'b00000000000000000000000001101100000000000000000001011010;
//
// shift amount: 1, Lanes IDs: [3, 4, 5, 6]
9'd55: rdata =   56'b00000000000000000000000000001101101101100000000001010001;
//
// read [False, True, False, False]
// ['r1(81,)', 'y1(81,)', 'r1(75,)', 'y1(57,)', 'r2(119,)', 'r1(79,)', 'y1(54,)', 'y1(82,)', 'y2(108,)', 'y2(123,)', 'y2(34,)', 'r1(25,)', 'y1(117,)', 'r1(60,)', 'y1(60,)', 'r1(64,)']
// Data values: [0, 3, 1, 2, 1, 0, 0, 4, 1, 2, 5, 0, 4, 0, 1, 1]
// Dest PEs: [58, 59, 2, 3, 23, 26, 27, 28, 29, 30, 31, 34, 27, 34, 35, 42]
9'd56: rdata =   56'b00000000000000000000000000000000000000000000000000000010;
//
// shift amount: 11, Lanes IDs: [10, 11, 12]
9'd57: rdata =   56'b00000000001101101100000000000000000000000000000001011011;
//
// shift amount: 13, Lanes IDs: [7]
9'd58: rdata =   56'b00000000000000000000000001100000000000000000000001011101;
//
// read [False, True, True, False]
// ['r1(81,)', 'y1(81,)', 'r1(75,)', 'y1(57,)', 'y1(112,)', 'y2(2,)', 'y1(34,)', 'r1(19,)', 'y2(108,)', 'y2(123,)', 'y2(34,)', 'r1(25,)', 'y1(117,)', 'r1(60,)', 'y1(60,)', 'r1(64,)']
// Data values: [0, 3, 1, 2, 5, 4, 4, 1, 1, 2, 5, 0, 4, 0, 1, 1]
// Dest PEs: [58, 59, 2, 3, 29, 30, 31, 34, 29, 30, 31, 34, 27, 34, 35, 42]
9'd59: rdata =   56'b00000000000000000000000000000000000000000000000000000110;
//
// shift amount: 5, Lanes IDs: [2]
9'd60: rdata =   56'b00000000000000000000000000000000000000010100000001010101;
//
// shift amount: 9, Lanes IDs: [2]
9'd61: rdata =   56'b00000000000000000000000000000000000000010100000001011001;
//
// shift amount: 7, Lanes IDs: [13, 14, 15]
9'd62: rdata =   56'b01101101100000000000000000000000000000000000000001010111;
//
// shift amount: 11, Lanes IDs: [13, 14, 15]
9'd63: rdata =   56'b01101101100000000000000000000000000000000000000001011011;
//
// read [False, True, True, False]
// ['r1(81,)', 'y1(81,)', 'r1(75,)', 'y1(57,)', 'y1(12,)', 'r1(28,)', 'y1(28,)', 'r1(13,)', 'y1(19,)', 'r1(41,)', 'y1(41,)', 'r1(16,)', 'y1(117,)', 'r1(60,)', 'y1(60,)', 'r1(64,)']
// Data values: [0, 3, 1, 2, 5, 1, 4, 0, 5, 1, 0, 0, 4, 0, 1, 1]
// Dest PEs: [58, 59, 2, 3, 35, 42, 43, 50, 35, 42, 43, 50, 27, 34, 35, 42]
9'd64: rdata =   56'b00000000000000000000000000000000000000000000000000000110;
//
// shift amount: 1, Lanes IDs: [3]
9'd65: rdata =   56'b00000000000000000000000000000000000010100000000001010001;
//
// shift amount: 5, Lanes IDs: [2, 3]
9'd66: rdata =   56'b00000000000000000000000000000000000010111100000001010101;
//
// shift amount: 9, Lanes IDs: [2]
9'd67: rdata =   56'b00000000000000000000000000000000000000011100000001011001;
//
// shift amount: 11, Lanes IDs: [10, 11]
9'd68: rdata =   56'b00000000000010110100000000000000000000000000000001011011;
//
// shift amount: 15, Lanes IDs: [10, 11]
9'd69: rdata =   56'b00000000000010110100000000000000000000000000000001011111;
//
// read [False, True, True, False]
// ['r1(81,)', 'y1(81,)', 'r1(75,)', 'y1(57,)', 'y1(13,)', 'r1(14,)', 'y1(14,)', 'r1(10,)', 'y1(16,)', 'r1(23,)', 'y1(23,)', 'r1(24,)', 'y1(117,)', 'r1(60,)', 'y1(60,)', 'r1(64,)']
// Data values: [0, 3, 1, 2, 1, 1, 0, 0, 0, 1, 0, 0, 4, 0, 1, 1]
// Dest PEs: [58, 59, 2, 3, 51, 58, 59, 2, 51, 58, 59, 2, 27, 34, 35, 42]
9'd70: rdata =   56'b00000000000000000000000000000000000000000000000000000110;
//
// shift amount: 1, Lanes IDs: [3]
9'd71: rdata =   56'b00000000000000000000000000000000000011100000000001010001;
//
// shift amount: 5, Lanes IDs: [2, 3]
9'd72: rdata =   56'b00000000000000000000000000000000000011100100000001010101;
//
// shift amount: 9, Lanes IDs: [2]
9'd73: rdata =   56'b00000000000000000000000000000000000000000100000001011001;
//
// shift amount: 11, Lanes IDs: [10, 11]
9'd74: rdata =   56'b00000000000011111100000000000000000000000000000001011011;
//
// shift amount: 15, Lanes IDs: [10, 11]
9'd75: rdata =   56'b00000000000011111100000000000000000000000000000001011111;
//
// read [False, True, False, False]
// ['r1(81,)', 'y1(81,)', 'r1(75,)', 'y1(57,)', 'y1(6,)', 'y1(30,)', 'r1(18,)', 'y1(5,)', 'y1(9,)', 'r1(31,)', 'y1(11,)', 'y2(88,)', 'y1(117,)', 'r1(60,)', 'y1(60,)', 'r1(64,)']
// Data values: [0, 3, 1, 2, 3, 1, 1, 4, 5, 1, 3, 0, 4, 0, 1, 1]
// Dest PEs: [58, 59, 2, 3, 3, 4, 10, 11, 3, 10, 11, 12, 27, 34, 35, 42]
9'd76: rdata =   56'b00000000000000000000000000000000000000000000000000000010;
//
// shift amount: 1, Lanes IDs: [3, 4]
9'd77: rdata =   56'b00000000000000000000000000000000000100100000000001010001;
//
// shift amount: 12, Lanes IDs: [10, 11]
9'd78: rdata =   56'b00000000000000100100000000000000000000000000000001011100;
//
// read [False, True, True, False]
// ['r1(81,)', 'y1(81,)', 'r1(75,)', 'y1(57,)', 'y1(135,)', 'y1(26,)', 'y1(39,)', 'r1(44,)', 'y1(9,)', 'r1(31,)', 'y1(11,)', 'y2(88,)', 'y1(117,)', 'r1(60,)', 'y1(60,)', 'r1(64,)']
// Data values: [0, 3, 1, 2, 4, 2, 1, 1, 5, 1, 3, 0, 4, 0, 1, 1]
// Dest PEs: [58, 59, 2, 3, 12, 13, 15, 18, 3, 10, 11, 12, 27, 34, 35, 42]
9'd79: rdata =   56'b00000000000000000000000000000000000000000000000000000110;
//
// shift amount: 8, Lanes IDs: [12, 13]
9'd80: rdata =   56'b00000000100100000000000000000000000000000000000001011000;
//
// shift amount: 15, Lanes IDs: [10, 11, 12]
9'd81: rdata =   56'b00000000000100100100000000000000000000000000000001011111;
//
// shift amount: 5, Lanes IDs: [2, 3]
9'd82: rdata =   56'b00000000000000000000000000000000000000101100000001010101;
//
// shift amount: 7, Lanes IDs: [15]
9'd83: rdata =   56'b00100000000000000000000000000000000000000000000001010111;
//
// read [False, True, True, False]
// ['r1(81,)', 'y1(81,)', 'r1(75,)', 'y1(57,)', 'r1(123,)', 'r2(12,)', 'r2(19,)', 'r1(131,)', 'y1(32,)', 'y1(56,)', 'r1(51,)', 'r1(124,)', 'y1(117,)', 'r1(60,)', 'y1(60,)', 'r1(64,)']
// Data values: [0, 3, 1, 2, 0, 1, 0, 1, 4, 4, 0, 1, 4, 0, 1, 1]
// Dest PEs: [58, 59, 2, 3, 19, 20, 21, 22, 13, 15, 18, 19, 27, 34, 35, 42]
9'd84: rdata =   56'b00000000000000000000000000000000000000000000000000000110;
//
// shift amount: 1, Lanes IDs: [3, 4, 5, 6]
9'd85: rdata =   56'b00000000000000000000000000001101101101100000000001010001;
//
// shift amount: 8, Lanes IDs: [2, 3]
9'd86: rdata =   56'b00000000000000000000000000000000000001101100000001011000;
//
// shift amount: 10, Lanes IDs: [15]
9'd87: rdata =   56'b00100000000000000000000000000000000000000000000001011010;
//
// shift amount: 11, Lanes IDs: [13]
9'd88: rdata =   56'b00000000100000000000000000000000000000000000000001011011;
//
// read [False, True, True, False]
// ['r1(81,)', 'y1(81,)', 'r1(75,)', 'y1(57,)', 'y2(119,)', 'r1(107,)', 'y1(71,)', 'y2(60,)', 'r2(122,)', 'r2(25,)', 'r2(48,)', 'r1(117,)', 'y1(117,)', 'r1(60,)', 'y1(60,)', 'r1(64,)']
// Data values: [0, 3, 1, 2, 5, 0, 2, 0, 1, 0, 0, 1, 4, 0, 1, 1]
// Dest PEs: [58, 59, 2, 3, 23, 26, 27, 28, 20, 21, 22, 26, 27, 34, 35, 42]
9'd89: rdata =   56'b00000000000000000000000000000000000000000000000000000110;
//
// shift amount: 11, Lanes IDs: [10, 11, 12]
9'd90: rdata =   56'b00000000001101101100000000000000000000000000000001011011;
//
// shift amount: 1, Lanes IDs: [10]
9'd91: rdata =   56'b00000000000000001100000000000000000000000000000001010001;
//
// shift amount: 4, Lanes IDs: [4, 5, 6]
9'd92: rdata =   56'b00000000000000000000000000001101101100000000000001010100;
//
// shift amount: 13, Lanes IDs: [7]
9'd93: rdata =   56'b00000000000000000000000001100000000000000000000001011101;
//
// read [False, False, True, False]
// ['r1(81,)', 'y1(81,)', 'r1(75,)', 'y1(57,)', 'y1(44,)', 'y2(78,)', 'y2(12,)', 'y2(19,)', 'y1(79,)', 'y2(120,)', 'y2(39,)', 'r1(42,)', 'y1(117,)', 'r1(60,)', 'y1(60,)', 'r1(64,)']
// Data values: [0, 3, 1, 2, 2, 3, 1, 3, 1, 1, 4, 0, 4, 0, 1, 1]
// Dest PEs: [58, 59, 2, 3, 19, 20, 21, 22, 27, 28, 31, 34, 27, 34, 35, 42]
9'd94: rdata =   56'b00000000000000000000000000000000000000000000000000000100;
//
// shift amount: 9, Lanes IDs: [2]
9'd95: rdata =   56'b00000000000000000000000000000000000000010100000001011001;
//
// shift amount: 11, Lanes IDs: [15]
9'd96: rdata =   56'b01100000000000000000000000000000000000000000000001011011;
//
// shift amount: 13, Lanes IDs: [11, 12]
9'd97: rdata =   56'b00000000001101100000000000000000000000000000000001011101;
//
// read [False, False, True, False]
// ['r1(81,)', 'y1(81,)', 'r1(75,)', 'y1(57,)', 'y1(44,)', 'y2(78,)', 'y2(12,)', 'y2(19,)', 'y1(42,)', 'r1(49,)', 'y1(49,)', 'r1(29,)', 'y1(117,)', 'r1(60,)', 'y1(60,)', 'r1(64,)']
// Data values: [0, 3, 1, 2, 2, 3, 1, 3, 3, 1, 0, 1, 4, 0, 1, 1]
// Dest PEs: [58, 59, 2, 3, 19, 20, 21, 22, 35, 42, 43, 50, 27, 34, 35, 42]
9'd98: rdata =   56'b00000000000000000000000000000000000000000000000000000100;
//
// shift amount: 9, Lanes IDs: [2]
9'd99: rdata =   56'b00000000000000000000000000000000000000011100000001011001;
//
// shift amount: 5, Lanes IDs: [3]
9'd100: rdata =  56'b00000000000000000000000000000000000010100000000001010101;
//
// shift amount: 15, Lanes IDs: [10, 11]
9'd101: rdata =  56'b00000000000010110100000000000000000000000000000001011111;
//
// read [False, False, True, False]
// ['r1(81,)', 'y1(81,)', 'r1(75,)', 'y1(57,)', 'y1(44,)', 'y2(78,)', 'y2(12,)', 'y2(19,)', 'y1(29,)', 'r1(37,)', 'y1(37,)', 'r1(40,)', 'y1(117,)', 'r1(60,)', 'y1(60,)', 'r1(64,)']
// Data values: [0, 3, 1, 2, 2, 3, 1, 3, 2, 1, 2, 0, 4, 0, 1, 1]
// Dest PEs: [58, 59, 2, 3, 19, 20, 21, 22, 51, 58, 59, 2, 27, 34, 35, 42]
9'd102: rdata =  56'b00000000000000000000000000000000000000000000000000000100;
//
// shift amount: 9, Lanes IDs: [2]
9'd103: rdata =  56'b00000000000000000000000000000000000000000100000001011001;
//
// shift amount: 5, Lanes IDs: [3]
9'd104: rdata =  56'b00000000000000000000000000000000000011100000000001010101;
//
// shift amount: 15, Lanes IDs: [10, 11]
9'd105: rdata =  56'b00000000000011111100000000000000000000000000000001011111;
//
// read [False, False, True, False]
// ['r1(81,)', 'y1(81,)', 'r1(75,)', 'y1(57,)', 'y1(44,)', 'y2(78,)', 'y2(12,)', 'y2(19,)', 'y1(10,)', 'r1(36,)', 'y1(18,)', 'r1(59,)', 'y1(117,)', 'r1(60,)', 'y1(60,)', 'r1(64,)']
// Data values: [0, 3, 1, 2, 2, 3, 1, 3, 5, 0, 1, 0, 4, 0, 1, 1]
// Dest PEs: [58, 59, 2, 3, 19, 20, 21, 22, 3, 10, 11, 18, 27, 34, 35, 42]
9'd106: rdata =  56'b00000000000000000000000000000000000000000000000000000100;
//
// shift amount: 9, Lanes IDs: [2]
9'd107: rdata =  56'b00000000000000000000000000000000000000001100000001011001;
//
// shift amount: 5, Lanes IDs: [3]
9'd108: rdata =  56'b00000000000000000000000000000000000000100000000001010101;
//
// shift amount: 15, Lanes IDs: [10, 11]
9'd109: rdata =  56'b00000000000000100100000000000000000000000000000001011111;
//
// read [False, False, True, False]
// ['r1(81,)', 'y1(81,)', 'r1(75,)', 'y1(57,)', 'y1(44,)', 'y2(78,)', 'y2(12,)', 'y2(19,)', 'r1(129,)', 'r2(126,)', 'r2(99,)', 'r2(121,)', 'y1(117,)', 'r1(60,)', 'y1(60,)', 'r1(64,)']
// Data values: [0, 3, 1, 2, 2, 3, 1, 3, 1, 1, 1, 0, 4, 0, 1, 1]
// Dest PEs: [58, 59, 2, 3, 19, 20, 21, 22, 19, 20, 21, 22, 27, 34, 35, 42]
9'd110: rdata =  56'b00000000000000000000000000000000000000000000000000000100;
//
// shift amount: 5, Lanes IDs: [3, 4, 5, 6]
9'd111: rdata =  56'b00000000000000000000000000001101101101100000000001010101;
//
// read [False, False, True, False]
// ['r1(81,)', 'y1(81,)', 'r1(75,)', 'y1(57,)', 'y1(44,)', 'y2(78,)', 'y2(12,)', 'y2(19,)', 'r2(7,)', 'y1(107,)', 'r1(48,)', 'y1(48,)', 'y1(117,)', 'r1(60,)', 'y1(60,)', 'r1(64,)']
// Data values: [0, 3, 1, 2, 2, 3, 1, 3, 0, 5, 1, 3, 4, 0, 1, 1]
// Dest PEs: [58, 59, 2, 3, 19, 20, 21, 22, 26, 27, 34, 35, 27, 34, 35, 42]
9'd112: rdata =  56'b00000000000000000000000000000000000000000000000000000100;
//
// shift amount: 8, Lanes IDs: [2, 3]
9'd113: rdata =  56'b00000000000000000000000000000000000010110100000001011000;
//
// shift amount: 14, Lanes IDs: [10, 11]
9'd114: rdata =  56'b00000000000001101100000000000000000000000000000001011110;
//
// read [False, False, True, True]
// ['r1(81,)', 'y1(81,)', 'r1(75,)', 'y1(57,)', 'y1(44,)', 'y2(78,)', 'y2(12,)', 'y2(19,)', 'r1(62,)', 'y1(62,)', 'r1(35,)', 'y1(35,)', 'y1(117,)', 'r1(60,)', 'y1(60,)', 'r1(64,)']
// Data values: [0, 3, 1, 2, 2, 3, 1, 3, 1, 1, 0, 5, 4, 0, 1, 1]
// Dest PEs: [58, 59, 2, 3, 19, 20, 21, 22, 42, 43, 50, 51, 27, 34, 35, 42]
9'd115: rdata =  56'b00000000000000000000000000000000000000000000000000001100;
//
// shift amount: 1, Lanes IDs: [11]
9'd116: rdata =  56'b00000000000001100000000000000000000000000000000001010001;
//
// shift amount: 8, Lanes IDs: [2, 3]
9'd117: rdata =  56'b00000000000000000000000000000000000011111100000001011000;
//
// shift amount: 11, Lanes IDs: [2, 3]
9'd118: rdata =  56'b00000000000000000000000000000000000010110100000001011011;
//
// shift amount: 14, Lanes IDs: [10, 11]
9'd119: rdata =  56'b00000000000010110100000000000000000000000000000001011110;
//
// shift amount: 5, Lanes IDs: [10]
9'd120: rdata =  56'b00000000000000010100000000000000000000000000000001010101;
//
// read [False, False, True, True]
// ['r1(81,)', 'y1(81,)', 'r1(75,)', 'y1(57,)', 'y1(44,)', 'y2(78,)', 'y2(12,)', 'y2(19,)', 'r1(47,)', 'y1(47,)', 'r1(43,)', 'y1(24,)', 'y1(64,)', 'r1(46,)', 'y1(46,)', 'r1(55,)']
// Data values: [0, 3, 1, 2, 2, 3, 1, 3, 0, 5, 1, 0, 1, 1, 5, 1]
// Dest PEs: [58, 59, 2, 3, 19, 20, 21, 22, 58, 59, 2, 3, 43, 50, 51, 58]
9'd121: rdata =  56'b00000000000000000000000000000000000000000000000000001100;
//
// shift amount: 1, Lanes IDs: [11]
9'd122: rdata =  56'b00000000000010100000000000000000000000000000000001010001;
//
// shift amount: 8, Lanes IDs: [2, 3]
9'd123: rdata =  56'b00000000000000000000000000000000000000100100000001011000;
//
// shift amount: 11, Lanes IDs: [2, 3]
9'd124: rdata =  56'b00000000000000000000000000000000000011111100000001011011;
//
// shift amount: 14, Lanes IDs: [10, 11]
9'd125: rdata =  56'b00000000000011111100000000000000000000000000000001011110;
//
// shift amount: 5, Lanes IDs: [10]
9'd126: rdata =  56'b00000000000000011100000000000000000000000000000001010101;
//
// read [False, False, True, True]
// ['r1(81,)', 'y1(81,)', 'r1(75,)', 'y1(57,)', 'y1(44,)', 'y2(78,)', 'y2(12,)', 'y2(19,)', 'r1(45,)', 'y1(31,)', 'r1(74,)', 'r2(6,)', 'y1(55,)', 'r1(52,)', 'y1(40,)', 'r1(50,)']
// Data values: [0, 3, 1, 2, 2, 3, 1, 3, 0, 1, 0, 1, 1, 1, 0, 0]
// Dest PEs: [58, 59, 2, 3, 19, 20, 21, 22, 10, 11, 18, 19, 59, 2, 3, 10]
9'd127: rdata =  56'b00000000000000000000000000000000000000000000000000001100;
//
// shift amount: 1, Lanes IDs: [11]
9'd128: rdata =  56'b00000000000011100000000000000000000000000000000001010001;
//
// shift amount: 8, Lanes IDs: [2, 3]
9'd129: rdata =  56'b00000000000000000000000000000000000001101100000001011000;
//
// shift amount: 11, Lanes IDs: [2, 3]
9'd130: rdata =  56'b00000000000000000000000000000000000000100100000001011011;
//
// shift amount: 14, Lanes IDs: [10, 11]
9'd131: rdata =  56'b00000000000000100100000000000000000000000000000001011110;
//
// shift amount: 5, Lanes IDs: [10]
9'd132: rdata =  56'b00000000000000000100000000000000000000000000000001010101;
//
// read [False, False, True, True]
// ['r1(81,)', 'y1(81,)', 'r1(75,)', 'y1(57,)', 'y1(44,)', 'y2(78,)', 'y2(12,)', 'y2(19,)', 'y1(58,)', 'r2(118,)', 'r2(124,)', 'r2(8,)', 'y1(36,)', 'r1(78,)', 'r2(66,)', 'y1(118,)']
// Data values: [0, 3, 1, 2, 2, 3, 1, 3, 3, 1, 0, 0, 0, 0, 1, 2]
// Dest PEs: [58, 59, 2, 3, 19, 20, 21, 22, 20, 21, 22, 26, 11, 18, 19, 20]
9'd133: rdata =  56'b00000000000000000000000000000000000000000000000000001100;
//
// shift amount: 1, Lanes IDs: [10, 11]
9'd134: rdata =  56'b00000000000000101100000000000000000000000000000001010001;
//
// shift amount: 4, Lanes IDs: [4, 5, 6]
9'd135: rdata =  56'b00000000000000000000000000001101101100000000000001010100;
//
// shift amount: 11, Lanes IDs: [2, 3, 4]
9'd136: rdata =  56'b00000000000000000000000000000000001101101100000001011011;
//
// read [False, False, False, True]
// ['r1(81,)', 'y1(81,)', 'r1(75,)', 'y1(57,)', 'y1(44,)', 'y2(78,)', 'y2(12,)', 'y2(19,)', 'r2(29,)', 'y2(29,)', 'r2(37,)', 'y2(37,)', 'r2(125,)', 'y1(22,)', 'r2(17,)', 'y2(7,)']
// Data values: [0, 3, 1, 2, 2, 3, 1, 3, 1, 5, 1, 1, 0, 4, 0, 2]
// Dest PEs: [58, 59, 2, 3, 19, 20, 21, 22, 50, 51, 58, 59, 21, 22, 26, 27]
9'd137: rdata =  56'b00000000000000000000000000000000000000000000000000001000;
//
// shift amount: 4, Lanes IDs: [10, 11]
9'd138: rdata =  56'b00000000000001101100000000000000000000000000000001010100;
//
// shift amount: 7, Lanes IDs: [5, 6]
9'd139: rdata =  56'b00000000000000000000000000001101100000000000000001010111;
//
// read [False, False, False, True]
// ['r1(81,)', 'y1(81,)', 'r1(75,)', 'y1(57,)', 'y1(44,)', 'y2(78,)', 'y2(12,)', 'y2(19,)', 'r2(29,)', 'y2(29,)', 'r2(37,)', 'y2(37,)', 'r1(80,)', 'y1(80,)', 'r1(72,)', 'y1(72,)']
// Data values: [0, 3, 1, 2, 2, 3, 1, 3, 1, 5, 1, 1, 0, 3, 1, 2]
// Dest PEs: [58, 59, 2, 3, 19, 20, 21, 22, 50, 51, 58, 59, 34, 35, 42, 43]
9'd140: rdata =  56'b00000000000000000000000000000000000000000000000000001000;
//
// shift amount: 10, Lanes IDs: [2, 3]
9'd141: rdata =  56'b00000000000000000000000000000000000010110100000001011010;
//
// shift amount: 4, Lanes IDs: [10, 11]
9'd142: rdata =  56'b00000000000010110100000000000000000000000000000001010100;
//
// read [False, False, False, True]
// ['r1(81,)', 'y1(81,)', 'r1(75,)', 'y1(57,)', 'y1(44,)', 'y2(78,)', 'y2(12,)', 'y2(19,)', 'r2(29,)', 'y2(29,)', 'r2(37,)', 'y2(37,)', 'r1(53,)', 'y1(53,)', 'r1(66,)', 'y1(66,)']
// Data values: [0, 3, 1, 2, 2, 3, 1, 3, 1, 5, 1, 1, 1, 3, 1, 3]
// Dest PEs: [58, 59, 2, 3, 19, 20, 21, 22, 50, 51, 58, 59, 50, 51, 58, 59]
9'd143: rdata =  56'b00000000000000000000000000000000000000000000000000001000;
//
// shift amount: 10, Lanes IDs: [2, 3]
9'd144: rdata =  56'b00000000000000000000000000000000000011111100000001011010;
//
// shift amount: 4, Lanes IDs: [10, 11]
9'd145: rdata =  56'b00000000000011111100000000000000000000000000000001010100;
//
// read [False, False, False, True]
// ['r1(81,)', 'y1(81,)', 'r1(75,)', 'y1(57,)', 'y1(44,)', 'y2(78,)', 'y2(12,)', 'y2(19,)', 'r2(29,)', 'y2(29,)', 'r2(37,)', 'y2(37,)', 'r1(57,)', 'y1(43,)', 'r1(63,)', 'y1(45,)']
// Data values: [0, 3, 1, 2, 2, 3, 1, 3, 1, 5, 1, 1, 1, 4, 0, 0]
// Dest PEs: [58, 59, 2, 3, 19, 20, 21, 22, 50, 51, 58, 59, 2, 3, 10, 11]
9'd146: rdata =  56'b00000000000000000000000000000000000000000000000000001000;
//
// shift amount: 10, Lanes IDs: [2, 3]
9'd147: rdata =  56'b00000000000000000000000000000000000000100100000001011010;
//
// shift amount: 4, Lanes IDs: [10, 11]
9'd148: rdata =  56'b00000000000000100100000000000000000000000000000001010100;
//
// read [False, False, False, True]
// ['r1(81,)', 'y1(81,)', 'r1(75,)', 'y1(57,)', 'y1(44,)', 'y2(78,)', 'y2(12,)', 'y2(19,)', 'r2(29,)', 'y2(29,)', 'r2(37,)', 'y2(37,)', 'r1(90,)', 'r2(78,)', 'y1(119,)', 'y1(61,)']
// Data values: [0, 3, 1, 2, 2, 3, 1, 3, 1, 5, 1, 1, 0, 1, 5, 2]
// Dest PEs: [58, 59, 2, 3, 19, 20, 21, 22, 50, 51, 58, 59, 18, 19, 20, 21]
9'd149: rdata =  56'b00000000000000000000000000000000000000000000000000001000;
//
// shift amount: 10, Lanes IDs: [2, 3, 4, 5]
9'd150: rdata =  56'b00000000000000000000000000000001101101101100000001011010;
//
// read [False, False, False, True]
// ['r1(81,)', 'y1(81,)', 'r1(75,)', 'y1(57,)', 'y1(44,)', 'y2(78,)', 'y2(12,)', 'y2(19,)', 'r2(29,)', 'y2(29,)', 'r2(37,)', 'y2(37,)', 'y1(73,)', 'r2(21,)', 'y2(8,)', 'r1(86,)']
// Data values: [0, 3, 1, 2, 2, 3, 1, 3, 1, 5, 1, 1, 1, 0, 1, 0]
// Dest PEs: [58, 59, 2, 3, 19, 20, 21, 22, 50, 51, 58, 59, 22, 26, 27, 34]
9'd151: rdata =  56'b00000000000000000000000000000000000000000000000000001000;
//
// shift amount: 3, Lanes IDs: [10, 11]
9'd152: rdata =  56'b00000000000001101100000000000000000000000000000001010011;
//
// shift amount: 13, Lanes IDs: [2]
9'd153: rdata =  56'b00000000000000000000000000000000000000010100000001011101;
//
// shift amount: 6, Lanes IDs: [6]
9'd154: rdata =  56'b00000000000000000000000000001100000000000000000001010110;
//
// read [False, False, False, True]
// ['r1(81,)', 'y1(81,)', 'r1(75,)', 'y1(57,)', 'y1(44,)', 'y2(78,)', 'y2(12,)', 'y2(19,)', 'r2(29,)', 'y2(29,)', 'r2(37,)', 'y2(37,)', 'y1(86,)', 'r1(88,)', 'y1(88,)', 'r1(65,)']
// Data values: [0, 3, 1, 2, 2, 3, 1, 3, 1, 5, 1, 1, 2, 1, 0, 1]
// Dest PEs: [58, 59, 2, 3, 19, 20, 21, 22, 50, 51, 58, 59, 35, 42, 43, 50]
9'd155: rdata =  56'b00000000000000000000000000000000000000000000000000001000;
//
// shift amount: 9, Lanes IDs: [3]
9'd156: rdata =  56'b00000000000000000000000000000000000010100000000001011001;
//
// shift amount: 3, Lanes IDs: [10, 11]
9'd157: rdata =  56'b00000000000010110100000000000000000000000000000001010011;
//
// shift amount: 13, Lanes IDs: [2]
9'd158: rdata =  56'b00000000000000000000000000000000000000011100000001011101;
//
// read [False, False, False, True]
// ['r1(81,)', 'y1(81,)', 'r1(75,)', 'y1(57,)', 'y1(44,)', 'y2(78,)', 'y2(12,)', 'y2(19,)', 'r2(29,)', 'y2(29,)', 'r2(37,)', 'y2(37,)', 'y1(65,)', 'r1(68,)', 'y1(68,)', 'r1(67,)']
// Data values: [0, 3, 1, 2, 2, 3, 1, 3, 1, 5, 1, 1, 3, 1, 2, 1]
// Dest PEs: [58, 59, 2, 3, 19, 20, 21, 22, 50, 51, 58, 59, 51, 58, 59, 2]
9'd159: rdata =  56'b00000000000000000000000000000000000000000000000000001000;
//
// shift amount: 9, Lanes IDs: [3]
9'd160: rdata =  56'b00000000000000000000000000000000000011100000000001011001;
//
// shift amount: 3, Lanes IDs: [10, 11]
9'd161: rdata =  56'b00000000000011111100000000000000000000000000000001010011;
//
// shift amount: 13, Lanes IDs: [2]
9'd162: rdata =  56'b00000000000000000000000000000000000000000100000001011101;
//
// read [False, False, False, True]
// ['r1(81,)', 'y1(81,)', 'r1(75,)', 'y1(57,)', 'y1(44,)', 'y2(78,)', 'y2(12,)', 'y2(19,)', 'r2(29,)', 'y2(29,)', 'r2(37,)', 'y2(37,)', 'y1(52,)', 'r1(69,)', 'y1(50,)', 'r1(96,)']
// Data values: [0, 3, 1, 2, 2, 3, 1, 3, 1, 5, 1, 1, 4, 1, 4, 1]
// Dest PEs: [58, 59, 2, 3, 19, 20, 21, 22, 50, 51, 58, 59, 3, 10, 11, 18]
9'd163: rdata =  56'b00000000000000000000000000000000000000000000000000001000;
//
// shift amount: 9, Lanes IDs: [3]
9'd164: rdata =  56'b00000000000000000000000000000000000000100000000001011001;
//
// shift amount: 3, Lanes IDs: [10, 11]
9'd165: rdata =  56'b00000000000000100100000000000000000000000000000001010011;
//
// shift amount: 13, Lanes IDs: [2]
9'd166: rdata =  56'b00000000000000000000000000000000000000001100000001011101;
//
// read [True, False, False, True]
// ['r1(81,)', 'y1(81,)', 'r1(75,)', 'y1(57,)', 'y1(44,)', 'y2(78,)', 'y2(12,)', 'y2(19,)', 'r2(29,)', 'y2(29,)', 'r2(37,)', 'y2(37,)', 'r2(127,)', 'y1(123,)', 'y1(100,)', 'y1(91,)']
// Data values: [0, 3, 1, 2, 2, 3, 1, 3, 1, 5, 1, 1, 1, 2, 0, 1]
// Dest PEs: [58, 59, 2, 3, 19, 20, 21, 22, 50, 51, 58, 59, 19, 20, 21, 22]
9'd167: rdata =  56'b00000000000000000000000000000000000000000000000000001001;
//
// shift amount: 0, Lanes IDs: [2, 3]
9'd168: rdata =  56'b00000000000000000000000000000000000000100100000001010000;
//
// shift amount: 9, Lanes IDs: [3, 4, 5, 6]
9'd169: rdata =  56'b00000000000000000000000000001101101101100000000001011001;
//
// shift amount: 6, Lanes IDs: [10, 11]
9'd170: rdata =  56'b00000000000011111100000000000000000000000000000001010110;
//
// read [True, False, False, True]
// ['r1(70,)', 'y1(63,)', 'r1(108,)', 'r2(128,)', 'y1(44,)', 'y2(78,)', 'y2(12,)', 'y2(19,)', 'r2(29,)', 'y2(29,)', 'r2(37,)', 'y2(37,)', 'r2(27,)', 'y2(17,)', 'r1(92,)', 'y1(92,)']
// Data values: [1, 0, 0, 0, 2, 3, 1, 3, 1, 5, 1, 1, 1, 5, 0, 2]
// Dest PEs: [10, 11, 18, 19, 19, 20, 21, 22, 50, 51, 58, 59, 26, 27, 34, 35]
9'd171: rdata =  56'b00000000000000000000000000000000000000000000000000001001;
//
// shift amount: 0, Lanes IDs: [2, 3]
9'd172: rdata =  56'b00000000000000000000000000000000000001101100000001010000;
//
// shift amount: 2, Lanes IDs: [10, 11]
9'd173: rdata =  56'b00000000000001101100000000000000000000000000000001010010;
//
// shift amount: 12, Lanes IDs: [2, 3]
9'd174: rdata =  56'b00000000000000000000000000000000000010110100000001011100;
//
// shift amount: 6, Lanes IDs: [10, 11]
9'd175: rdata =  56'b00000000000000100100000000000000000000000000000001010110;
//
// read [True, False, False, True]
// ['y1(124,)', 'y1(108,)', 'y1(121,)', 'r2(32,)', 'y1(44,)', 'y2(78,)', 'y2(12,)', 'y2(19,)', 'r2(29,)', 'y2(29,)', 'r2(37,)', 'y2(37,)', 'r1(93,)', 'y1(93,)', 'r1(87,)', 'y1(87,)']
// Data values: [2, 2, 2, 0, 2, 3, 1, 3, 1, 5, 1, 1, 0, 2, 0, 3]
// Dest PEs: [20, 21, 22, 26, 19, 20, 21, 22, 50, 51, 58, 59, 42, 43, 50, 51]
9'd176: rdata =  56'b00000000000000000000000000000000000000000000000000001001;
//
// shift amount: 9, Lanes IDs: [10]
9'd177: rdata =  56'b00000000000000001100000000000000000000000000000001011001;
//
// shift amount: 2, Lanes IDs: [10, 11]
9'd178: rdata =  56'b00000000000010110100000000000000000000000000000001010010;
//
// shift amount: 12, Lanes IDs: [2, 3, 4, 5, 6]
9'd179: rdata =  56'b00000000000000000000000000001101101111111100000001011100;
//
// read [True, False, False, False]
// ['y2(21,)', 'r1(99,)', 'y1(99,)', 'r1(98,)', 'y1(44,)', 'y2(78,)', 'y2(12,)', 'y2(19,)', 'r2(29,)', 'y2(29,)', 'r2(37,)', 'y2(37,)', 'r2(61,)', 'y2(42,)', 'r2(51,)', 'y1(137,)']
// Data values: [5, 1, 3, 0, 2, 3, 1, 3, 1, 5, 1, 1, 0, 4, 0, 4]
// Dest PEs: [27, 34, 35, 42, 19, 20, 21, 22, 50, 51, 58, 59, 2, 3, 10, 11]
9'd180: rdata =  56'b00000000000000000000000000000000000000000000000000000001;
//
// shift amount: 9, Lanes IDs: [10]
9'd181: rdata =  56'b00000000000000010100000000000000000000000000000001011001;
//
// shift amount: 5, Lanes IDs: [11]
9'd182: rdata =  56'b00000000000001100000000000000000000000000000000001010101;
//
// shift amount: 15, Lanes IDs: [2, 3]
9'd183: rdata =  56'b00000000000000000000000000000000000010110100000001011111;
//
// read [True, False, False, False]
// ['y1(98,)', 'r1(94,)', 'y1(94,)', 'r1(95,)', 'y1(44,)', 'y2(78,)', 'y2(12,)', 'y2(19,)', 'r2(29,)', 'y2(29,)', 'r2(37,)', 'y2(37,)', 'r2(61,)', 'y2(42,)', 'r2(51,)', 'y1(137,)']
// Data values: [0, 0, 4, 0, 2, 3, 1, 3, 1, 5, 1, 1, 0, 4, 0, 4]
// Dest PEs: [43, 50, 51, 58, 19, 20, 21, 22, 50, 51, 58, 59, 2, 3, 10, 11]
9'd184: rdata =  56'b00000000000000000000000000000000000000000000000000000001;
//
// shift amount: 9, Lanes IDs: [10]
9'd185: rdata =  56'b00000000000000011100000000000000000000000000000001011001;
//
// shift amount: 5, Lanes IDs: [11]
9'd186: rdata =  56'b00000000000010100000000000000000000000000000000001010101;
//
// shift amount: 15, Lanes IDs: [2, 3]
9'd187: rdata =  56'b00000000000000000000000000000000000011111100000001011111;
//
// read [True, False, False, False]
// ['y1(95,)', 'r1(89,)', 'y1(67,)', 'r1(76,)', 'y1(44,)', 'y2(78,)', 'y2(12,)', 'y2(19,)', 'r2(29,)', 'y2(29,)', 'r2(37,)', 'y2(37,)', 'r2(61,)', 'y2(42,)', 'r2(51,)', 'y1(137,)']
// Data values: [0, 1, 5, 0, 2, 3, 1, 3, 1, 5, 1, 1, 0, 4, 0, 4]
// Dest PEs: [59, 2, 3, 10, 19, 20, 21, 22, 50, 51, 58, 59, 2, 3, 10, 11]
9'd188: rdata =  56'b00000000000000000000000000000000000000000000000000000001;
//
// shift amount: 9, Lanes IDs: [10]
9'd189: rdata =  56'b00000000000000000100000000000000000000000000000001011001;
//
// shift amount: 5, Lanes IDs: [11]
9'd190: rdata =  56'b00000000000011100000000000000000000000000000000001010101;
//
// shift amount: 15, Lanes IDs: [2, 3]
9'd191: rdata =  56'b00000000000000000000000000000000000000100100000001011111;
//
// read [True, False, False, False]
// ['y1(69,)', 'r1(118,)', 'r2(129,)', 'y1(129,)', 'y1(44,)', 'y2(78,)', 'y2(12,)', 'y2(19,)', 'r2(29,)', 'y2(29,)', 'r2(37,)', 'y2(37,)', 'r2(61,)', 'y2(42,)', 'r2(51,)', 'y1(137,)']
// Data values: [1, 0, 0, 3, 2, 3, 1, 3, 1, 5, 1, 1, 0, 4, 0, 4]
// Dest PEs: [11, 18, 19, 20, 19, 20, 21, 22, 50, 51, 58, 59, 2, 3, 10, 11]
9'd192: rdata =  56'b00000000000000000000000000000000000000000000000000000001;
//
// shift amount: 5, Lanes IDs: [11]
9'd193: rdata =  56'b00000000000000100000000000000000000000000000000001010101;
//
// shift amount: 15, Lanes IDs: [2, 3, 4]
9'd194: rdata =  56'b00000000000000000000000000000000001101101100000001011111;
//
// read [True, False, False, False]
// ['y1(130,)', 'y1(131,)', 'r2(54,)', 'y2(27,)', 'y1(44,)', 'y2(78,)', 'y2(12,)', 'y2(19,)', 'r2(29,)', 'y2(29,)', 'r2(37,)', 'y2(37,)', 'r2(61,)', 'y2(42,)', 'r2(51,)', 'y1(137,)']
// Data values: [4, 4, 1, 3, 2, 3, 1, 3, 1, 5, 1, 1, 0, 4, 0, 4]
// Dest PEs: [21, 22, 26, 27, 19, 20, 21, 22, 50, 51, 58, 59, 2, 3, 10, 11]
9'd195: rdata =  56'b00000000000000000000000000000000000000000000000000000001;
//
// shift amount: 8, Lanes IDs: [10, 11]
9'd196: rdata =  56'b00000000000001101100000000000000000000000000000001011000;
//
// shift amount: 11, Lanes IDs: [5, 6]
9'd197: rdata =  56'b00000000000000000000000000001101100000000000000001011011;
//
// read [True, False, False, False]
// ['r1(110,)', 'y1(110,)', 'r1(109,)', 'y1(109,)', 'y1(44,)', 'y2(78,)', 'y2(12,)', 'y2(19,)', 'r2(29,)', 'y2(29,)', 'r2(37,)', 'y2(37,)', 'r2(61,)', 'y2(42,)', 'r2(51,)', 'y1(137,)']
// Data values: [1, 4, 0, 1, 2, 3, 1, 3, 1, 5, 1, 1, 0, 4, 0, 4]
// Dest PEs: [34, 35, 42, 43, 19, 20, 21, 22, 50, 51, 58, 59, 2, 3, 10, 11]
9'd198: rdata =  56'b00000000000000000000000000000000000000000000000000000001;
//
// shift amount: 8, Lanes IDs: [10, 11]
9'd199: rdata =  56'b00000000000010110100000000000000000000000000000001011000;
//
// shift amount: 14, Lanes IDs: [2, 3]
9'd200: rdata =  56'b00000000000000000000000000000000000010110100000001011110;
//
// read [True, False, False, False]
// ['r1(101,)', 'y1(101,)', 'r1(106,)', 'y1(106,)', 'y1(44,)', 'y2(78,)', 'y2(12,)', 'y2(19,)', 'r2(29,)', 'y2(29,)', 'r2(37,)', 'y2(37,)', 'r2(61,)', 'y2(42,)', 'r2(51,)', 'y1(137,)']
// Data values: [0, 0, 0, 1, 2, 3, 1, 3, 1, 5, 1, 1, 0, 4, 0, 4]
// Dest PEs: [50, 51, 58, 59, 19, 20, 21, 22, 50, 51, 58, 59, 2, 3, 10, 11]
9'd201: rdata =  56'b00000000000000000000000000000000000000000000000000000001;
//
// shift amount: 8, Lanes IDs: [10, 11]
9'd202: rdata =  56'b00000000000011111100000000000000000000000000000001011000;
//
// shift amount: 14, Lanes IDs: [2, 3]
9'd203: rdata =  56'b00000000000000000000000000000000000011111100000001011110;
//
// read [True, False, False, False]
// ['r1(97,)', 'y1(75,)', 'r1(83,)', 'y1(70,)', 'y1(44,)', 'y2(78,)', 'y2(12,)', 'y2(19,)', 'r2(29,)', 'y2(29,)', 'r2(37,)', 'y2(37,)', 'r2(61,)', 'y2(42,)', 'r2(51,)', 'y1(137,)']
// Data values: [1, 2, 0, 0, 2, 3, 1, 3, 1, 5, 1, 1, 0, 4, 0, 4]
// Dest PEs: [2, 3, 10, 11, 19, 20, 21, 22, 50, 51, 58, 59, 2, 3, 10, 11]
9'd204: rdata =  56'b00000000000000000000000000000000000000000000000000000001;
//
// shift amount: 8, Lanes IDs: [10, 11]
9'd205: rdata =  56'b00000000000000100100000000000000000000000000000001011000;
//
// shift amount: 14, Lanes IDs: [2, 3]
9'd206: rdata =  56'b00000000000000000000000000000000000000100100000001011110;
//
// read [True, False, False, False]
// ['r1(121,)', 'y1(27,)', 'y2(66,)', 'y2(6,)', 'y1(44,)', 'y2(78,)', 'y2(12,)', 'y2(19,)', 'r2(29,)', 'y2(29,)', 'r2(37,)', 'y2(37,)', 'r2(61,)', 'y2(42,)', 'r2(51,)', 'y1(137,)']
// Data values: [0, 4, 3, 0, 2, 3, 1, 3, 1, 5, 1, 1, 0, 4, 0, 4]
// Dest PEs: [18, 19, 20, 21, 19, 20, 21, 22, 50, 51, 58, 59, 2, 3, 10, 11]
9'd207: rdata =  56'b00000000000000000000000000000000000000000000000000000001;
//
// shift amount: 14, Lanes IDs: [2, 3, 4, 5]
9'd208: rdata =  56'b00000000000000000000000000000001101101101100000001011110;
//
// read [True, True, False, False]
// ['y2(18,)', 'r2(94,)', 'y2(32,)', 'r1(127,)', 'y1(44,)', 'y2(78,)', 'y2(12,)', 'y2(19,)', 'r2(29,)', 'y2(29,)', 'r2(37,)', 'y2(37,)', 'r2(61,)', 'y2(42,)', 'r2(51,)', 'y1(137,)']
// Data values: [2, 1, 0, 1, 2, 3, 1, 3, 1, 5, 1, 1, 0, 4, 0, 4]
// Dest PEs: [22, 26, 27, 34, 19, 20, 21, 22, 50, 51, 58, 59, 2, 3, 10, 11]
9'd209: rdata =  56'b00000000000000000000000000000000000000000000000000000011;
//
// shift amount: 10, Lanes IDs: [6]
9'd210: rdata =  56'b00000000000000000000000000001100000000000000000001011010;
//
// shift amount: 1, Lanes IDs: [2, 3, 4, 5, 6]
9'd211: rdata =  56'b00000000000000000000000000001101101101110100000001010001;
//
// shift amount: 7, Lanes IDs: [10, 11]
9'd212: rdata =  56'b00000000000001101100000000000000000000000000000001010111;
//
// read [True, True, False, False]
// ['y1(127,)', 'r1(116,)', 'y1(116,)', 'r1(113,)', 'r2(105,)', 'y2(94,)', 'r2(3,)', 'y2(3,)', 'r2(29,)', 'y2(29,)', 'r2(37,)', 'y2(37,)', 'r2(61,)', 'y2(42,)', 'r2(51,)', 'y1(137,)']
// Data values: [2, 1, 3, 1, 0, 1, 1, 5, 1, 5, 1, 1, 0, 4, 0, 4]
// Dest PEs: [35, 42, 43, 50, 26, 27, 34, 35, 50, 51, 58, 59, 2, 3, 10, 11]
9'd213: rdata =  56'b00000000000000000000000000000000000000000000000000000011;
//
// shift amount: 1, Lanes IDs: [2]
9'd214: rdata =  56'b00000000000000000000000000000000000000011100000001010001;
//
// shift amount: 7, Lanes IDs: [10, 11]
9'd215: rdata =  56'b00000000000010110100000000000000000000000000000001010111;
//
// shift amount: 10, Lanes IDs: [10, 11]
9'd216: rdata =  56'b00000000000001101100000000000000000000000000000001011010;
//
// shift amount: 13, Lanes IDs: [3]
9'd217: rdata =  56'b00000000000000000000000000000000000010100000000001011101;
//
// shift amount: 4, Lanes IDs: [2, 3]
9'd218: rdata =  56'b00000000000000000000000000000000000010110100000001010100;
//
// read [True, True, False, False]
// ['y1(113,)', 'r1(114,)', 'y1(114,)', 'r1(104,)', 'r2(1,)', 'y2(1,)', 'r1(120,)', 'y1(120,)', 'r2(29,)', 'y2(29,)', 'r2(37,)', 'y2(37,)', 'r2(61,)', 'y2(42,)', 'r2(51,)', 'y1(137,)']
// Data values: [2, 1, 1, 0, 1, 4, 1, 1, 1, 5, 1, 1, 0, 4, 0, 4]
// Dest PEs: [51, 58, 59, 2, 42, 43, 50, 51, 50, 51, 58, 59, 2, 3, 10, 11]
9'd219: rdata =  56'b00000000000000000000000000000000000000000000000000000011;
//
// shift amount: 1, Lanes IDs: [2]
9'd220: rdata =  56'b00000000000000000000000000000000000000000100000001010001;
//
// shift amount: 7, Lanes IDs: [10, 11]
9'd221: rdata =  56'b00000000000011111100000000000000000000000000000001010111;
//
// shift amount: 10, Lanes IDs: [10, 11]
9'd222: rdata =  56'b00000000000010110100000000000000000000000000000001011010;
//
// shift amount: 13, Lanes IDs: [3]
9'd223: rdata =  56'b00000000000000000000000000000000000011100000000001011101;
//
// shift amount: 4, Lanes IDs: [2, 3]
9'd224: rdata =  56'b00000000000000000000000000000000000011111100000001010100;
//
// read [True, True, False, False]
// ['y1(89,)', 'r1(103,)', 'y1(76,)', 'r1(128,)', 'r1(134,)', 'y1(134,)', 'r1(115,)', 'y1(97,)', 'r2(29,)', 'y2(29,)', 'r2(37,)', 'y2(37,)', 'r2(61,)', 'y2(42,)', 'r2(51,)', 'y1(137,)']
// Data values: [0, 1, 1, 0, 1, 5, 1, 3, 1, 5, 1, 1, 0, 4, 0, 4]
// Dest PEs: [3, 10, 11, 18, 58, 59, 2, 3, 50, 51, 58, 59, 2, 3, 10, 11]
9'd225: rdata =  56'b00000000000000000000000000000000000000000000000000000011;
//
// shift amount: 1, Lanes IDs: [2]
9'd226: rdata =  56'b00000000000000000000000000000000000000001100000001010001;
//
// shift amount: 7, Lanes IDs: [10, 11]
9'd227: rdata =  56'b00000000000000100100000000000000000000000000000001010111;
//
// shift amount: 10, Lanes IDs: [10, 11]
9'd228: rdata =  56'b00000000000011111100000000000000000000000000000001011010;
//
// shift amount: 13, Lanes IDs: [3]
9'd229: rdata =  56'b00000000000000000000000000000000000000100000000001011101;
//
// shift amount: 4, Lanes IDs: [2, 3]
9'd230: rdata =  56'b00000000000000000000000000000000000000100100000001010100;
//
// read [False, True, False, False]
// ['r2(107,)', 'y2(107,)', 'r2(106,)', 'y2(106,)', 'r1(111,)', 'y1(83,)', 'r2(18,)', 'y1(59,)', 'r2(29,)', 'y2(29,)', 'r2(37,)', 'y2(37,)', 'r2(61,)', 'y2(42,)', 'r2(51,)', 'y1(137,)']
// Data values: [1, 0, 1, 0, 1, 5, 1, 4, 1, 5, 1, 1, 0, 4, 0, 4]
// Dest PEs: [42, 43, 50, 51, 10, 11, 18, 19, 50, 51, 58, 59, 2, 3, 10, 11]
9'd231: rdata =  56'b00000000000000000000000000000000000000000000000000000010;
//
// shift amount: 10, Lanes IDs: [10, 11]
9'd232: rdata =  56'b00000000000000100100000000000000000000000000000001011010;
//
// shift amount: 4, Lanes IDs: [2, 3]
9'd233: rdata =  56'b00000000000000000000000000000000000001101100000001010100;
//
// read [False, True, False, False]
// ['r2(107,)', 'y2(107,)', 'r2(106,)', 'y2(106,)', 'y2(128,)', 'y2(25,)', 'y2(48,)', 'r2(117,)', 'r2(29,)', 'y2(29,)', 'r2(37,)', 'y2(37,)', 'r2(61,)', 'y2(42,)', 'r2(51,)', 'y1(137,)']
// Data values: [1, 0, 1, 0, 2, 5, 1, 0, 1, 5, 1, 1, 0, 4, 0, 4]
// Dest PEs: [42, 43, 50, 51, 20, 21, 22, 26, 50, 51, 58, 59, 2, 3, 10, 11]
9'd234: rdata =  56'b00000000000000000000000000000000000000000000000000000010;
//
// shift amount: 0, Lanes IDs: [4, 5, 6]
9'd235: rdata =  56'b00000000000000000000000000001101101100000000000001010000;
//
// shift amount: 13, Lanes IDs: [10]
9'd236: rdata =  56'b00000000000000001100000000000000000000000000000001011101;
//
// read [False, True, False, False]
// ['r2(107,)', 'y2(107,)', 'r2(106,)', 'y2(106,)', 'y2(105,)', 'r2(5,)', 'y2(5,)', 'r2(9,)', 'r2(29,)', 'y2(29,)', 'r2(37,)', 'y2(37,)', 'r2(61,)', 'y2(42,)', 'r2(51,)', 'y1(137,)']
// Data values: [1, 0, 1, 0, 1, 0, 0, 1, 1, 5, 1, 1, 0, 4, 0, 4]
// Dest PEs: [42, 43, 50, 51, 27, 34, 35, 42, 50, 51, 58, 59, 2, 3, 10, 11]
9'd237: rdata =  56'b00000000000000000000000000000000000000000000000000000010;
//
// shift amount: 9, Lanes IDs: [11]
9'd238: rdata =  56'b00000000000001100000000000000000000000000000000001011001;
//
// shift amount: 3, Lanes IDs: [2, 3]
9'd239: rdata =  56'b00000000000000000000000000000000000010110100000001010011;
//
// shift amount: 13, Lanes IDs: [10]
9'd240: rdata =  56'b00000000000000010100000000000000000000000000000001011101;
//
// read [False, True, False, False]
// ['r2(107,)', 'y2(107,)', 'r2(106,)', 'y2(106,)', 'y2(9,)', 'r2(4,)', 'y2(4,)', 'r2(14,)', 'r2(29,)', 'y2(29,)', 'r2(37,)', 'y2(37,)', 'r2(61,)', 'y2(42,)', 'r2(51,)', 'y1(137,)']
// Data values: [1, 0, 1, 0, 5, 1, 2, 1, 1, 5, 1, 1, 0, 4, 0, 4]
// Dest PEs: [42, 43, 50, 51, 43, 50, 51, 58, 50, 51, 58, 59, 2, 3, 10, 11]
9'd241: rdata =  56'b00000000000000000000000000000000000000000000000000000010;
//
// shift amount: 9, Lanes IDs: [11]
9'd242: rdata =  56'b00000000000010100000000000000000000000000000000001011001;
//
// shift amount: 3, Lanes IDs: [2, 3]
9'd243: rdata =  56'b00000000000000000000000000000000000011111100000001010011;
//
// shift amount: 13, Lanes IDs: [10]
9'd244: rdata =  56'b00000000000000011100000000000000000000000000000001011101;
//
// read [False, True, False, False]
// ['r2(107,)', 'y2(107,)', 'r2(106,)', 'y2(106,)', 'y2(14,)', 'r2(0,)', 'y1(104,)', 'r1(122,)', 'r2(29,)', 'y2(29,)', 'r2(37,)', 'y2(37,)', 'r2(61,)', 'y2(42,)', 'r2(51,)', 'y1(137,)']
// Data values: [1, 0, 1, 0, 0, 1, 1, 1, 1, 5, 1, 1, 0, 4, 0, 4]
// Dest PEs: [42, 43, 50, 51, 59, 2, 3, 10, 50, 51, 58, 59, 2, 3, 10, 11]
9'd245: rdata =  56'b00000000000000000000000000000000000000000000000000000010;
//
// shift amount: 9, Lanes IDs: [11]
9'd246: rdata =  56'b00000000000011100000000000000000000000000000000001011001;
//
// shift amount: 3, Lanes IDs: [2, 3]
9'd247: rdata =  56'b00000000000000000000000000000000000000100100000001010011;
//
// shift amount: 13, Lanes IDs: [10]
9'd248: rdata =  56'b00000000000000000100000000000000000000000000000001011101;
//
// read [False, True, False, False]
// ['r2(107,)', 'y2(107,)', 'r2(106,)', 'y2(106,)', 'y1(103,)', 'r2(28,)', 'y1(74,)', 'y2(129,)', 'r2(29,)', 'y2(29,)', 'r2(37,)', 'y2(37,)', 'r2(61,)', 'y2(42,)', 'r2(51,)', 'y1(137,)']
// Data values: [1, 0, 1, 0, 2, 1, 4, 1, 1, 5, 1, 1, 0, 4, 0, 4]
// Dest PEs: [42, 43, 50, 51, 11, 18, 19, 20, 50, 51, 58, 59, 2, 3, 10, 11]
9'd249: rdata =  56'b00000000000000000000000000000000000000000000000000000010;
//
// shift amount: 9, Lanes IDs: [11]
9'd250: rdata =  56'b00000000000000100000000000000000000000000000000001011001;
//
// shift amount: 3, Lanes IDs: [2, 3, 4]
9'd251: rdata =  56'b00000000000000000000000000000000001101101100000001010011;
//
// read [False, True, False, False]
// ['r2(107,)', 'y2(107,)', 'r2(106,)', 'y2(106,)', 'y2(99,)', 'y2(118,)', 'y2(54,)', 'y2(117,)', 'r2(29,)', 'y2(29,)', 'r2(37,)', 'y2(37,)', 'r2(61,)', 'y2(42,)', 'r2(51,)', 'y1(137,)']
// Data values: [1, 0, 1, 0, 2, 3, 1, 4, 1, 5, 1, 1, 0, 4, 0, 4]
// Dest PEs: [42, 43, 50, 51, 21, 22, 26, 27, 50, 51, 58, 59, 2, 3, 10, 11]
9'd252: rdata =  56'b00000000000000000000000000000000000000000000000000000010;
//
// shift amount: 12, Lanes IDs: [10, 11]
9'd253: rdata =  56'b00000000000001101100000000000000000000000000000001011100;
//
// shift amount: 15, Lanes IDs: [5, 6]
9'd254: rdata =  56'b00000000000000000000000000001101100000000000000001011111;
//
// read [False, True, False, False]
// ['r2(107,)', 'y2(107,)', 'r2(106,)', 'y2(106,)', 'r2(24,)', 'y2(24,)', 'r2(13,)', 'y2(13,)', 'r2(29,)', 'y2(29,)', 'r2(37,)', 'y2(37,)', 'r2(61,)', 'y2(42,)', 'r2(51,)', 'y1(137,)']
// Data values: [1, 0, 1, 0, 0, 2, 1, 1, 1, 5, 1, 1, 0, 4, 0, 4]
// Dest PEs: [42, 43, 50, 51, 34, 35, 42, 43, 50, 51, 58, 59, 2, 3, 10, 11]
9'd255: rdata =  56'b00000000000000000000000000000000000000000000000000000010;
//
// shift amount: 2, Lanes IDs: [2, 3]
9'd256: rdata =  56'b00000000000000000000000000000000000010110100000001010010;
//
// shift amount: 12, Lanes IDs: [10, 11]
9'd257: rdata =  56'b00000000000010110100000000000000000000000000000001011100;
//
// read [False, True, True, False]
// ['r2(107,)', 'y2(107,)', 'r2(106,)', 'y2(106,)', 'r2(20,)', 'y2(20,)', 'r2(15,)', 'y2(15,)', 'r2(29,)', 'y2(29,)', 'r2(37,)', 'y2(37,)', 'r2(61,)', 'y2(42,)', 'r2(51,)', 'y1(137,)']
// Data values: [1, 0, 1, 0, 1, 5, 0, 0, 1, 5, 1, 1, 0, 4, 0, 4]
// Dest PEs: [42, 43, 50, 51, 50, 51, 58, 59, 50, 51, 58, 59, 2, 3, 10, 11]
9'd258: rdata =  56'b00000000000000000000000000000000000000000000000000000110;
//
// shift amount: 2, Lanes IDs: [2, 3]
9'd259: rdata =  56'b00000000000000000000000000000000000011111100000001010010;
//
// shift amount: 12, Lanes IDs: [10, 11]
9'd260: rdata =  56'b00000000000011111100000000000000000000000000000001011100;
//
// shift amount: 0, Lanes IDs: [10, 11]
9'd261: rdata =  56'b00000000000011111100000000000000000000000000000001010000;
//
// shift amount: 6, Lanes IDs: [2, 3]
9'd262: rdata =  56'b00000000000000000000000000000000000011111100000001010110;
//
// read [False, True, True, False]
// ['r2(107,)', 'y2(107,)', 'r2(106,)', 'y2(106,)', 'r2(16,)', 'y1(115,)', 'r1(125,)', 'y1(111,)', 'r2(22,)', 'y2(0,)', 'r1(132,)', 'y1(122,)', 'r2(61,)', 'y2(42,)', 'r2(51,)', 'y1(137,)']
// Data values: [1, 0, 1, 0, 1, 2, 1, 3, 0, 2, 0, 3, 0, 4, 0, 4]
// Dest PEs: [42, 43, 50, 51, 2, 3, 10, 11, 2, 3, 10, 11, 2, 3, 10, 11]
9'd263: rdata =  56'b00000000000000000000000000000000000000000000000000000110;
//
// shift amount: 2, Lanes IDs: [2, 3]
9'd264: rdata =  56'b00000000000000000000000000000000000000100100000001010010;
//
// shift amount: 12, Lanes IDs: [10, 11]
9'd265: rdata =  56'b00000000000000100100000000000000000000000000000001011100;
//
// shift amount: 0, Lanes IDs: [10, 11]
9'd266: rdata =  56'b00000000000000100100000000000000000000000000000001010000;
//
// shift amount: 6, Lanes IDs: [2, 3]
9'd267: rdata =  56'b00000000000000000000000000000000000000100100000001010110;
//
// read [False, True, True, False]
// ['r2(107,)', 'y2(107,)', 'r2(106,)', 'y2(106,)', 'r2(38,)', 'y1(78,)', 'y2(122,)', 'y2(121,)', 'r2(47,)', 'y1(84,)', 'y2(125,)', 'y2(124,)', 'r2(61,)', 'y2(42,)', 'r2(51,)', 'y1(137,)']
// Data values: [1, 0, 1, 0, 0, 5, 3, 1, 0, 3, 1, 2, 0, 4, 0, 4]
// Dest PEs: [42, 43, 50, 51, 18, 19, 21, 22, 18, 19, 21, 22, 2, 3, 10, 11]
9'd268: rdata =  56'b00000000000000000000000000000000000000000000000000000110;
//
// shift amount: 1, Lanes IDs: [5, 6]
9'd269: rdata =  56'b00000000000000000000000000001101100000000000000001010001;
//
// shift amount: 2, Lanes IDs: [2, 3]
9'd270: rdata =  56'b00000000000000000000000000000000000001101100000001010010;
//
// shift amount: 5, Lanes IDs: [5, 6]
9'd271: rdata =  56'b00000000000000000000000000001101100000000000000001010101;
//
// shift amount: 6, Lanes IDs: [2, 3]
9'd272: rdata =  56'b00000000000000000000000000000000000001101100000001010110;
//
// read [False, True, True, False]
// ['r2(107,)', 'y2(107,)', 'r2(106,)', 'y2(106,)', 'r2(31,)', 'y2(31,)', 'r2(23,)', 'y2(23,)', 'r2(35,)', 'y2(35,)', 'r2(33,)', 'y2(33,)', 'r2(61,)', 'y2(42,)', 'r2(51,)', 'y1(137,)']
// Data values: [1, 0, 1, 0, 1, 1, 1, 2, 0, 1, 0, 5, 0, 4, 0, 4]
// Dest PEs: [42, 43, 50, 51, 34, 35, 42, 43, 34, 35, 42, 43, 2, 3, 10, 11]
9'd273: rdata =  56'b00000000000000000000000000000000000000000000000000000110;
//
// shift amount: 2, Lanes IDs: [2, 3]
9'd274: rdata =  56'b00000000000000000000000000000000000010110100000001010010;
//
// shift amount: 12, Lanes IDs: [10, 11]
9'd275: rdata =  56'b00000000000010110100000000000000000000000000000001011100;
//
// shift amount: 0, Lanes IDs: [10, 11]
9'd276: rdata =  56'b00000000000010110100000000000000000000000000000001010000;
//
// shift amount: 6, Lanes IDs: [2, 3]
9'd277: rdata =  56'b00000000000000000000000000000000000010110100000001010110;
//
// read [False, False, True, False]
// ['r2(107,)', 'y2(107,)', 'r2(106,)', 'y2(106,)', None, None, None, None, 'r2(36,)', 'y2(36,)', 'r2(46,)', 'y2(46,)', 'r2(61,)', 'y2(42,)', 'r2(51,)', 'y1(137,)']
// Data values: [1, 0, 1, 0, None, None, None, None, 0, 4, 0, 4, 0, 4, 0, 4]
// Dest PEs: [42, 43, 50, 51, None, None, None, None, 50, 51, 58, 59, 2, 3, 10, 11]
9'd278: rdata =  56'b00000000000000000000000000000000000000000000000000000100;
//
// shift amount: 0, Lanes IDs: [10, 11]
9'd279: rdata =  56'b00000000000011111100000000000000000000000000000001010000;
//
// shift amount: 6, Lanes IDs: [2, 3]
9'd280: rdata =  56'b00000000000000000000000000000000000011111100000001010110;
//
// read [False, False, True, False]
// ['r2(107,)', 'y2(107,)', 'r2(106,)', 'y2(106,)', None, None, None, None, 'r2(30,)', 'y2(16,)', 'r1(136,)', 'y1(125,)', 'r2(61,)', 'y2(42,)', 'r2(51,)', 'y1(137,)']
// Data values: [1, 0, 1, 0, None, None, None, None, 1, 1, 0, 3, 0, 4, 0, 4]
// Dest PEs: [42, 43, 50, 51, None, None, None, None, 2, 3, 10, 11, 2, 3, 10, 11]
9'd281: rdata =  56'b00000000000000000000000000000000000000000000000000000100;
//
// shift amount: 0, Lanes IDs: [10, 11]
9'd282: rdata =  56'b00000000000000100100000000000000000000000000000001010000;
//
// shift amount: 6, Lanes IDs: [2, 3]
9'd283: rdata =  56'b00000000000000000000000000000000000000100100000001010110;
//
// read [False, False, True, False]
// ['r2(107,)', 'y2(107,)', 'r2(106,)', 'y2(106,)', None, None, None, None, 'r2(52,)', 'y1(90,)', 'y2(126,)', 'y2(127,)', 'r2(61,)', 'y2(42,)', 'r2(51,)', 'y1(137,)']
// Data values: [1, 0, 1, 0, None, None, None, None, 0, 1, 2, 1, 0, 4, 0, 4]
// Dest PEs: [42, 43, 50, 51, None, None, None, None, 18, 19, 21, 22, 2, 3, 10, 11]
9'd284: rdata =  56'b00000000000000000000000000000000000000000000000000000100;
//
// shift amount: 5, Lanes IDs: [5, 6]
9'd285: rdata =  56'b00000000000000000000000000001101100000000000000001010101;
//
// shift amount: 6, Lanes IDs: [2, 3]
9'd286: rdata =  56'b00000000000000000000000000000000000001101100000001010110;
//
// read [False, False, True, False]
// ['r2(107,)', 'y2(107,)', 'r2(106,)', 'y2(106,)', None, None, None, None, 'r2(40,)', 'y2(40,)', 'r2(41,)', 'y2(41,)', 'r2(61,)', 'y2(42,)', 'r2(51,)', 'y1(137,)']
// Data values: [1, 0, 1, 0, None, None, None, None, 0, 3, 0, 2, 0, 4, 0, 4]
// Dest PEs: [42, 43, 50, 51, None, None, None, None, 34, 35, 42, 43, 2, 3, 10, 11]
9'd287: rdata =  56'b00000000000000000000000000000000000000000000000000000100;
//
// shift amount: 0, Lanes IDs: [10, 11]
9'd288: rdata =  56'b00000000000010110100000000000000000000000000000001010000;
//
// shift amount: 6, Lanes IDs: [2, 3]
9'd289: rdata =  56'b00000000000000000000000000000000000010110100000001010110;
//
// read [False, False, True, False]
// ['r2(107,)', 'y2(107,)', 'r2(106,)', 'y2(106,)', None, None, None, None, 'r2(45,)', 'y2(45,)', 'r2(59,)', 'y2(59,)', 'r2(61,)', 'y2(42,)', 'r2(51,)', 'y1(137,)']
// Data values: [1, 0, 1, 0, None, None, None, None, 1, 3, 0, 5, 0, 4, 0, 4]
// Dest PEs: [42, 43, 50, 51, None, None, None, None, 50, 51, 58, 59, 2, 3, 10, 11]
9'd290: rdata =  56'b00000000000000000000000000000000000000000000000000000100;
//
// shift amount: 0, Lanes IDs: [10, 11]
9'd291: rdata =  56'b00000000000011111100000000000000000000000000000001010000;
//
// shift amount: 6, Lanes IDs: [2, 3]
9'd292: rdata =  56'b00000000000000000000000000000000000011111100000001010110;
//
// read [False, False, True, False]
// ['r2(107,)', 'y2(107,)', 'r2(106,)', 'y2(106,)', None, None, None, None, 'r2(42,)', 'y2(22,)', 'r1(137,)', 'y1(132,)', 'r2(61,)', 'y2(42,)', 'r2(51,)', 'y1(137,)']
// Data values: [1, 0, 1, 0, None, None, None, None, 0, 0, 0, 2, 0, 4, 0, 4]
// Dest PEs: [42, 43, 50, 51, None, None, None, None, 2, 3, 10, 11, 2, 3, 10, 11]
9'd293: rdata =  56'b00000000000000000000000000000000000000000000000000000100;
//
// shift amount: 0, Lanes IDs: [10, 11]
9'd294: rdata =  56'b00000000000000100100000000000000000000000000000001010000;
//
// shift amount: 6, Lanes IDs: [2, 3]
9'd295: rdata =  56'b00000000000000000000000000000000000000100100000001010110;
//
// read [False, False, True, False]
// ['r2(107,)', 'y2(107,)', 'r2(106,)', 'y2(106,)', None, None, None, None, 'r2(58,)', 'y1(96,)', 'r2(49,)', 'y2(49,)', 'r2(61,)', 'y2(42,)', 'r2(51,)', 'y1(137,)']
// Data values: [1, 0, 1, 0, None, None, None, None, 0, 3, 0, 4, 0, 4, 0, 4]
// Dest PEs: [42, 43, 50, 51, None, None, None, None, 18, 19, 34, 35, 2, 3, 10, 11]
9'd296: rdata =  56'b00000000000000000000000000000000000000000000000000000100;
//
// shift amount: 8, Lanes IDs: [2, 3]
9'd297: rdata =  56'b00000000000000000000000000000000000010110100000001011000;
//
// shift amount: 6, Lanes IDs: [2, 3]
9'd298: rdata =  56'b00000000000000000000000000000000000001101100000001010110;
//
// read [False, False, True, False]
// ['r2(107,)', 'y2(107,)', 'r2(106,)', 'y2(106,)', None, None, None, None, 'r2(44,)', 'y2(44,)', 'r2(56,)', 'y2(56,)', 'r2(61,)', 'y2(42,)', 'r2(51,)', 'y1(137,)']
// Data values: [1, 0, 1, 0, None, None, None, None, 0, 4, 1, 2, 0, 4, 0, 4]
// Dest PEs: [42, 43, 50, 51, None, None, None, None, 42, 43, 50, 51, 2, 3, 10, 11]
9'd299: rdata =  56'b00000000000000000000000000000000000000000000000000000100;
//
// shift amount: 8, Lanes IDs: [2, 3]
9'd300: rdata =  56'b00000000000000000000000000000000000011111100000001011000;
//
// shift amount: 14, Lanes IDs: [10, 11]
9'd301: rdata =  56'b00000000000010110100000000000000000000000000000001011110;
//
// read [False, False, True, False]
// ['r2(107,)', 'y2(107,)', 'r2(106,)', 'y2(106,)', None, None, None, None, 'r2(65,)', 'y2(65,)', 'r2(50,)', 'y2(30,)', 'r2(61,)', 'y2(42,)', 'r2(51,)', 'y1(137,)']
// Data values: [1, 0, 1, 0, None, None, None, None, 0, 3, 1, 1, 0, 4, 0, 4]
// Dest PEs: [42, 43, 50, 51, None, None, None, None, 58, 59, 2, 3, 2, 3, 10, 11]
9'd302: rdata =  56'b00000000000000000000000000000000000000000000000000000100;
//
// shift amount: 8, Lanes IDs: [2, 3]
9'd303: rdata =  56'b00000000000000000000000000000000000000100100000001011000;
//
// shift amount: 14, Lanes IDs: [10, 11]
9'd304: rdata =  56'b00000000000011111100000000000000000000000000000001011110;
//
// read [False, False, True, True]
// ['r2(107,)', 'y2(107,)', 'r2(106,)', 'y2(106,)', None, None, None, None, 'r2(43,)', 'y1(136,)', 'r2(70,)', 'y2(28,)', 'r2(61,)', 'y2(42,)', 'r2(51,)', 'y1(137,)']
// Data values: [1, 0, 1, 0, None, None, None, None, 1, 3, 0, 2, 0, 4, 0, 4]
// Dest PEs: [42, 43, 50, 51, None, None, None, None, 10, 11, 18, 19, 2, 3, 10, 11]
9'd305: rdata =  56'b00000000000000000000000000000000000000000000000000001100;
//
// shift amount: 8, Lanes IDs: [2, 3]
9'd306: rdata =  56'b00000000000000000000000000000000000001101100000001011000;
//
// shift amount: 10, Lanes IDs: [2, 3]
9'd307: rdata =  56'b00000000000000000000000000000000000000100100000001011010;
//
// shift amount: 14, Lanes IDs: [10, 11]
9'd308: rdata =  56'b00000000000000100100000000000000000000000000000001011110;
//
// shift amount: 4, Lanes IDs: [10, 11]
9'd309: rdata =  56'b00000000000000100100000000000000000000000000000001010100;
//
// read [False, False, True, True]
// ['r2(107,)', 'y2(107,)', 'r2(106,)', 'y2(106,)', None, None, None, None, 'r2(53,)', 'y2(53,)', 'r2(55,)', 'y2(55,)', 'r2(76,)', 'y2(38,)', 'r2(57,)', 'y2(57,)']
// Data values: [1, 0, 1, 0, None, None, None, None, 1, 0, 0, 3, 0, 3, 1, 1]
// Dest PEs: [42, 43, 50, 51, None, None, None, None, 34, 35, 42, 43, 18, 19, 34, 35]
9'd310: rdata =  56'b00000000000000000000000000000000000000000000000000001100;
//
// shift amount: 0, Lanes IDs: [10, 11]
9'd311: rdata =  56'b00000000000010110100000000000000000000000000000001010000;
//
// shift amount: 10, Lanes IDs: [2, 3]
9'd312: rdata =  56'b00000000000000000000000000000000000001101100000001011010;
//
// shift amount: 6, Lanes IDs: [2, 3]
9'd313: rdata =  56'b00000000000000000000000000000000000010110100000001010110;
//
// shift amount: 12, Lanes IDs: [2, 3]
9'd314: rdata =  56'b00000000000000000000000000000000000010110100000001011100;
//
// read [False, False, True, True]
// ['r2(107,)', 'y2(107,)', 'r2(106,)', 'y2(106,)', None, None, None, None, 'r2(64,)', 'y2(64,)', 'r2(75,)', 'y2(75,)', 'r2(63,)', 'y2(63,)', 'r2(73,)', 'y2(73,)']
// Data values: [1, 0, 1, 0, None, None, None, None, 1, 1, 1, 1, 0, 0, 0, 3]
// Dest PEs: [42, 43, 50, 51, None, None, None, None, 50, 51, 58, 59, 42, 43, 50, 51]
9'd315: rdata =  56'b00000000000000000000000000000000000000000000000000001100;
//
// shift amount: 0, Lanes IDs: [10, 11]
9'd316: rdata =  56'b00000000000011111100000000000000000000000000000001010000;
//
// shift amount: 2, Lanes IDs: [10, 11]
9'd317: rdata =  56'b00000000000010110100000000000000000000000000000001010010;
//
// shift amount: 6, Lanes IDs: [2, 3]
9'd318: rdata =  56'b00000000000000000000000000000000000011111100000001010110;
//
// shift amount: 12, Lanes IDs: [2, 3]
9'd319: rdata =  56'b00000000000000000000000000000000000011111100000001011100;
//
// read [False, False, False, True]
// ['r2(107,)', 'y2(107,)', 'r2(106,)', 'y2(106,)', None, None, None, None, None, None, None, None, 'r2(85,)', 'y2(85,)', 'r2(69,)', 'y2(50,)']
// Data values: [1, 0, 1, 0, None, None, None, None, None, None, None, None, 0, 2, 0, 3]
// Dest PEs: [42, 43, 50, 51, None, None, None, None, None, None, None, None, 58, 59, 2, 3]
9'd320: rdata =  56'b00000000000000000000000000000000000000000000000000001000;
//
// shift amount: 2, Lanes IDs: [10, 11]
9'd321: rdata =  56'b00000000000011111100000000000000000000000000000001010010;
//
// shift amount: 12, Lanes IDs: [2, 3]
9'd322: rdata =  56'b00000000000000000000000000000000000000100100000001011100;
//
// read [False, False, False, True]
// ['r2(107,)', 'y2(107,)', 'r2(106,)', 'y2(106,)', None, None, None, None, None, None, None, None, 'r2(62,)', 'y2(43,)', 'r2(77,)', 'y2(47,)']
// Data values: [1, 0, 1, 0, None, None, None, None, None, None, None, None, 1, 0, 0, 4]
// Dest PEs: [42, 43, 50, 51, None, None, None, None, None, None, None, None, 10, 11, 18, 19]
9'd323: rdata =  56'b00000000000000000000000000000000000000000000000000001000;
//
// shift amount: 2, Lanes IDs: [10, 11]
9'd324: rdata =  56'b00000000000000100100000000000000000000000000000001010010;
//
// shift amount: 12, Lanes IDs: [2, 3]
9'd325: rdata =  56'b00000000000000000000000000000000000001101100000001011100;
//
// read [False, False, False, True]
// ['r2(107,)', 'y2(107,)', 'r2(106,)', 'y2(106,)', None, None, None, None, None, None, None, None, 'r2(68,)', 'y2(68,)', 'r2(74,)', 'y2(74,)']
// Data values: [1, 0, 1, 0, None, None, None, None, None, None, None, None, 0, 2, 1, 5]
// Dest PEs: [42, 43, 50, 51, None, None, None, None, None, None, None, None, 34, 35, 42, 43]
9'd326: rdata =  56'b00000000000000000000000000000000000000000000000000001000;
//
// shift amount: 10, Lanes IDs: [2, 3]
9'd327: rdata =  56'b00000000000000000000000000000000000010110100000001011010;
//
// shift amount: 4, Lanes IDs: [10, 11]
9'd328: rdata =  56'b00000000000010110100000000000000000000000000000001010100;
//
// read [False, False, False, True]
// ['r2(107,)', 'y2(107,)', 'r2(106,)', 'y2(106,)', None, None, None, None, None, None, None, None, 'r2(80,)', 'y2(80,)', 'r2(93,)', 'y2(93,)']
// Data values: [1, 0, 1, 0, None, None, None, None, None, None, None, None, 0, 2, 0, 5]
// Dest PEs: [42, 43, 50, 51, None, None, None, None, None, None, None, None, 50, 51, 58, 59]
9'd329: rdata =  56'b00000000000000000000000000000000000000000000000000001000;
//
// shift amount: 10, Lanes IDs: [2, 3]
9'd330: rdata =  56'b00000000000000000000000000000000000011111100000001011010;
//
// shift amount: 4, Lanes IDs: [10, 11]
9'd331: rdata =  56'b00000000000011111100000000000000000000000000000001010100;
//
// read [False, False, False, True]
// ['r2(107,)', 'y2(107,)', 'r2(106,)', 'y2(106,)', None, None, None, None, None, None, None, None, 'r2(72,)', 'y2(61,)', 'r2(67,)', 'y2(51,)']
// Data values: [1, 0, 1, 0, None, None, None, None, None, None, None, None, 0, 0, 0, 4]
// Dest PEs: [42, 43, 50, 51, None, None, None, None, None, None, None, None, 2, 3, 10, 11]
9'd332: rdata =  56'b00000000000000000000000000000000000000000000000000001000;
//
// shift amount: 10, Lanes IDs: [2, 3]
9'd333: rdata =  56'b00000000000000000000000000000000000000100100000001011010;
//
// shift amount: 4, Lanes IDs: [10, 11]
9'd334: rdata =  56'b00000000000000100100000000000000000000000000000001010100;
//
// read [False, False, False, True]
// ['r2(107,)', 'y2(107,)', 'r2(106,)', 'y2(106,)', None, None, None, None, None, None, None, None, 'r2(83,)', 'y2(52,)', 'r2(71,)', 'y2(71,)']
// Data values: [1, 0, 1, 0, None, None, None, None, None, None, None, None, 0, 1, 1, 3]
// Dest PEs: [42, 43, 50, 51, None, None, None, None, None, None, None, None, 18, 19, 34, 35]
9'd335: rdata =  56'b00000000000000000000000000000000000000000000000000001000;
//
// shift amount: 10, Lanes IDs: [2, 3]
9'd336: rdata =  56'b00000000000000000000000000000000000001101100000001011010;
//
// shift amount: 12, Lanes IDs: [2, 3]
9'd337: rdata =  56'b00000000000000000000000000000000000010110100000001011100;
//
// read [False, False, False, True]
// ['r2(107,)', 'y2(107,)', 'r2(106,)', 'y2(106,)', None, None, None, None, None, None, None, None, 'r2(84,)', 'y2(84,)', 'r2(89,)', 'y2(89,)']
// Data values: [1, 0, 1, 0, None, None, None, None, None, None, None, None, 0, 4, 0, 4]
// Dest PEs: [42, 43, 50, 51, None, None, None, None, None, None, None, None, 42, 43, 50, 51]
9'd338: rdata =  56'b00000000000000000000000000000000000000000000000000001000;
//
// shift amount: 2, Lanes IDs: [10, 11]
9'd339: rdata =  56'b00000000000010110100000000000000000000000000000001010010;
//
// shift amount: 12, Lanes IDs: [2, 3]
9'd340: rdata =  56'b00000000000000000000000000000000000011111100000001011100;
//
// read [False, False, False, True]
// ['r2(107,)', 'y2(107,)', 'r2(106,)', 'y2(106,)', None, None, None, None, None, None, None, None, 'r2(100,)', 'y2(100,)', 'r2(81,)', 'y2(69,)']
// Data values: [1, 0, 1, 0, None, None, None, None, None, None, None, None, 1, 3, 0, 4]
// Dest PEs: [42, 43, 50, 51, None, None, None, None, None, None, None, None, 58, 59, 2, 3]
9'd341: rdata =  56'b00000000000000000000000000000000000000000000000000001000;
//
// shift amount: 2, Lanes IDs: [10, 11]
9'd342: rdata =  56'b00000000000011111100000000000000000000000000000001010010;
//
// shift amount: 12, Lanes IDs: [2, 3]
9'd343: rdata =  56'b00000000000000000000000000000000000000100100000001011100;
//
// read [False, False, False, True]
// ['r2(107,)', 'y2(107,)', 'r2(106,)', 'y2(106,)', None, None, None, None, None, None, None, None, 'r2(82,)', 'y2(62,)', 'r2(87,)', 'y2(58,)']
// Data values: [1, 0, 1, 0, None, None, None, None, None, None, None, None, 1, 2, 1, 5]
// Dest PEs: [42, 43, 50, 51, None, None, None, None, None, None, None, None, 10, 11, 18, 19]
9'd344: rdata =  56'b00000000000000000000000000000000000000000000000000001000;
//
// shift amount: 2, Lanes IDs: [10, 11]
9'd345: rdata =  56'b00000000000000100100000000000000000000000000000001010010;
//
// shift amount: 12, Lanes IDs: [2, 3]
9'd346: rdata =  56'b00000000000000000000000000000000000001101100000001011100;
//
// read [False, False, False, True]
// ['r2(107,)', 'y2(107,)', 'r2(106,)', 'y2(106,)', None, None, None, None, None, None, None, None, 'r2(79,)', 'y2(79,)', 'r2(95,)', 'y2(95,)']
// Data values: [1, 0, 1, 0, None, None, None, None, None, None, None, None, 0, 3, 1, 2]
// Dest PEs: [42, 43, 50, 51, None, None, None, None, None, None, None, None, 34, 35, 42, 43]
9'd347: rdata =  56'b00000000000000000000000000000000000000000000000000001000;
//
// shift amount: 10, Lanes IDs: [2, 3]
9'd348: rdata =  56'b00000000000000000000000000000000000010110100000001011010;
//
// shift amount: 4, Lanes IDs: [10, 11]
9'd349: rdata =  56'b00000000000010110100000000000000000000000000000001010100;
//
// read [False, False, False, True]
// ['r2(107,)', 'y2(107,)', 'r2(106,)', 'y2(106,)', None, None, None, None, None, None, None, None, 'r2(97,)', 'y2(97,)', 'r2(112,)', 'y2(112,)']
// Data values: [1, 0, 1, 0, None, None, None, None, None, None, None, None, 1, 0, 1, 1]
// Dest PEs: [42, 43, 50, 51, None, None, None, None, None, None, None, None, 50, 51, 58, 59]
9'd350: rdata =  56'b00000000000000000000000000000000000000000000000000001000;
//
// shift amount: 10, Lanes IDs: [2, 3]
9'd351: rdata =  56'b00000000000000000000000000000000000011111100000001011010;
//
// shift amount: 4, Lanes IDs: [10, 11]
9'd352: rdata =  56'b00000000000011111100000000000000000000000000000001010100;
//
// read [True, False, False, True]
// ['r2(107,)', 'y2(107,)', 'r2(106,)', 'y2(106,)', None, None, None, None, None, None, None, None, 'r2(90,)', 'y2(72,)', 'r2(92,)', 'y2(67,)']
// Data values: [1, 0, 1, 0, None, None, None, None, None, None, None, None, 1, 4, 0, 5]
// Dest PEs: [42, 43, 50, 51, None, None, None, None, None, None, None, None, 2, 3, 10, 11]
9'd353: rdata =  56'b00000000000000000000000000000000000000000000000000001001;
//
// shift amount: 0, Lanes IDs: [2, 3]
9'd354: rdata =  56'b00000000000000000000000000000000000011111100000001010000;
//
// shift amount: 10, Lanes IDs: [2, 3]
9'd355: rdata =  56'b00000000000000000000000000000000000000100100000001011010;
//
// shift amount: 4, Lanes IDs: [10, 11]
9'd356: rdata =  56'b00000000000000100100000000000000000000000000000001010100;
//
// shift amount: 6, Lanes IDs: [10, 11]
9'd357: rdata =  56'b00000000000010110100000000000000000000000000000001010110;
//
// read [True, False, False, True]
// ['r2(101,)', 'y2(81,)', 'r2(102,)', 'y2(82,)', None, None, None, None, None, None, None, None, 'r2(98,)', 'y2(70,)', 'r2(86,)', 'y2(86,)']
// Data values: [0, 4, 0, 1, None, None, None, None, None, None, None, None, 0, 5, 0, 0]
// Dest PEs: [2, 3, 10, 11, None, None, None, None, None, None, None, None, 18, 19, 34, 35]
9'd358: rdata =  56'b00000000000000000000000000000000000000000000000000001001;
//
// shift amount: 8, Lanes IDs: [10, 11]
9'd359: rdata =  56'b00000000000000100100000000000000000000000000000001011000;
//
// shift amount: 10, Lanes IDs: [2, 3]
9'd360: rdata =  56'b00000000000000000000000000000000000001101100000001011010;
//
// shift amount: 12, Lanes IDs: [2, 3]
9'd361: rdata =  56'b00000000000000000000000000000000000010110100000001011100;
//
// shift amount: 14, Lanes IDs: [2, 3]
9'd362: rdata =  56'b00000000000000000000000000000000000000100100000001011110;
//
// read [True, False, False, False]
// ['r2(109,)', 'y2(76,)', 'r2(91,)', 'y2(91,)', None, None, None, None, None, None, None, None, None, None, None, None]
// Data values: [0, 3, 0, 5, None, None, None, None, None, None, None, None, None, None, None, None]
// Dest PEs: [18, 19, 34, 35, None, None, None, None, None, None, None, None, None, None, None, None]
9'd363: rdata =  56'b00000000000000000000000000000000000000000000000000000001;
//
// shift amount: 0, Lanes IDs: [2, 3]
9'd364: rdata =  56'b00000000000000000000000000000000000010110100000001010000;
//
// shift amount: 14, Lanes IDs: [2, 3]
9'd365: rdata =  56'b00000000000000000000000000000000000001101100000001011110;
//
// read [True, False, False, False]
// ['r2(114,)', 'y2(114,)', 'r2(111,)', 'y2(111,)', None, None, None, None, None, None, None, None, None, None, None, None]
// Data values: [0, 1, 1, 4, None, None, None, None, None, None, None, None, None, None, None, None]
// Dest PEs: [42, 43, 50, 51, None, None, None, None, None, None, None, None, None, None, None, None]
9'd366: rdata =  56'b00000000000000000000000000000000000000000000000000000001;
//
// shift amount: 0, Lanes IDs: [2, 3]
9'd367: rdata =  56'b00000000000000000000000000000000000011111100000001010000;
//
// shift amount: 6, Lanes IDs: [10, 11]
9'd368: rdata =  56'b00000000000010110100000000000000000000000000000001010110;
//
// read [True, False, False, False]
// ['r2(113,)', 'y2(90,)', 'r2(116,)', 'y2(92,)', None, None, None, None, None, None, None, None, None, None, None, None]
// Data values: [1, 4, 0, 3, None, None, None, None, None, None, None, None, None, None, None, None]
// Dest PEs: [2, 3, 10, 11, None, None, None, None, None, None, None, None, None, None, None, None]
9'd369: rdata =  56'b00000000000000000000000000000000000000000000000000000001;
//
// shift amount: 8, Lanes IDs: [10, 11]
9'd370: rdata =  56'b00000000000000100100000000000000000000000000000001011000;
//
// shift amount: 14, Lanes IDs: [2, 3]
9'd371: rdata =  56'b00000000000000000000000000000000000000100100000001011110;
//
// read [True, False, False, False]
// ['r2(110,)', 'y2(77,)', 'r2(96,)', 'y2(96,)', None, None, None, None, None, None, None, None, None, None, None, None]
// Data values: [0, 2, 0, 5, None, None, None, None, None, None, None, None, None, None, None, None]
// Dest PEs: [18, 19, 34, 35, None, None, None, None, None, None, None, None, None, None, None, None]
9'd372: rdata =  56'b00000000000000000000000000000000000000000000000000000001;
//
// shift amount: 0, Lanes IDs: [2, 3]
9'd373: rdata =  56'b00000000000000000000000000000000000010110100000001010000;
//
// shift amount: 14, Lanes IDs: [2, 3]
9'd374: rdata =  56'b00000000000000000000000000000000000001101100000001011110;
//
// read [True, False, False, False]
// ['y2(113,)', 'y2(101,)', 'y2(102,)', 'r2(115,)', None, None, None, None, None, None, None, None, None, None, None, None]
// Data values: [0, 2, 0, 1, None, None, None, None, None, None, None, None, None, None, None, None]
// Dest PEs: [2, 3, 11, 18, None, None, None, None, None, None, None, None, None, None, None, None]
9'd375: rdata =  56'b00000000000000000000000000000000000000000000000000000001;
//
// shift amount: 1, Lanes IDs: [2]
9'd376: rdata =  56'b00000000000000000000000000000000000000001100000001010001;
//
// shift amount: 14, Lanes IDs: [2, 3]
9'd377: rdata =  56'b00000000000000000000000000000000000000100100000001011110;
//
// shift amount: 7, Lanes IDs: [11]
9'd378: rdata =  56'b00000000000000100000000000000000000000000000000001010111;
//
// read [True, False, False, False]
// ['y2(83,)', 'r2(103,)', 'y2(103,)', 'y2(116,)', None, None, None, None, None, None, None, None, None, None, None, None]
// Data values: [5, 1, 3, 5, None, None, None, None, None, None, None, None, None, None, None, None]
// Dest PEs: [19, 34, 35, 11, None, None, None, None, None, None, None, None, None, None, None, None]
9'd379: rdata =  56'b00000000000000000000000000000000000000000000000000000001;
//
// shift amount: 8, Lanes IDs: [11]
9'd380: rdata =  56'b00000000000000100000000000000000000000000000000001011000;
//
// shift amount: 13, Lanes IDs: [3]
9'd381: rdata =  56'b00000000000000000000000000000000000001100000000001011101;
//
// shift amount: 15, Lanes IDs: [2, 3]
9'd382: rdata =  56'b00000000000000000000000000000000000010110100000001011111;
//
// read [True, False, False, False]
// ['y1(33,)', 'y2(87,)', 'r2(104,)', 'y2(104,)', None, None, None, None, None, None, None, None, None, None, None, None]
// Data values: [2, 4, 0, 5, None, None, None, None, None, None, None, None, None, None, None, None]
// Dest PEs: [18, 19, 34, 35, None, None, None, None, None, None, None, None, None, None, None, None]
9'd383: rdata =  56'b00000000000000000000000000000000000000000000000000000001;
//
// shift amount: 0, Lanes IDs: [2, 3]
9'd384: rdata =  56'b00000000000000000000000000000000000010110100000001010000;
//
// shift amount: 14, Lanes IDs: [2, 3]
9'd385: rdata =  56'b00000000000000000000000000000000000001101100000001011110;
//
// read [True, False, False, False]
// ['y1(38,)', 'y2(98,)', 'y1(25,)', 'y1(51,)', None, None, None, None, None, None, None, None, None, None, None, None]
// Data values: [5, 1, 0, 4, None, None, None, None, None, None, None, None, None, None, None, None]
// Dest PEs: [18, 19, 34, 18, None, None, None, None, None, None, None, None, None, None, None, None]
9'd386: rdata =  56'b00000000000000000000000000000000000000000000000000000001;
//
// shift amount: 0, Lanes IDs: [2]
9'd387: rdata =  56'b00000000000000000000000000000000000000010100000001010000;
//
// shift amount: 14, Lanes IDs: [2, 3]
9'd388: rdata =  56'b00000000000000000000000000000000000001101100000001011110;
//
// shift amount: 1, Lanes IDs: [2]
9'd389: rdata =  56'b00000000000000000000000000000000000000001100000001010001;
//
// read [True, False, False, False]
// ['y2(109,)', 'y1(128,)', 'y2(110,)', 'y2(115,)', None, None, None, None, None, None, None, None, None, None, None, None]
// Data values: [2, 2, 2, 2, None, None, None, None, None, None, None, None, None, None, None, None]
// Dest PEs: [19, 18, 19, 19, None, None, None, None, None, None, None, None, None, None, None, None]
9'd390: rdata =  56'b00000000000000000000000000000000000000000000000000000001;
//
// shift amount: 13, Lanes IDs: [3]
9'd391: rdata =  56'b00000000000000000000000000000000000001100000000001011101;
//
// shift amount: 15, Lanes IDs: [2, 3]
9'd392: rdata =  56'b00000000000000000000000000000000000001101100000001011111;
//
// shift amount: 0, Lanes IDs: [3]
9'd393: rdata =  56'b00000000000000000000000000000000000001100000000001010000;
//
// wfi
9'd394: rdata =  56'b00000000000000000000000000000000000000000000000001100000;
//
// loop
9'd395: rdata =  56'b00000000000000000000000000000000000000000000000001110000;/****************************************************************************************/
default: rdata = 56'b00000000000000000000000000000000000000000000000001110000;

	endcase
	end

    //reg     [ADDR_WIDTH-1:0]        address;

// ******************************************************************
// Read Logic
// ******************************************************************

    always @ (posedge CLK)
    begin : READ_VALID
        if (RESET) begin
            DATA_OUT_VALID <= 1'b0;
        end else if (ENABLE) begin
            DATA_OUT_VALID <= 1'b1;
        end
    end



 always @(posedge CLK) begin
    if (ENABLE)
        DATA_OUT <= rdata;
end

endmodule
