
`timescale 1ns/1ps
module instruction_memory #(
    parameter integer addrLen = 5,
    parameter integer dataLen = 32,
    parameter integer peId  = 1
)(
    input clk,
    input rstn,
    
    input stall,
    input start,
    input restart,
    
    output reg [dataLen - 1: 0] data_out
);
//--------------------------------------------------------------------------------------
//reg [dataLen - 1: 0] mem  [0: (1 << addrLen) - 1];
reg [addrLen-1:0]        address;
reg enable;
reg [dataLen - 1: 0] rdata;
wire end_of_instruction;
always @(posedge clk or negedge rstn)
    if(~rstn)
        enable <= 1'b0;
    else if(start)
        enable <= 1'b1;
    else if(end_of_instruction)
       enable <= 1'b0;
always @(posedge clk or negedge rstn) begin
    if(~rstn)
        address <= {addrLen{1'b0}};
    else begin
        if(end_of_instruction)
            address <= {addrLen{1'b0}};
        else if(~stall && enable )
            address <= address + {{addrLen-1{1'b0}},1'b1};   
    end     
end
always @(posedge clk or negedge rstn) begin
    if(~rstn)
        data_out <= {1'b1,{dataLen-1{1'b0}}};
    else if((~stall && enable && ~end_of_instruction)||(end_of_instruction && start))
       data_out <= rdata;
end
    
assign end_of_instruction = (data_out[dataLen-1:dataLen-5] == 5'b0);
/****************************************************************************/
generate
if(peId == 0) begin
	always @(*) begin
		case(address)
			// PEs: 7 -> 8
			// srcs: (3, 0)(120) 2 --> (120) 2:PENB, pass, PUNB
			6'd0 : rdata = 41'b11000110111111100000000000000001000000000;
			// PEs: 56 -> 0
			// srcs: (8, 3)(146) 6 --> (146) 6:PUNB, pass, NI0
			6'd1 : rdata = 41'b11000110111111110000000000010000000000000;
			// PEs: 6 -> 16
			// srcs: (9, 1)(170) -3 --> (170) -3:PEGB6, pass, PUGB2
			6'd2 : rdata = 41'b11000111000011000000000000000000000001010;
			// PEs: 24 -> 1
			// srcs: (11, 2)(196) -1 --> (196) -1:PUGB3, pass, PENB
			6'd3 : rdata = 41'b11000111000001110000000000000000100000000;
			// PEs: 1 -> 48
			// srcs: (17, 5)(169) 13 --> (169) 13:PEGB1, pass, PUGB6
			6'd4 : rdata = 41'b11000111000000100000000000000000000001110;
			// PEs: 0 -> 1
			// srcs: (18, 4)(146) 6 --> (146) 6:NI0, pass, PENB
			6'd5 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 1 -> 8
			// srcs: (25, 6)(197) 5 --> (197) 5:PEGB1, pass, PUNB
			6'd6 : rdata = 41'b11000111000000100000000000000001000000000;
			// PEs: 40 -> 0
			// srcs: (30, 7)(211) 1 --> (211) 1:PUGB5, pass, NI0
			6'd7 : rdata = 41'b11000111000010110000000000010000000000000;
			// PEs: 56 -> 1
			// srcs: (41, 8)(216) 0 --> (216) 0:PUNB, pass, PENB
			6'd8 : rdata = 41'b11000110111111110000000000000000100000000;
			// PEs: 0 -> 1
			// srcs: (51, 9)(211) 1 --> (211) 1:NI0, pass, PENB
			6'd9 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 1 -> 24
			// srcs: (58, 10)(217) 1 --> (217) 1:PEGB1, pass, PUGB3
			6'd10 : rdata = 41'b11000111000000100000000000000000000001011;
			// PEs: 56 -> 1
			// srcs: (121, 11)(225) 0 --> (225) 0:PUNB, pass, PENB
			6'd11 : rdata = 41'b11000110111111110000000000000000100000000;
			// PEs: 56 -> 2
			// srcs: (125, 12)(225) 0 --> (225) 0:PUNB, pass, PEGB2
			6'd12 : rdata = 41'b11000110111111110000000000000000010100000;
			// PEs: 56 -> 3
			// srcs: (126, 13)(225) 0 --> (225) 0:PUNB, pass, PEGB3
			6'd13 : rdata = 41'b11000110111111110000000000000000010110000;
			// PEs: 56 -> 4
			// srcs: (127, 14)(225) 0 --> (225) 0:PUNB, pass, PEGB4
			6'd14 : rdata = 41'b11000110111111110000000000000000011000000;
			// PEs: 56 -> 5
			// srcs: (128, 15)(225) 0 --> (225) 0:PUNB, pass, PEGB5
			6'd15 : rdata = 41'b11000110111111110000000000000000011010000;
			// PEs: 56 -> 6
			// srcs: (129, 16)(225) 0 --> (225) 0:PUNB, pass, PEGB6
			6'd16 : rdata = 41'b11000110111111110000000000000000011100000;
			// PEs: 56 -> 7
			// srcs: (131, 17)(225) 0 --> (225) 0:PUNB, pass, PEGB7
			6'd17 : rdata = 41'b11000110111111110000000000000000011110000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 1) begin
	always @(*) begin
		case(address)
			// PEs: 1, 1 -> 2
			// srcs: (1, 0)(4) 2, (59) 2 --> (113) 4:ND0, NW0, *, PENB
			6'd0 : rdata = 41'b00011011000000000100000000000000100000000;
			// PEs: 4 -> 
			// srcs: (9, 1)(168) 9 --> (168) 9:PEGB4, pass, 
			6'd1 : rdata = 41'b11000111000010000000000000000000000000000;
			// PEs: 2, 1 -> 0
			// srcs: (12, 2)(167) 4, (168) 9 --> (169) 13:PEGB2, ALU, +, PEGB0
			6'd2 : rdata = 41'b00001111000001000011111111100000010000000;
			// PEs: 0 -> 
			// srcs: (13, 3)(196) -1 --> (196) -1:PENB, pass, 
			6'd3 : rdata = 41'b11000110111111100000000000000000000000000;
			// PEs: 1, 0 -> 0
			// srcs: (20, 4)(196) -1, (146) 6 --> (197) 5:ALU, PENB, +, PEGB0
			6'd4 : rdata = 41'b00001001111111111101111111000000010000000;
			// PEs: 0 -> 
			// srcs: (43, 5)(216) 0 --> (216) 0:PENB, pass, 
			6'd5 : rdata = 41'b11000110111111100000000000000000000000000;
			// PEs: 0, 1 -> 0
			// srcs: (53, 6)(211) 1, (216) 0 --> (217) 1:PENB, ALU, +, PEGB0
			6'd6 : rdata = 41'b00001110111111100011111111100000010000000;
			// PEs: 0, 1 -> 2
			// srcs: (124, 7)(225) 0, (4) 2 --> (226) 0:PENB, ND0, *, PENB
			6'd7 : rdata = 41'b00011110111111100110000000000000100000000;
			// PEs: 1, 2 -> 1
			// srcs: (133, 8)(59) 2, (280) 0 --> (334) 2:NW0, PEGB2, -, NW0
			6'd8 : rdata = 41'b00010010000000001110000010000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 2) begin
	always @(*) begin
		case(address)
			// PEs: 2, 2 -> 
			// srcs: (1, 0)(5) 2, (60) 0 --> (114) 0:ND0, NW0, *, 
			6'd0 : rdata = 41'b00011011000000000100000000000000000000000;
			// PEs: 1, 2 -> 1
			// srcs: (4, 1)(113) 4, (114) 0 --> (167) 4:PENB, ALU, +, PEGB1
			6'd1 : rdata = 41'b00001110111111100011111111100000010010000;
			// PEs: 2, 1 -> 1
			// srcs: (127, 3)(3) 1, (226) 0 --> (280) 0:NM0, PENB, *, PEGB1
			6'd2 : rdata = 41'b00011100000000001101111111000000010010000;
			// PEs: 0, 2 -> 3
			// srcs: (130, 2)(225) 0, (5) 2 --> (227) 0:PEGB0, ND0, *, PENB
			6'd3 : rdata = 41'b00011111000000000110000000000000100000000;
			// PEs: 2, 3 -> 2
			// srcs: (139, 4)(60) 0, (281) 0 --> (335) 0:NW0, PEGB3, -, NW0
			6'd4 : rdata = 41'b00010010000000001110000011000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 3) begin
	always @(*) begin
		case(address)
			// PEs: 3, 3 -> 4
			// srcs: (1, 0)(6) -2, (61) 0 --> (115) 0:ND0, NW0, *, PENB
			6'd0 : rdata = 41'b00011011000000000100000000000000100000000;
			// PEs: 0, 3 -> 3
			// srcs: (131, 1)(225) 0, (6) -2 --> (228) 0:PEGB0, ND0, *, NI0
			6'd1 : rdata = 41'b00011111000000000110000000010000000000000;
			// PEs: 3, 2 -> 2
			// srcs: (133, 2)(3) 1, (227) 0 --> (281) 0:NM0, PENB, *, PEGB2
			6'd2 : rdata = 41'b00011100000000001101111111000000010100000;
			// PEs: 3, 3 -> 
			// srcs: (134, 3)(3) 1, (228) 0 --> (282) 0:NM0, NI0, *, 
			6'd3 : rdata = 41'b00011100000000001010000000000000000000000;
			// PEs: 3, 3 -> 3
			// srcs: (137, 4)(61) 0, (282) 0 --> (336) 0:NW0, ALU, -, NW0
			6'd4 : rdata = 41'b00010010000000000011111111100100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 4) begin
	always @(*) begin
		case(address)
			// PEs: 4, 4 -> 
			// srcs: (1, 0)(7) -3, (62) -3 --> (116) 9:ND0, NW0, *, 
			6'd0 : rdata = 41'b00011011000000000100000000000000000000000;
			// PEs: 3, 4 -> 1
			// srcs: (4, 1)(115) 0, (116) 9 --> (168) 9:PENB, ALU, +, PEGB1
			6'd1 : rdata = 41'b00001110111111100011111111100000010010000;
			// PEs: 0, 4 -> 5
			// srcs: (132, 2)(225) 0, (7) -3 --> (229) 0:PEGB0, ND0, *, PENB
			6'd2 : rdata = 41'b00011111000000000110000000000000100000000;
			// PEs: 4, 5 -> 4
			// srcs: (141, 3)(62) -3, (283) 0 --> (337) -3:NW0, PEGB5, -, NW0
			6'd3 : rdata = 41'b00010010000000001110000101000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 5) begin
	always @(*) begin
		case(address)
			// PEs: 5, 5 -> 6
			// srcs: (1, 0)(8) 2, (63) -1 --> (117) -2:ND0, NW0, *, PENB
			6'd0 : rdata = 41'b00011011000000000100000000000000100000000;
			// PEs: 0, 5 -> 5
			// srcs: (133, 1)(225) 0, (8) 2 --> (230) 0:PEGB0, ND0, *, NI0
			6'd1 : rdata = 41'b00011111000000000110000000010000000000000;
			// PEs: 5, 4 -> 4
			// srcs: (135, 2)(3) 1, (229) 0 --> (283) 0:NM0, PENB, *, PEGB4
			6'd2 : rdata = 41'b00011100000000001101111111000000011000000;
			// PEs: 5, 5 -> 
			// srcs: (136, 3)(3) 1, (230) 0 --> (284) 0:NM0, NI0, *, 
			6'd3 : rdata = 41'b00011100000000001010000000000000000000000;
			// PEs: 5, 5 -> 5
			// srcs: (139, 4)(63) -1, (284) 0 --> (338) -1:NW0, ALU, -, NW0
			6'd4 : rdata = 41'b00010010000000000011111111100100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 6) begin
	always @(*) begin
		case(address)
			// PEs: 6, 6 -> 
			// srcs: (1, 0)(9) 1, (64) -1 --> (118) -1:ND0, NW0, *, 
			6'd0 : rdata = 41'b00011011000000000100000000000000000000000;
			// PEs: 5, 6 -> 0
			// srcs: (4, 1)(117) -2, (118) -1 --> (170) -3:PENB, ALU, +, PEGB0
			6'd1 : rdata = 41'b00001110111111100011111111100000010000000;
			// PEs: 0, 6 -> 7
			// srcs: (134, 2)(225) 0, (9) 1 --> (231) 0:PEGB0, ND0, *, PENB
			6'd2 : rdata = 41'b00011111000000000110000000000000100000000;
			// PEs: 6, 7 -> 6
			// srcs: (143, 3)(64) -1, (285) 0 --> (339) -1:NW0, PEGB7, -, NW0
			6'd3 : rdata = 41'b00010010000000001110000111000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 7) begin
	always @(*) begin
		case(address)
			// PEs: 7, 7 -> 0
			// srcs: (1, 0)(11) -1, (66) -2 --> (120) 2:ND0, NW0, *, PENB
			6'd0 : rdata = 41'b00011011000000000100000000000000100000000;
			// PEs: 0, 7 -> 7
			// srcs: (136, 1)(225) 0, (11) -1 --> (233) 0:PEGB0, ND0, *, NI0
			6'd1 : rdata = 41'b00011111000000000110000000010000000000000;
			// PEs: 7, 6 -> 6
			// srcs: (137, 2)(3) 1, (231) 0 --> (285) 0:NM0, PENB, *, PEGB6
			6'd2 : rdata = 41'b00011100000000001101111111000000011100000;
			// PEs: 7, 7 -> 
			// srcs: (139, 3)(3) 1, (233) 0 --> (287) 0:NM0, NI0, *, 
			6'd3 : rdata = 41'b00011100000000001010000000000000000000000;
			// PEs: 7, 7 -> 7
			// srcs: (142, 4)(66) -2, (287) 0 --> (341) -2:NW0, ALU, -, NW0
			6'd4 : rdata = 41'b00010010000000000011111111100100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 8) begin
	always @(*) begin
		case(address)
			// PEs: 0 -> 9
			// srcs: (5, 0)(120) 2 --> (120) 2:PUNB, pass, PENB
			6'd0 : rdata = 41'b11000110111111110000000000000000100000000;
			// PEs: 15 -> 16
			// srcs: (6, 2)(180) 2 --> (180) 2:PENB, pass, PUNB
			6'd1 : rdata = 41'b11000110111111100000000000000001000000000;
			// PEs: 13 -> 32
			// srcs: (9, 1)(176) -5 --> (176) -5:PEGB5, pass, PUGB4
			6'd2 : rdata = 41'b11000111000010100000000000000000000001100;
			// PEs: 32 -> 8
			// srcs: (14, 3)(202) -1 --> (202) -1:PUGB4, pass, NI0
			6'd3 : rdata = 41'b11000111000010010000000000010000000000000;
			// PEs: 56 -> 9
			// srcs: (15, 4)(153) 9 --> (153) 9:PUGB7, pass, PENB
			6'd4 : rdata = 41'b11000111000011110000000000000000100000000;
			// PEs: 10 -> 24
			// srcs: (19, 6)(175) 5 --> (175) 5:PEGB2, pass, PUGB3
			6'd5 : rdata = 41'b11000111000001000000000000000000000001011;
			// PEs: 8 -> 9
			// srcs: (21, 5)(202) -1 --> (202) -1:NI0, pass, PENB
			6'd6 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 24 -> 8
			// srcs: (22, 7)(195) 17 --> (195) 17:PUGB3, pass, NI0
			6'd7 : rdata = 41'b11000111000001110000000000010000000000000;
			// PEs: 0 -> 9
			// srcs: (27, 8)(197) 5 --> (197) 5:PUNB, pass, PENB
			6'd8 : rdata = 41'b11000110111111110000000000000000100000000;
			// PEs: 9 -> 16
			// srcs: (28, 10)(203) 8 --> (203) 8:PEGB1, pass, PUNB
			6'd9 : rdata = 41'b11000111000000100000000000000001000000000;
			// PEs: 8 -> 9
			// srcs: (37, 9)(195) 17 --> (195) 17:NI0, pass, PENB
			6'd10 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 9 -> 16
			// srcs: (44, 11)(198) 22 --> (198) 22:PEGB1, pass, PUNB
			6'd11 : rdata = 41'b11000111000000100000000000000001000000000;
			// PEs: 56 -> 9
			// srcs: (135, 12)(225) 0 --> (225) 0:PUGB7, pass, PENB
			6'd12 : rdata = 41'b11000111000011110000000000000000100000000;
			// PEs: 56 -> 10
			// srcs: (136, 13)(225) 0 --> (225) 0:PUGB7, pass, PEGB2
			6'd13 : rdata = 41'b11000111000011110000000000000000010100000;
			// PEs: 56 -> 11
			// srcs: (137, 14)(225) 0 --> (225) 0:PUGB7, pass, PEGB3
			6'd14 : rdata = 41'b11000111000011110000000000000000010110000;
			// PEs: 56 -> 12
			// srcs: (138, 15)(225) 0 --> (225) 0:PUGB7, pass, PEGB4
			6'd15 : rdata = 41'b11000111000011110000000000000000011000000;
			// PEs: 56 -> 13
			// srcs: (139, 16)(225) 0 --> (225) 0:PUGB7, pass, PEGB5
			6'd16 : rdata = 41'b11000111000011110000000000000000011010000;
			// PEs: 56 -> 14
			// srcs: (141, 17)(225) 0 --> (225) 0:PUGB7, pass, PEGB6
			6'd17 : rdata = 41'b11000111000011110000000000000000011100000;
			// PEs: 56 -> 15
			// srcs: (142, 18)(225) 0 --> (225) 0:PUGB7, pass, PEGB7
			6'd18 : rdata = 41'b11000111000011110000000000000000011110000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 9) begin
	always @(*) begin
		case(address)
			// PEs: 9, 9 -> 
			// srcs: (1, 0)(12) -2, (67) 0 --> (121) 0:ND0, NW0, *, 
			6'd0 : rdata = 41'b00011011000000000100000000000000000000000;
			// PEs: 8, 9 -> 10
			// srcs: (8, 1)(120) 2, (121) 0 --> (173) 2:PENB, ALU, +, PENB
			6'd1 : rdata = 41'b00001110111111100011111111100000100000000;
			// PEs: 8 -> 
			// srcs: (17, 2)(153) 9 --> (153) 9:PENB, pass, 
			6'd2 : rdata = 41'b11000110111111100000000000000000000000000;
			// PEs: 8, 9 -> 8
			// srcs: (23, 3)(202) -1, (153) 9 --> (203) 8:PENB, ALU, +, PEGB0
			6'd3 : rdata = 41'b00001110111111100011111111100000010000000;
			// PEs: 8 -> 
			// srcs: (29, 4)(197) 5 --> (197) 5:PENB, pass, 
			6'd4 : rdata = 41'b11000110111111100000000000000000000000000;
			// PEs: 8, 9 -> 8
			// srcs: (39, 5)(195) 17, (197) 5 --> (198) 22:PENB, ALU, +, PEGB0
			6'd5 : rdata = 41'b00001110111111100011111111100000010000000;
			// PEs: 8, 9 -> 10
			// srcs: (137, 6)(225) 0, (12) -2 --> (234) 0:PENB, ND0, *, PENB
			6'd6 : rdata = 41'b00011110111111100110000000000000100000000;
			// PEs: 9, 10 -> 9
			// srcs: (146, 7)(67) 0, (288) 0 --> (342) 0:NW0, PEGB2, -, NW0
			6'd7 : rdata = 41'b00010010000000001110000010000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 10) begin
	always @(*) begin
		case(address)
			// PEs: 10, 10 -> 11
			// srcs: (1, 0)(13) 2, (68) 1 --> (122) 2:ND0, NW0, *, PENB
			6'd0 : rdata = 41'b00011011000000000100000000000000100000000;
			// PEs: 9, 11 -> 8
			// srcs: (14, 1)(173) 2, (174) 3 --> (175) 5:PENB, PEGB3, +, PEGB0
			6'd1 : rdata = 41'b00001110111111101110000011000000010000000;
			// PEs: 10, 9 -> 9
			// srcs: (140, 3)(3) 1, (234) 0 --> (288) 0:NM0, PENB, *, PEGB1
			6'd2 : rdata = 41'b00011100000000001101111111000000010010000;
			// PEs: 8, 10 -> 11
			// srcs: (141, 2)(225) 0, (13) 2 --> (235) 0:PEGB0, ND0, *, PENB
			6'd3 : rdata = 41'b00011111000000000110000000000000100000000;
			// PEs: 10, 11 -> 10
			// srcs: (150, 4)(68) 1, (289) 0 --> (343) 1:NW0, PEGB3, -, NW0
			6'd4 : rdata = 41'b00010010000000001110000011000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 11) begin
	always @(*) begin
		case(address)
			// PEs: 11, 11 -> 
			// srcs: (1, 0)(14) 1, (69) 1 --> (123) 1:ND0, NW0, *, 
			6'd0 : rdata = 41'b00011011000000000100000000000000000000000;
			// PEs: 10, 11 -> 10
			// srcs: (4, 1)(122) 2, (123) 1 --> (174) 3:PENB, ALU, +, PEGB2
			6'd1 : rdata = 41'b00001110111111100011111111100000010100000;
			// PEs: 8, 11 -> 12
			// srcs: (142, 2)(225) 0, (14) 1 --> (236) 0:PEGB0, ND0, *, PENB
			6'd2 : rdata = 41'b00011111000000000110000000000000100000000;
			// PEs: 11, 10 -> 10
			// srcs: (144, 3)(3) 1, (235) 0 --> (289) 0:NM0, PENB, *, PEGB2
			6'd3 : rdata = 41'b00011100000000001101111111000000010100000;
			// PEs: 11, 12 -> 11
			// srcs: (151, 4)(69) 1, (290) 0 --> (344) 1:NW0, PEGB4, -, NW0
			6'd4 : rdata = 41'b00010010000000001110000100000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 12) begin
	always @(*) begin
		case(address)
			// PEs: 12, 12 -> 13
			// srcs: (1, 0)(15) -1, (70) 1 --> (124) -1:ND0, NW0, *, PENB
			6'd0 : rdata = 41'b00011011000000000100000000000000100000000;
			// PEs: 8, 12 -> 12
			// srcs: (143, 1)(225) 0, (15) -1 --> (237) 0:PEGB0, ND0, *, NI0
			6'd1 : rdata = 41'b00011111000000000110000000010000000000000;
			// PEs: 12, 11 -> 11
			// srcs: (145, 2)(3) 1, (236) 0 --> (290) 0:NM0, PENB, *, PEGB3
			6'd2 : rdata = 41'b00011100000000001101111111000000010110000;
			// PEs: 12, 12 -> 
			// srcs: (146, 3)(3) 1, (237) 0 --> (291) 0:NM0, NI0, *, 
			6'd3 : rdata = 41'b00011100000000001010000000000000000000000;
			// PEs: 12, 12 -> 12
			// srcs: (149, 4)(70) 1, (291) 0 --> (345) 1:NW0, ALU, -, NW0
			6'd4 : rdata = 41'b00010010000000000011111111100100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 13) begin
	always @(*) begin
		case(address)
			// PEs: 13, 13 -> 
			// srcs: (1, 0)(16) 2, (71) -2 --> (125) -4:ND0, NW0, *, 
			6'd0 : rdata = 41'b00011011000000000100000000000000000000000;
			// PEs: 12, 13 -> 8
			// srcs: (4, 1)(124) -1, (125) -4 --> (176) -5:PENB, ALU, +, PEGB0
			6'd1 : rdata = 41'b00001110111111100011111111100000010000000;
			// PEs: 8, 13 -> 14
			// srcs: (144, 2)(225) 0, (16) 2 --> (238) 0:PEGB0, ND0, *, PENB
			6'd2 : rdata = 41'b00011111000000000110000000000000100000000;
			// PEs: 13, 14 -> 13
			// srcs: (153, 3)(71) -2, (292) 0 --> (346) -2:NW0, PEGB6, -, NW0
			6'd3 : rdata = 41'b00010010000000001110000110000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 14) begin
	always @(*) begin
		case(address)
			// PEs: 14, 14 -> 15
			// srcs: (1, 0)(18) -1, (73) -2 --> (127) 2:ND0, NW0, *, PENB
			6'd0 : rdata = 41'b00011011000000000100000000000000100000000;
			// PEs: 8, 14 -> 14
			// srcs: (146, 1)(225) 0, (18) -1 --> (240) 0:PEGB0, ND0, *, NI0
			6'd1 : rdata = 41'b00011111000000000110000000010000000000000;
			// PEs: 14, 13 -> 13
			// srcs: (147, 2)(3) 1, (238) 0 --> (292) 0:NM0, PENB, *, PEGB5
			6'd2 : rdata = 41'b00011100000000001101111111000000011010000;
			// PEs: 14, 14 -> 
			// srcs: (149, 3)(3) 1, (240) 0 --> (294) 0:NM0, NI0, *, 
			6'd3 : rdata = 41'b00011100000000001010000000000000000000000;
			// PEs: 14, 14 -> 14
			// srcs: (152, 4)(73) -2, (294) 0 --> (348) -2:NW0, ALU, -, NW0
			6'd4 : rdata = 41'b00010010000000000011111111100100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 15) begin
	always @(*) begin
		case(address)
			// PEs: 15, 15 -> 
			// srcs: (1, 0)(19) -2, (74) 0 --> (128) 0:ND0, NW0, *, 
			6'd0 : rdata = 41'b00011011000000000100000000000000000000000;
			// PEs: 14, 15 -> 8
			// srcs: (4, 1)(127) 2, (128) 0 --> (180) 2:PENB, ALU, +, PENB
			6'd1 : rdata = 41'b00001110111111100011111111100000100000000;
			// PEs: 8, 15 -> 
			// srcs: (147, 2)(225) 0, (19) -2 --> (241) 0:PEGB0, ND0, *, 
			6'd2 : rdata = 41'b00011111000000000110000000000000000000000;
			// PEs: 15, 15 -> 
			// srcs: (150, 3)(3) 1, (241) 0 --> (295) 0:NM0, ALU, *, 
			6'd3 : rdata = 41'b00011100000000000011111111100000000000000;
			// PEs: 15, 15 -> 15
			// srcs: (153, 4)(74) 0, (295) 0 --> (349) 0:NW0, ALU, -, NW0
			6'd4 : rdata = 41'b00010010000000000011111111100100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 16) begin
	always @(*) begin
		case(address)
			// PEs: 23 -> 24
			// srcs: (3, 0)(137) 0 --> (137) 0:PENB, pass, PUNB
			6'd0 : rdata = 41'b11000110111111100000000000000001000000000;
			// PEs: 20 -> 48
			// srcs: (9, 5)(183) 9 --> (183) 9:PEGB4, pass, PUGB6
			6'd1 : rdata = 41'b11000111000010000000000000000000000001110;
			// PEs: 22 -> 56
			// srcs: (10, 6)(186) 5 --> (186) 5:PEGB6, pass, PUGB7
			6'd2 : rdata = 41'b11000111000011000000000000000000000001111;
			// PEs: 48 -> 16
			// srcs: (11, 2)(119) -2 --> (119) -2:PUGB6, pass, NI0
			6'd3 : rdata = 41'b11000111000011010000000000010000000000000;
			// PEs: 0 -> 17
			// srcs: (14, 1)(170) -3 --> (170) -3:PUGB0, pass, PENB
			6'd4 : rdata = 41'b11000111000000010000000000000000100000000;
			// PEs: 16 -> 17
			// srcs: (21, 3)(119) -2 --> (119) -2:NI0, pass, PENB
			6'd5 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 8 -> 17
			// srcs: (22, 4)(180) 2 --> (180) 2:PUNB, pass, PENB
			6'd6 : rdata = 41'b11000110111111110000000000000000100000000;
			// PEs: 32 -> 16
			// srcs: (23, 9)(201) 13 --> (201) 13:PUGB4, pass, NI0
			6'd7 : rdata = 41'b11000111000010010000000000010000000000000;
			// PEs: 17 -> 48
			// srcs: (28, 7)(171) -5 --> (171) -5:PEGB1, pass, PUGB6
			6'd8 : rdata = 41'b11000111000000100000000000000000000001110;
			// PEs: 17 -> 32
			// srcs: (29, 8)(182) 2 --> (182) 2:PEGB1, pass, PUGB4
			6'd9 : rdata = 41'b11000111000000100000000000000000000001100;
			// PEs: 8 -> 17
			// srcs: (30, 10)(203) 8 --> (203) 8:PUNB, pass, PENB
			6'd10 : rdata = 41'b11000110111111110000000000000000100000000;
			// PEs: 16 -> 17
			// srcs: (40, 11)(201) 13 --> (201) 13:NI0, pass, PENB
			6'd11 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 8 -> 17
			// srcs: (46, 12)(198) 22 --> (198) 22:PUNB, pass, PENB
			6'd12 : rdata = 41'b11000110111111110000000000000000100000000;
			// PEs: 17 -> 24
			// srcs: (57, 13)(205) 43 --> (205) 43:PEGB1, pass, PUNB
			6'd13 : rdata = 41'b11000111000000100000000000000001000000000;
			// PEs: 56 -> 17
			// srcs: (143, 14)(225) 0 --> (225) 0:PUGB7, pass, PENB
			6'd14 : rdata = 41'b11000111000011110000000000000000100000000;
			// PEs: 56 -> 18
			// srcs: (144, 15)(225) 0 --> (225) 0:PUGB7, pass, PEGB2
			6'd15 : rdata = 41'b11000111000011110000000000000000010100000;
			// PEs: 56 -> 19
			// srcs: (145, 16)(225) 0 --> (225) 0:PUGB7, pass, PEGB3
			6'd16 : rdata = 41'b11000111000011110000000000000000010110000;
			// PEs: 56 -> 20
			// srcs: (146, 17)(225) 0 --> (225) 0:PUGB7, pass, PEGB4
			6'd17 : rdata = 41'b11000111000011110000000000000000011000000;
			// PEs: 56 -> 21
			// srcs: (148, 18)(225) 0 --> (225) 0:PUGB7, pass, PEGB5
			6'd18 : rdata = 41'b11000111000011110000000000000000011010000;
			// PEs: 56 -> 22
			// srcs: (149, 19)(225) 0 --> (225) 0:PUGB7, pass, PEGB6
			6'd19 : rdata = 41'b11000111000011110000000000000000011100000;
			// PEs: 56 -> 23
			// srcs: (151, 20)(225) 0 --> (225) 0:PUGB7, pass, PEGB7
			6'd20 : rdata = 41'b11000111000011110000000000000000011110000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 17) begin
	always @(*) begin
		case(address)
			// PEs: 17, 17 -> 18
			// srcs: (1, 0)(20) -1, (75) 0 --> (129) 0:ND0, NW0, *, PENB
			6'd0 : rdata = 41'b00011011000000000100000000000000100000000;
			// PEs: 16 -> 
			// srcs: (16, 1)(170) -3 --> (170) -3:PENB, pass, 
			6'd1 : rdata = 41'b11000110111111100000000000000000000000000;
			// PEs: 17, 16 -> 16
			// srcs: (23, 2)(170) -3, (119) -2 --> (171) -5:ALU, PENB, +, PEGB0
			6'd2 : rdata = 41'b00001001111111111101111111000000010000000;
			// PEs: 16, 18 -> 16
			// srcs: (24, 3)(180) 2, (181) 0 --> (182) 2:PENB, PEGB2, +, PEGB0
			6'd3 : rdata = 41'b00001110111111101110000010000000010000000;
			// PEs: 16 -> 
			// srcs: (32, 4)(203) 8 --> (203) 8:PENB, pass, 
			6'd4 : rdata = 41'b11000110111111100000000000000000000000000;
			// PEs: 16, 17 -> 
			// srcs: (42, 5)(201) 13, (203) 8 --> (204) 21:PENB, ALU, +, 
			6'd5 : rdata = 41'b00001110111111100011111111100000000000000;
			// PEs: 16, 17 -> 16
			// srcs: (52, 6)(198) 22, (204) 21 --> (205) 43:PENB, ALU, +, PEGB0
			6'd6 : rdata = 41'b00001110111111100011111111100000010000000;
			// PEs: 16, 17 -> 18
			// srcs: (145, 7)(225) 0, (20) -1 --> (242) 0:PENB, ND0, *, PENB
			6'd7 : rdata = 41'b00011110111111100110000000000000100000000;
			// PEs: 17, 18 -> 17
			// srcs: (154, 8)(75) 0, (296) 0 --> (350) 0:NW0, PEGB2, -, NW0
			6'd8 : rdata = 41'b00010010000000001110000010000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 18) begin
	always @(*) begin
		case(address)
			// PEs: 18, 18 -> 
			// srcs: (1, 0)(21) -2, (76) 0 --> (130) 0:ND0, NW0, *, 
			6'd0 : rdata = 41'b00011011000000000100000000000000000000000;
			// PEs: 17, 18 -> 17
			// srcs: (4, 1)(129) 0, (130) 0 --> (181) 0:PENB, ALU, +, PEGB1
			6'd1 : rdata = 41'b00001110111111100011111111100000010010000;
			// PEs: 18, 17 -> 17
			// srcs: (148, 3)(3) 1, (242) 0 --> (296) 0:NM0, PENB, *, PEGB1
			6'd2 : rdata = 41'b00011100000000001101111111000000010010000;
			// PEs: 16, 18 -> 19
			// srcs: (149, 2)(225) 0, (21) -2 --> (243) 0:PEGB0, ND0, *, PENB
			6'd3 : rdata = 41'b00011111000000000110000000000000100000000;
			// PEs: 18, 19 -> 18
			// srcs: (158, 4)(76) 0, (297) 0 --> (351) 0:NW0, PEGB3, -, NW0
			6'd4 : rdata = 41'b00010010000000001110000011000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 19) begin
	always @(*) begin
		case(address)
			// PEs: 19, 19 -> 20
			// srcs: (1, 0)(22) -3, (77) -3 --> (131) 9:ND0, NW0, *, PENB
			6'd0 : rdata = 41'b00011011000000000100000000000000100000000;
			// PEs: 16, 19 -> 19
			// srcs: (150, 1)(225) 0, (22) -3 --> (244) 0:PEGB0, ND0, *, NI0
			6'd1 : rdata = 41'b00011111000000000110000000010000000000000;
			// PEs: 19, 18 -> 18
			// srcs: (152, 2)(3) 1, (243) 0 --> (297) 0:NM0, PENB, *, PEGB2
			6'd2 : rdata = 41'b00011100000000001101111111000000010100000;
			// PEs: 19, 19 -> 
			// srcs: (153, 3)(3) 1, (244) 0 --> (298) 0:NM0, NI0, *, 
			6'd3 : rdata = 41'b00011100000000001010000000000000000000000;
			// PEs: 19, 19 -> 19
			// srcs: (156, 4)(77) -3, (298) 0 --> (352) -3:NW0, ALU, -, NW0
			6'd4 : rdata = 41'b00010010000000000011111111100100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 20) begin
	always @(*) begin
		case(address)
			// PEs: 20, 20 -> 
			// srcs: (1, 0)(23) 0, (78) -3 --> (132) 0:ND0, NW0, *, 
			6'd0 : rdata = 41'b00011011000000000100000000000000000000000;
			// PEs: 19, 20 -> 16
			// srcs: (4, 1)(131) 9, (132) 0 --> (183) 9:PENB, ALU, +, PEGB0
			6'd1 : rdata = 41'b00001110111111100011111111100000010000000;
			// PEs: 16, 20 -> 21
			// srcs: (151, 2)(225) 0, (23) 0 --> (245) 0:PEGB0, ND0, *, PENB
			6'd2 : rdata = 41'b00011111000000000110000000000000100000000;
			// PEs: 20, 21 -> 20
			// srcs: (160, 3)(78) -3, (299) 0 --> (353) -3:NW0, PEGB5, -, NW0
			6'd3 : rdata = 41'b00010010000000001110000101000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 21) begin
	always @(*) begin
		case(address)
			// PEs: 21, 21 -> 22
			// srcs: (1, 0)(25) -3, (80) -3 --> (134) 9:ND0, NW0, *, PENB
			6'd0 : rdata = 41'b00011011000000000100000000000000100000000;
			// PEs: 16, 21 -> 21
			// srcs: (153, 1)(225) 0, (25) -3 --> (247) 0:PEGB0, ND0, *, NI0
			6'd1 : rdata = 41'b00011111000000000110000000010000000000000;
			// PEs: 21, 20 -> 20
			// srcs: (154, 2)(3) 1, (245) 0 --> (299) 0:NM0, PENB, *, PEGB4
			6'd2 : rdata = 41'b00011100000000001101111111000000011000000;
			// PEs: 21, 21 -> 
			// srcs: (156, 3)(3) 1, (247) 0 --> (301) 0:NM0, NI0, *, 
			6'd3 : rdata = 41'b00011100000000001010000000000000000000000;
			// PEs: 21, 21 -> 21
			// srcs: (159, 4)(80) -3, (301) 0 --> (355) -3:NW0, ALU, -, NW0
			6'd4 : rdata = 41'b00010010000000000011111111100100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 22) begin
	always @(*) begin
		case(address)
			// PEs: 22, 22 -> 
			// srcs: (1, 0)(26) 2, (81) -2 --> (135) -4:ND0, NW0, *, 
			6'd0 : rdata = 41'b00011011000000000100000000000000000000000;
			// PEs: 21, 22 -> 16
			// srcs: (4, 1)(134) 9, (135) -4 --> (186) 5:PENB, ALU, +, PEGB0
			6'd1 : rdata = 41'b00001110111111100011111111100000010000000;
			// PEs: 16, 22 -> 23
			// srcs: (154, 2)(225) 0, (26) 2 --> (248) 0:PEGB0, ND0, *, PENB
			6'd2 : rdata = 41'b00011111000000000110000000000000100000000;
			// PEs: 22, 23 -> 22
			// srcs: (163, 3)(81) -2, (302) 0 --> (356) -2:NW0, PEGB7, -, NW0
			6'd3 : rdata = 41'b00010010000000001110000111000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 23) begin
	always @(*) begin
		case(address)
			// PEs: 23, 23 -> 16
			// srcs: (1, 0)(28) -3, (83) 0 --> (137) 0:ND0, NW0, *, PENB
			6'd0 : rdata = 41'b00011011000000000100000000000000100000000;
			// PEs: 16, 23 -> 23
			// srcs: (156, 1)(225) 0, (28) -3 --> (250) 0:PEGB0, ND0, *, NI0
			6'd1 : rdata = 41'b00011111000000000110000000010000000000000;
			// PEs: 23, 22 -> 22
			// srcs: (157, 2)(3) 1, (248) 0 --> (302) 0:NM0, PENB, *, PEGB6
			6'd2 : rdata = 41'b00011100000000001101111111000000011100000;
			// PEs: 23, 23 -> 
			// srcs: (159, 3)(3) 1, (250) 0 --> (304) 0:NM0, NI0, *, 
			6'd3 : rdata = 41'b00011100000000001010000000000000000000000;
			// PEs: 23, 23 -> 23
			// srcs: (162, 4)(83) 0, (304) 0 --> (358) 0:NW0, ALU, -, NW0
			6'd4 : rdata = 41'b00010010000000000011111111100100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 24) begin
	always @(*) begin
		case(address)
			// PEs: 16 -> 25
			// srcs: (5, 0)(137) 0 --> (137) 0:PUNB, pass, PENB
			6'd0 : rdata = 41'b11000110111111110000000000000000100000000;
			// PEs: 31 -> 0
			// srcs: (6, 2)(196) -1 --> (196) -1:PENB, pass, PUGB0
			6'd1 : rdata = 41'b11000110111111100000000000000000000001000;
			// PEs: 48 -> 25
			// srcs: (8, 1)(139) 0 --> (139) 0:PUGB6, pass, PENB
			6'd2 : rdata = 41'b11000111000011010000000000000000100000000;
			// PEs: 26 -> 8
			// srcs: (17, 7)(195) 17 --> (195) 17:PEGB2, pass, PUGB1
			6'd3 : rdata = 41'b11000111000001000000000000000000000001001;
			// PEs: 25 -> 40
			// srcs: (23, 6)(189) 2 --> (189) 2:PEGB1, pass, PUGB5
			6'd4 : rdata = 41'b11000111000000100000000000000000000001101;
			// PEs: 8 -> 24
			// srcs: (24, 3)(175) 5 --> (175) 5:PUGB1, pass, NI0
			6'd5 : rdata = 41'b11000111000000110000000000010000000000000;
			// PEs: 32 -> 25
			// srcs: (33, 4)(177) -1 --> (177) -1:PUGB4, pass, PENB
			6'd6 : rdata = 41'b11000111000010010000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (40, 5)(175) 5 --> (175) 5:NI0, pass, PENB
			6'd7 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 25 -> 48
			// srcs: (47, 8)(178) 4 --> (178) 4:PEGB1, pass, PUGB6
			6'd8 : rdata = 41'b11000111000000100000000000000000000001110;
			// PEs: 16 -> 24
			// srcs: (59, 9)(205) 43 --> (205) 43:PUNB, pass, NI0
			6'd9 : rdata = 41'b11000110111111110000000000010000000000000;
			// PEs: 0 -> 25
			// srcs: (63, 10)(217) 1 --> (217) 1:PUGB0, pass, PENB
			6'd10 : rdata = 41'b11000111000000010000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (70, 11)(205) 43 --> (205) 43:NI0, pass, PENB
			6'd11 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 25 -> 32
			// srcs: (77, 12)(218) 44 --> (218) 44:PEGB1, pass, PUNB
			6'd12 : rdata = 41'b11000111000000100000000000000001000000000;
			// PEs: 56 -> 25
			// srcs: (152, 13)(225) 0 --> (225) 0:PUGB7, pass, PENB
			6'd13 : rdata = 41'b11000111000011110000000000000000100000000;
			// PEs: 56 -> 26
			// srcs: (154, 14)(225) 0 --> (225) 0:PUGB7, pass, PEGB2
			6'd14 : rdata = 41'b11000111000011110000000000000000010100000;
			// PEs: 56 -> 27
			// srcs: (155, 15)(225) 0 --> (225) 0:PUGB7, pass, PEGB3
			6'd15 : rdata = 41'b11000111000011110000000000000000010110000;
			// PEs: 56 -> 28
			// srcs: (156, 16)(225) 0 --> (225) 0:PUGB7, pass, PEGB4
			6'd16 : rdata = 41'b11000111000011110000000000000000011000000;
			// PEs: 56 -> 29
			// srcs: (157, 17)(225) 0 --> (225) 0:PUGB7, pass, PEGB5
			6'd17 : rdata = 41'b11000111000011110000000000000000011010000;
			// PEs: 56 -> 30
			// srcs: (158, 18)(225) 0 --> (225) 0:PUGB7, pass, PEGB6
			6'd18 : rdata = 41'b11000111000011110000000000000000011100000;
			// PEs: 56 -> 31
			// srcs: (159, 19)(225) 0 --> (225) 0:PUGB7, pass, PEGB7
			6'd19 : rdata = 41'b11000111000011110000000000000000011110000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 25) begin
	always @(*) begin
		case(address)
			// PEs: 25, 25 -> 
			// srcs: (1, 0)(29) -2, (84) -1 --> (138) 2:ND0, NW0, *, 
			6'd0 : rdata = 41'b00011011000000000100000000000000000000000;
			// PEs: 24, 25 -> 
			// srcs: (8, 1)(137) 0, (138) 2 --> (188) 2:PENB, ALU, +, 
			6'd1 : rdata = 41'b00001110111111100011111111100000000000000;
			// PEs: 25, 24 -> 24
			// srcs: (18, 2)(188) 2, (139) 0 --> (189) 2:ALU, PENB, +, PEGB0
			6'd2 : rdata = 41'b00001001111111111101111111000000010000000;
			// PEs: 24 -> 
			// srcs: (35, 3)(177) -1 --> (177) -1:PENB, pass, 
			6'd3 : rdata = 41'b11000110111111100000000000000000000000000;
			// PEs: 24, 25 -> 24
			// srcs: (42, 4)(175) 5, (177) -1 --> (178) 4:PENB, ALU, +, PEGB0
			6'd4 : rdata = 41'b00001110111111100011111111100000010000000;
			// PEs: 24 -> 
			// srcs: (65, 5)(217) 1 --> (217) 1:PENB, pass, 
			6'd5 : rdata = 41'b11000110111111100000000000000000000000000;
			// PEs: 24, 25 -> 24
			// srcs: (72, 6)(205) 43, (217) 1 --> (218) 44:PENB, ALU, +, PEGB0
			6'd6 : rdata = 41'b00001110111111100011111111100000010000000;
			// PEs: 24, 25 -> 26
			// srcs: (154, 7)(225) 0, (29) -2 --> (251) 0:PENB, ND0, *, PENB
			6'd7 : rdata = 41'b00011110111111100110000000000000100000000;
			// PEs: 25, 26 -> 25
			// srcs: (163, 8)(84) -1, (305) 0 --> (359) -1:NW0, PEGB2, -, NW0
			6'd8 : rdata = 41'b00010010000000001110000010000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 26) begin
	always @(*) begin
		case(address)
			// PEs: 26, 26 -> 27
			// srcs: (1, 0)(31) 1, (86) 1 --> (140) 1:ND0, NW0, *, PENB
			6'd0 : rdata = 41'b00011011000000000100000000000000100000000;
			// PEs: 29 -> 
			// srcs: (9, 1)(194) 10 --> (194) 10:PEGB5, pass, 
			6'd1 : rdata = 41'b11000111000010100000000000000000000000000;
			// PEs: 27, 26 -> 24
			// srcs: (12, 2)(193) 7, (194) 10 --> (195) 17:PEGB3, ALU, +, PEGB0
			6'd2 : rdata = 41'b00001111000001100011111111100000010000000;
			// PEs: 26, 25 -> 25
			// srcs: (157, 4)(3) 1, (251) 0 --> (305) 0:NM0, PENB, *, PEGB1
			6'd3 : rdata = 41'b00011100000000001101111111000000010010000;
			// PEs: 24, 26 -> 27
			// srcs: (159, 3)(225) 0, (31) 1 --> (253) 0:PEGB0, ND0, *, PENB
			6'd4 : rdata = 41'b00011111000000000110000000000000100000000;
			// PEs: 26, 27 -> 26
			// srcs: (168, 5)(86) 1, (307) 0 --> (361) 1:NW0, PEGB3, -, NW0
			6'd5 : rdata = 41'b00010010000000001110000011000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 27) begin
	always @(*) begin
		case(address)
			// PEs: 27, 27 -> 
			// srcs: (1, 0)(32) -3, (87) -2 --> (141) 6:ND0, NW0, *, 
			6'd0 : rdata = 41'b00011011000000000100000000000000000000000;
			// PEs: 26, 27 -> 26
			// srcs: (4, 1)(140) 1, (141) 6 --> (193) 7:PENB, ALU, +, PEGB2
			6'd1 : rdata = 41'b00001110111111100011111111100000010100000;
			// PEs: 24, 27 -> 28
			// srcs: (160, 2)(225) 0, (32) -3 --> (254) 0:PEGB0, ND0, *, PENB
			6'd2 : rdata = 41'b00011111000000000110000000000000100000000;
			// PEs: 27, 26 -> 26
			// srcs: (162, 3)(3) 1, (253) 0 --> (307) 0:NM0, PENB, *, PEGB2
			6'd3 : rdata = 41'b00011100000000001101111111000000010100000;
			// PEs: 27, 28 -> 27
			// srcs: (169, 4)(87) -2, (308) 0 --> (362) -2:NW0, PEGB4, -, NW0
			6'd4 : rdata = 41'b00010010000000001110000100000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 28) begin
	always @(*) begin
		case(address)
			// PEs: 28, 28 -> 29
			// srcs: (1, 0)(33) -3, (88) -2 --> (142) 6:ND0, NW0, *, PENB
			6'd0 : rdata = 41'b00011011000000000100000000000000100000000;
			// PEs: 24, 28 -> 28
			// srcs: (161, 1)(225) 0, (33) -3 --> (255) 0:PEGB0, ND0, *, NI0
			6'd1 : rdata = 41'b00011111000000000110000000010000000000000;
			// PEs: 28, 27 -> 27
			// srcs: (163, 2)(3) 1, (254) 0 --> (308) 0:NM0, PENB, *, PEGB3
			6'd2 : rdata = 41'b00011100000000001101111111000000010110000;
			// PEs: 28, 28 -> 
			// srcs: (164, 3)(3) 1, (255) 0 --> (309) 0:NM0, NI0, *, 
			6'd3 : rdata = 41'b00011100000000001010000000000000000000000;
			// PEs: 28, 28 -> 28
			// srcs: (167, 4)(88) -2, (309) 0 --> (363) -2:NW0, ALU, -, NW0
			6'd4 : rdata = 41'b00010010000000000011111111100100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 29) begin
	always @(*) begin
		case(address)
			// PEs: 29, 29 -> 
			// srcs: (1, 0)(34) 2, (89) 2 --> (143) 4:ND0, NW0, *, 
			6'd0 : rdata = 41'b00011011000000000100000000000000000000000;
			// PEs: 28, 29 -> 26
			// srcs: (4, 1)(142) 6, (143) 4 --> (194) 10:PENB, ALU, +, PEGB2
			6'd1 : rdata = 41'b00001110111111100011111111100000010100000;
			// PEs: 24, 29 -> 30
			// srcs: (162, 2)(225) 0, (34) 2 --> (256) 0:PEGB0, ND0, *, PENB
			6'd2 : rdata = 41'b00011111000000000110000000000000100000000;
			// PEs: 29, 30 -> 29
			// srcs: (171, 3)(89) 2, (310) 0 --> (364) 2:NW0, PEGB6, -, NW0
			6'd3 : rdata = 41'b00010010000000001110000110000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 30) begin
	always @(*) begin
		case(address)
			// PEs: 30, 30 -> 31
			// srcs: (1, 0)(35) -1, (90) 1 --> (144) -1:ND0, NW0, *, PENB
			6'd0 : rdata = 41'b00011011000000000100000000000000100000000;
			// PEs: 24, 30 -> 30
			// srcs: (163, 1)(225) 0, (35) -1 --> (257) 0:PEGB0, ND0, *, NI0
			6'd1 : rdata = 41'b00011111000000000110000000010000000000000;
			// PEs: 30, 29 -> 29
			// srcs: (165, 2)(3) 1, (256) 0 --> (310) 0:NM0, PENB, *, PEGB5
			6'd2 : rdata = 41'b00011100000000001101111111000000011010000;
			// PEs: 30, 30 -> 
			// srcs: (166, 3)(3) 1, (257) 0 --> (311) 0:NM0, NI0, *, 
			6'd3 : rdata = 41'b00011100000000001010000000000000000000000;
			// PEs: 30, 30 -> 30
			// srcs: (169, 4)(90) 1, (311) 0 --> (365) 1:NW0, ALU, -, NW0
			6'd4 : rdata = 41'b00010010000000000011111111100100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 31) begin
	always @(*) begin
		case(address)
			// PEs: 31, 31 -> 
			// srcs: (1, 0)(36) 0, (91) -1 --> (145) 0:ND0, NW0, *, 
			6'd0 : rdata = 41'b00011011000000000100000000000000000000000;
			// PEs: 30, 31 -> 24
			// srcs: (4, 1)(144) -1, (145) 0 --> (196) -1:PENB, ALU, +, PENB
			6'd1 : rdata = 41'b00001110111111100011111111100000100000000;
			// PEs: 24, 31 -> 
			// srcs: (164, 2)(225) 0, (36) 0 --> (258) 0:PEGB0, ND0, *, 
			6'd2 : rdata = 41'b00011111000000000110000000000000000000000;
			// PEs: 31, 31 -> 
			// srcs: (167, 3)(3) 1, (258) 0 --> (312) 0:NM0, ALU, *, 
			6'd3 : rdata = 41'b00011100000000000011111111100000000000000;
			// PEs: 31, 31 -> 31
			// srcs: (170, 4)(91) -1, (312) 0 --> (366) -1:NW0, ALU, -, NW0
			6'd4 : rdata = 41'b00010010000000000011111111100100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 32) begin
	always @(*) begin
		case(address)
			// PEs: 39 -> 40
			// srcs: (3, 0)(154) -2 --> (154) -2:PENB, pass, PUNB
			6'd0 : rdata = 41'b11000110111111100000000000000001000000000;
			// PEs: 38 -> 8
			// srcs: (9, 4)(202) -1 --> (202) -1:PEGB6, pass, PUGB1
			6'd1 : rdata = 41'b11000111000011000000000000000000000001001;
			// PEs: 48 -> 32
			// srcs: (12, 2)(126) 4 --> (126) 4:PUGB6, pass, NI0
			6'd2 : rdata = 41'b11000111000011010000000000010000000000000;
			// PEs: 8 -> 33
			// srcs: (14, 1)(176) -5 --> (176) -5:PUGB1, pass, PENB
			6'd3 : rdata = 41'b11000111000000110000000000000000100000000;
			// PEs: 35 -> 16
			// srcs: (15, 9)(201) 13 --> (201) 13:PEGB3, pass, PUGB2
			6'd4 : rdata = 41'b11000111000001100000000000000000000001010;
			// PEs: 32 -> 33
			// srcs: (21, 3)(126) 4 --> (126) 4:NI0, pass, PENB
			6'd5 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 33 -> 24
			// srcs: (28, 5)(177) -1 --> (177) -1:PEGB1, pass, PUGB3
			6'd6 : rdata = 41'b11000111000000100000000000000000000001011;
			// PEs: 16 -> 32
			// srcs: (34, 6)(182) 2 --> (182) 2:PUGB2, pass, NI0
			6'd7 : rdata = 41'b11000111000001010000000000010000000000000;
			// PEs: 48 -> 33
			// srcs: (35, 7)(184) 7 --> (184) 7:PUGB6, pass, PENB
			6'd8 : rdata = 41'b11000111000011010000000000000000100000000;
			// PEs: 32 -> 33
			// srcs: (41, 8)(182) 2 --> (182) 2:NI0, pass, PENB
			6'd9 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 33 -> 40
			// srcs: (48, 10)(185) 9 --> (185) 9:PEGB1, pass, PUNB
			6'd10 : rdata = 41'b11000111000000100000000000000001000000000;
			// PEs: 48 -> 32
			// srcs: (75, 11)(192) 32 --> (192) 32:PUGB6, pass, NI0
			6'd11 : rdata = 41'b11000111000011010000000000010000000000000;
			// PEs: 24 -> 33
			// srcs: (79, 12)(218) 44 --> (218) 44:PUNB, pass, PENB
			6'd12 : rdata = 41'b11000110111111110000000000000000100000000;
			// PEs: 32 -> 33
			// srcs: (89, 13)(192) 32 --> (192) 32:NI0, pass, PENB
			6'd13 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 33 -> 56
			// srcs: (96, 14)(219) 76 --> (219) 76:PEGB1, pass, PUGB7
			6'd14 : rdata = 41'b11000111000000100000000000000000000001111;
			// PEs: 56 -> 33
			// srcs: (160, 15)(225) 0 --> (225) 0:PUGB7, pass, PENB
			6'd15 : rdata = 41'b11000111000011110000000000000000100000000;
			// PEs: 56 -> 34
			// srcs: (161, 16)(225) 0 --> (225) 0:PUGB7, pass, PEGB2
			6'd16 : rdata = 41'b11000111000011110000000000000000010100000;
			// PEs: 56 -> 35
			// srcs: (162, 17)(225) 0 --> (225) 0:PUGB7, pass, PEGB3
			6'd17 : rdata = 41'b11000111000011110000000000000000010110000;
			// PEs: 56 -> 36
			// srcs: (163, 18)(225) 0 --> (225) 0:PUGB7, pass, PEGB4
			6'd18 : rdata = 41'b11000111000011110000000000000000011000000;
			// PEs: 56 -> 37
			// srcs: (164, 19)(225) 0 --> (225) 0:PUGB7, pass, PEGB5
			6'd19 : rdata = 41'b11000111000011110000000000000000011010000;
			// PEs: 56 -> 38
			// srcs: (165, 20)(225) 0 --> (225) 0:PUGB7, pass, PEGB6
			6'd20 : rdata = 41'b11000111000011110000000000000000011100000;
			// PEs: 56 -> 39
			// srcs: (167, 21)(225) 0 --> (225) 0:PUGB7, pass, PEGB7
			6'd21 : rdata = 41'b11000111000011110000000000000000011110000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 33) begin
	always @(*) begin
		case(address)
			// PEs: 33, 33 -> 34
			// srcs: (1, 0)(38) 2, (93) 2 --> (147) 4:ND0, NW0, *, PENB
			6'd0 : rdata = 41'b00011011000000000100000000000000100000000;
			// PEs: 32 -> 
			// srcs: (16, 1)(176) -5 --> (176) -5:PENB, pass, 
			6'd1 : rdata = 41'b11000110111111100000000000000000000000000;
			// PEs: 33, 32 -> 32
			// srcs: (23, 2)(176) -5, (126) 4 --> (177) -1:ALU, PENB, +, PEGB0
			6'd2 : rdata = 41'b00001001111111111101111111000000010000000;
			// PEs: 32 -> 
			// srcs: (37, 3)(184) 7 --> (184) 7:PENB, pass, 
			6'd3 : rdata = 41'b11000110111111100000000000000000000000000;
			// PEs: 32, 33 -> 32
			// srcs: (43, 4)(182) 2, (184) 7 --> (185) 9:PENB, ALU, +, PEGB0
			6'd4 : rdata = 41'b00001110111111100011111111100000010000000;
			// PEs: 32 -> 
			// srcs: (81, 5)(218) 44 --> (218) 44:PENB, pass, 
			6'd5 : rdata = 41'b11000110111111100000000000000000000000000;
			// PEs: 32, 33 -> 32
			// srcs: (91, 6)(192) 32, (218) 44 --> (219) 76:PENB, ALU, +, PEGB0
			6'd6 : rdata = 41'b00001110111111100011111111100000010000000;
			// PEs: 32, 33 -> 34
			// srcs: (162, 7)(225) 0, (38) 2 --> (260) 0:PENB, ND0, *, PENB
			6'd7 : rdata = 41'b00011110111111100110000000000000100000000;
			// PEs: 33, 34 -> 33
			// srcs: (171, 8)(93) 2, (314) 0 --> (368) 2:NW0, PEGB2, -, NW0
			6'd8 : rdata = 41'b00010010000000001110000010000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 34) begin
	always @(*) begin
		case(address)
			// PEs: 34, 34 -> 
			// srcs: (1, 0)(39) -3, (94) -1 --> (148) 3:ND0, NW0, *, 
			6'd0 : rdata = 41'b00011011000000000100000000000000000000000;
			// PEs: 33, 34 -> 35
			// srcs: (4, 1)(147) 4, (148) 3 --> (199) 7:PENB, ALU, +, PENB
			6'd1 : rdata = 41'b00001110111111100011111111100000100000000;
			// PEs: 34, 33 -> 33
			// srcs: (165, 3)(3) 1, (260) 0 --> (314) 0:NM0, PENB, *, PEGB1
			6'd2 : rdata = 41'b00011100000000001101111111000000010010000;
			// PEs: 32, 34 -> 35
			// srcs: (166, 2)(225) 0, (39) -3 --> (261) 0:PEGB0, ND0, *, PENB
			6'd3 : rdata = 41'b00011111000000000110000000000000100000000;
			// PEs: 34, 35 -> 34
			// srcs: (175, 4)(94) -1, (315) 0 --> (369) -1:NW0, PEGB3, -, NW0
			6'd4 : rdata = 41'b00010010000000001110000011000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 35) begin
	always @(*) begin
		case(address)
			// PEs: 35, 35 -> 36
			// srcs: (1, 0)(40) -3, (95) -2 --> (149) 6:ND0, NW0, *, PENB
			6'd0 : rdata = 41'b00011011000000000100000000000000100000000;
			// PEs: 34, 36 -> 32
			// srcs: (10, 1)(199) 7, (200) 6 --> (201) 13:PENB, PEGB4, +, PEGB0
			6'd1 : rdata = 41'b00001110111111101110000100000000010000000;
			// PEs: 32, 35 -> 36
			// srcs: (167, 2)(225) 0, (40) -3 --> (262) 0:PEGB0, ND0, *, PENB
			6'd2 : rdata = 41'b00011111000000000110000000000000100000000;
			// PEs: 35, 34 -> 34
			// srcs: (169, 3)(3) 1, (261) 0 --> (315) 0:NM0, PENB, *, PEGB2
			6'd3 : rdata = 41'b00011100000000001101111111000000010100000;
			// PEs: 35, 36 -> 35
			// srcs: (176, 4)(95) -2, (316) 0 --> (370) -2:NW0, PEGB4, -, NW0
			6'd4 : rdata = 41'b00010010000000001110000100000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 36) begin
	always @(*) begin
		case(address)
			// PEs: 36, 36 -> 
			// srcs: (1, 0)(41) -3, (96) 0 --> (150) 0:ND0, NW0, *, 
			6'd0 : rdata = 41'b00011011000000000100000000000000000000000;
			// PEs: 35, 36 -> 35
			// srcs: (4, 1)(149) 6, (150) 0 --> (200) 6:PENB, ALU, +, PEGB3
			6'd1 : rdata = 41'b00001110111111100011111111100000010110000;
			// PEs: 32, 36 -> 37
			// srcs: (168, 2)(225) 0, (41) -3 --> (263) 0:PEGB0, ND0, *, PENB
			6'd2 : rdata = 41'b00011111000000000110000000000000100000000;
			// PEs: 36, 35 -> 35
			// srcs: (170, 3)(3) 1, (262) 0 --> (316) 0:NM0, PENB, *, PEGB3
			6'd3 : rdata = 41'b00011100000000001101111111000000010110000;
			// PEs: 36, 37 -> 36
			// srcs: (177, 4)(96) 0, (317) 0 --> (371) 0:NW0, PEGB5, -, NW0
			6'd4 : rdata = 41'b00010010000000001110000101000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 37) begin
	always @(*) begin
		case(address)
			// PEs: 37, 37 -> 38
			// srcs: (1, 0)(42) 0, (97) 2 --> (151) 0:ND0, NW0, *, PENB
			6'd0 : rdata = 41'b00011011000000000100000000000000100000000;
			// PEs: 32, 37 -> 37
			// srcs: (169, 1)(225) 0, (42) 0 --> (264) 0:PEGB0, ND0, *, NI0
			6'd1 : rdata = 41'b00011111000000000110000000010000000000000;
			// PEs: 37, 36 -> 36
			// srcs: (171, 2)(3) 1, (263) 0 --> (317) 0:NM0, PENB, *, PEGB4
			6'd2 : rdata = 41'b00011100000000001101111111000000011000000;
			// PEs: 37, 37 -> 
			// srcs: (172, 3)(3) 1, (264) 0 --> (318) 0:NM0, NI0, *, 
			6'd3 : rdata = 41'b00011100000000001010000000000000000000000;
			// PEs: 37, 37 -> 37
			// srcs: (175, 4)(97) 2, (318) 0 --> (372) 2:NW0, ALU, -, NW0
			6'd4 : rdata = 41'b00010010000000000011111111100100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 38) begin
	always @(*) begin
		case(address)
			// PEs: 38, 38 -> 
			// srcs: (1, 0)(43) 1, (98) -1 --> (152) -1:ND0, NW0, *, 
			6'd0 : rdata = 41'b00011011000000000100000000000000000000000;
			// PEs: 37, 38 -> 32
			// srcs: (4, 1)(151) 0, (152) -1 --> (202) -1:PENB, ALU, +, PEGB0
			6'd1 : rdata = 41'b00001110111111100011111111100000010000000;
			// PEs: 32, 38 -> 39
			// srcs: (170, 2)(225) 0, (43) 1 --> (265) 0:PEGB0, ND0, *, PENB
			6'd2 : rdata = 41'b00011111000000000110000000000000100000000;
			// PEs: 38, 39 -> 38
			// srcs: (179, 3)(98) -1, (319) 0 --> (373) -1:NW0, PEGB7, -, NW0
			6'd3 : rdata = 41'b00010010000000001110000111000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 39) begin
	always @(*) begin
		case(address)
			// PEs: 39, 39 -> 32
			// srcs: (1, 0)(45) 2, (100) -1 --> (154) -2:ND0, NW0, *, PENB
			6'd0 : rdata = 41'b00011011000000000100000000000000100000000;
			// PEs: 32, 39 -> 39
			// srcs: (172, 1)(225) 0, (45) 2 --> (267) 0:PEGB0, ND0, *, NI0
			6'd1 : rdata = 41'b00011111000000000110000000010000000000000;
			// PEs: 39, 38 -> 38
			// srcs: (173, 2)(3) 1, (265) 0 --> (319) 0:NM0, PENB, *, PEGB6
			6'd2 : rdata = 41'b00011100000000001101111111000000011100000;
			// PEs: 39, 39 -> 
			// srcs: (175, 3)(3) 1, (267) 0 --> (321) 0:NM0, NI0, *, 
			6'd3 : rdata = 41'b00011100000000001010000000000000000000000;
			// PEs: 39, 39 -> 39
			// srcs: (178, 4)(100) -1, (321) 0 --> (375) -1:NW0, ALU, -, NW0
			6'd4 : rdata = 41'b00010010000000000011111111100100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 40) begin
	always @(*) begin
		case(address)
			// PEs: 32 -> 41
			// srcs: (5, 0)(154) -2 --> (154) -2:PUNB, pass, PENB
			6'd0 : rdata = 41'b11000110111111110000000000000000100000000;
			// PEs: 47 -> 56
			// srcs: (6, 2)(212) 0 --> (212) 0:PENB, pass, PUGB7
			6'd1 : rdata = 41'b11000110111111100000000000000000000001111;
			// PEs: 56 -> 41
			// srcs: (13, 1)(160) 2 --> (160) 2:PUGB7, pass, PENB
			6'd2 : rdata = 41'b11000111000011110000000000000000100000000;
			// PEs: 42 -> 0
			// srcs: (25, 7)(211) 1 --> (211) 1:PEGB2, pass, PUGB0
			6'd3 : rdata = 41'b11000111000001000000000000000000000001000;
			// PEs: 56 -> 40
			// srcs: (33, 3)(187) 9 --> (187) 9:PUGB7, pass, NI0
			6'd4 : rdata = 41'b11000111000011110000000000010000000000000;
			// PEs: 24 -> 41
			// srcs: (34, 4)(189) 2 --> (189) 2:PUGB3, pass, PENB
			6'd5 : rdata = 41'b11000111000001110000000000000000100000000;
			// PEs: 40 -> 41
			// srcs: (40, 5)(187) 9 --> (187) 9:NI0, pass, PENB
			6'd6 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 32 -> 41
			// srcs: (50, 6)(185) 9 --> (185) 9:PUNB, pass, PENB
			6'd7 : rdata = 41'b11000110111111110000000000000000100000000;
			// PEs: 41 -> 48
			// srcs: (58, 8)(191) 20 --> (191) 20:PEGB1, pass, PUNB
			6'd8 : rdata = 41'b11000111000000100000000000000001000000000;
			// PEs: 56 -> 41
			// srcs: (168, 9)(225) 0 --> (225) 0:PUGB7, pass, PENB
			6'd9 : rdata = 41'b11000111000011110000000000000000100000000;
			// PEs: 56 -> 42
			// srcs: (169, 10)(225) 0 --> (225) 0:PUGB7, pass, PEGB2
			6'd10 : rdata = 41'b11000111000011110000000000000000010100000;
			// PEs: 56 -> 43
			// srcs: (170, 11)(225) 0 --> (225) 0:PUGB7, pass, PEGB3
			6'd11 : rdata = 41'b11000111000011110000000000000000010110000;
			// PEs: 56 -> 44
			// srcs: (171, 12)(225) 0 --> (225) 0:PUGB7, pass, PEGB4
			6'd12 : rdata = 41'b11000111000011110000000000000000011000000;
			// PEs: 56 -> 45
			// srcs: (172, 13)(225) 0 --> (225) 0:PUGB7, pass, PEGB5
			6'd13 : rdata = 41'b11000111000011110000000000000000011010000;
			// PEs: 56 -> 46
			// srcs: (174, 14)(225) 0 --> (225) 0:PUGB7, pass, PEGB6
			6'd14 : rdata = 41'b11000111000011110000000000000000011100000;
			// PEs: 56 -> 47
			// srcs: (175, 15)(225) 0 --> (225) 0:PUGB7, pass, PEGB7
			6'd15 : rdata = 41'b11000111000011110000000000000000011110000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 41) begin
	always @(*) begin
		case(address)
			// PEs: 41, 41 -> 
			// srcs: (1, 0)(46) -1, (101) 0 --> (155) 0:ND0, NW0, *, 
			6'd0 : rdata = 41'b00011011000000000100000000000000000000000;
			// PEs: 40, 41 -> 42
			// srcs: (8, 1)(154) -2, (155) 0 --> (206) -2:PENB, ALU, +, PENB
			6'd1 : rdata = 41'b00001110111111100011111111100000100000000;
			// PEs: 45, 40 -> 42
			// srcs: (17, 2)(209) -2, (160) 2 --> (210) 0:PEGB5, PENB, +, PENB
			6'd2 : rdata = 41'b00001111000010101101111111000000100000000;
			// PEs: 40 -> 
			// srcs: (36, 3)(189) 2 --> (189) 2:PENB, pass, 
			6'd3 : rdata = 41'b11000110111111100000000000000000000000000;
			// PEs: 40, 41 -> 
			// srcs: (42, 4)(187) 9, (189) 2 --> (190) 11:PENB, ALU, +, 
			6'd4 : rdata = 41'b00001110111111100011111111100000000000000;
			// PEs: 40, 41 -> 40
			// srcs: (53, 5)(185) 9, (190) 11 --> (191) 20:PENB, ALU, +, PEGB0
			6'd5 : rdata = 41'b00001110111111100011111111100000010000000;
			// PEs: 40, 41 -> 42
			// srcs: (170, 6)(225) 0, (46) -1 --> (268) 0:PENB, ND0, *, PENB
			6'd6 : rdata = 41'b00011110111111100110000000000000100000000;
			// PEs: 41, 42 -> 41
			// srcs: (179, 7)(101) 0, (322) 0 --> (376) 0:NW0, PEGB2, -, NW0
			6'd7 : rdata = 41'b00010010000000001110000010000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 42) begin
	always @(*) begin
		case(address)
			// PEs: 42, 42 -> 43
			// srcs: (1, 0)(47) 0, (102) 1 --> (156) 0:ND0, NW0, *, PENB
			6'd0 : rdata = 41'b00011011000000000100000000000000100000000;
			// PEs: 41, 43 -> 
			// srcs: (14, 1)(206) -2, (207) 3 --> (208) 1:PENB, PEGB3, +, 
			6'd1 : rdata = 41'b00001110111111101110000011000000000000000;
			// PEs: 42, 41 -> 40
			// srcs: (20, 2)(208) 1, (210) 0 --> (211) 1:ALU, PENB, +, PEGB0
			6'd2 : rdata = 41'b00001001111111111101111111000000010000000;
			// PEs: 42, 41 -> 41
			// srcs: (173, 4)(3) 1, (268) 0 --> (322) 0:NM0, PENB, *, PEGB1
			6'd3 : rdata = 41'b00011100000000001101111111000000010010000;
			// PEs: 40, 42 -> 43
			// srcs: (174, 3)(225) 0, (47) 0 --> (269) 0:PEGB0, ND0, *, PENB
			6'd4 : rdata = 41'b00011111000000000110000000000000100000000;
			// PEs: 42, 43 -> 42
			// srcs: (183, 5)(102) 1, (323) 0 --> (377) 1:NW0, PEGB3, -, NW0
			6'd5 : rdata = 41'b00010010000000001110000011000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 43) begin
	always @(*) begin
		case(address)
			// PEs: 43, 43 -> 
			// srcs: (1, 0)(48) -1, (103) -3 --> (157) 3:ND0, NW0, *, 
			6'd0 : rdata = 41'b00011011000000000100000000000000000000000;
			// PEs: 42, 43 -> 42
			// srcs: (4, 1)(156) 0, (157) 3 --> (207) 3:PENB, ALU, +, PEGB2
			6'd1 : rdata = 41'b00001110111111100011111111100000010100000;
			// PEs: 40, 43 -> 44
			// srcs: (175, 2)(225) 0, (48) -1 --> (270) 0:PEGB0, ND0, *, PENB
			6'd2 : rdata = 41'b00011111000000000110000000000000100000000;
			// PEs: 43, 42 -> 42
			// srcs: (177, 3)(3) 1, (269) 0 --> (323) 0:NM0, PENB, *, PEGB2
			6'd3 : rdata = 41'b00011100000000001101111111000000010100000;
			// PEs: 43, 44 -> 43
			// srcs: (184, 4)(103) -3, (324) 0 --> (378) -3:NW0, PEGB4, -, NW0
			6'd4 : rdata = 41'b00010010000000001110000100000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 44) begin
	always @(*) begin
		case(address)
			// PEs: 44, 44 -> 45
			// srcs: (1, 0)(49) 2, (104) -3 --> (158) -6:ND0, NW0, *, PENB
			6'd0 : rdata = 41'b00011011000000000100000000000000100000000;
			// PEs: 40, 44 -> 44
			// srcs: (176, 1)(225) 0, (49) 2 --> (271) 0:PEGB0, ND0, *, NI0
			6'd1 : rdata = 41'b00011111000000000110000000010000000000000;
			// PEs: 44, 43 -> 43
			// srcs: (178, 2)(3) 1, (270) 0 --> (324) 0:NM0, PENB, *, PEGB3
			6'd2 : rdata = 41'b00011100000000001101111111000000010110000;
			// PEs: 44, 44 -> 
			// srcs: (179, 3)(3) 1, (271) 0 --> (325) 0:NM0, NI0, *, 
			6'd3 : rdata = 41'b00011100000000001010000000000000000000000;
			// PEs: 44, 44 -> 44
			// srcs: (182, 4)(104) -3, (325) 0 --> (379) -3:NW0, ALU, -, NW0
			6'd4 : rdata = 41'b00010010000000000011111111100100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 45) begin
	always @(*) begin
		case(address)
			// PEs: 45, 45 -> 
			// srcs: (1, 0)(50) -2, (105) -2 --> (159) 4:ND0, NW0, *, 
			6'd0 : rdata = 41'b00011011000000000100000000000000000000000;
			// PEs: 44, 45 -> 41
			// srcs: (4, 1)(158) -6, (159) 4 --> (209) -2:PENB, ALU, +, PEGB1
			6'd1 : rdata = 41'b00001110111111100011111111100000010010000;
			// PEs: 40, 45 -> 46
			// srcs: (177, 2)(225) 0, (50) -2 --> (272) 0:PEGB0, ND0, *, PENB
			6'd2 : rdata = 41'b00011111000000000110000000000000100000000;
			// PEs: 45, 46 -> 45
			// srcs: (186, 3)(105) -2, (326) 0 --> (380) -2:NW0, PEGB6, -, NW0
			6'd3 : rdata = 41'b00010010000000001110000110000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 46) begin
	always @(*) begin
		case(address)
			// PEs: 46, 46 -> 47
			// srcs: (1, 0)(52) -3, (107) 0 --> (161) 0:ND0, NW0, *, PENB
			6'd0 : rdata = 41'b00011011000000000100000000000000100000000;
			// PEs: 40, 46 -> 46
			// srcs: (179, 1)(225) 0, (52) -3 --> (274) 0:PEGB0, ND0, *, NI0
			6'd1 : rdata = 41'b00011111000000000110000000010000000000000;
			// PEs: 46, 45 -> 45
			// srcs: (180, 2)(3) 1, (272) 0 --> (326) 0:NM0, PENB, *, PEGB5
			6'd2 : rdata = 41'b00011100000000001101111111000000011010000;
			// PEs: 46, 46 -> 
			// srcs: (182, 3)(3) 1, (274) 0 --> (328) 0:NM0, NI0, *, 
			6'd3 : rdata = 41'b00011100000000001010000000000000000000000;
			// PEs: 46, 46 -> 46
			// srcs: (185, 4)(107) 0, (328) 0 --> (382) 0:NW0, ALU, -, NW0
			6'd4 : rdata = 41'b00010010000000000011111111100100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 47) begin
	always @(*) begin
		case(address)
			// PEs: 47, 47 -> 
			// srcs: (1, 0)(53) 0, (108) -1 --> (162) 0:ND0, NW0, *, 
			6'd0 : rdata = 41'b00011011000000000100000000000000000000000;
			// PEs: 46, 47 -> 40
			// srcs: (4, 1)(161) 0, (162) 0 --> (212) 0:PENB, ALU, +, PENB
			6'd1 : rdata = 41'b00001110111111100011111111100000100000000;
			// PEs: 40, 47 -> 
			// srcs: (180, 2)(225) 0, (53) 0 --> (275) 0:PEGB0, ND0, *, 
			6'd2 : rdata = 41'b00011111000000000110000000000000000000000;
			// PEs: 47, 47 -> 
			// srcs: (183, 3)(3) 1, (275) 0 --> (329) 0:NM0, ALU, *, 
			6'd3 : rdata = 41'b00011100000000000011111111100000000000000;
			// PEs: 47, 47 -> 47
			// srcs: (186, 4)(108) -1, (329) 0 --> (383) -1:NW0, ALU, -, NW0
			6'd4 : rdata = 41'b00010010000000000011111111100100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 48) begin
	always @(*) begin
		case(address)
			// PEs: 55 -> 24
			// srcs: (3, 4)(139) 0 --> (139) 0:PENB, pass, PUGB3
			6'd0 : rdata = 41'b11000110111111100000000000000000000001011;
			// PEs: 51 -> 16
			// srcs: (6, 0)(119) -2 --> (119) -2:PEGB3, pass, PUGB2
			6'd1 : rdata = 41'b11000111000001100000000000000000000001010;
			// PEs: 52 -> 32
			// srcs: (7, 1)(126) 4 --> (126) 4:PEGB4, pass, PUGB4
			6'd2 : rdata = 41'b11000111000010000000000000000000000001100;
			// PEs: 54 -> 56
			// srcs: (8, 3)(136) 4 --> (136) 4:PEGB6, pass, PUNB
			6'd3 : rdata = 41'b11000111000011000000000000000001000000000;
			// PEs: 50 -> 56
			// srcs: (9, 5)(214) 4 --> (214) 4:PEGB2, pass, PUNB
			6'd4 : rdata = 41'b11000111000001000000000000000001000000000;
			// PEs: 16 -> 49
			// srcs: (14, 2)(183) 9 --> (183) 9:PUGB2, pass, PENB
			6'd5 : rdata = 41'b11000111000001010000000000000000100000000;
			// PEs: 0 -> 48
			// srcs: (22, 6)(169) 13 --> (169) 13:PUGB0, pass, NI0
			6'd6 : rdata = 41'b11000111000000010000000000010000000000000;
			// PEs: 49 -> 32
			// srcs: (23, 9)(184) 7 --> (184) 7:PEGB1, pass, PUGB4
			6'd7 : rdata = 41'b11000111000000100000000000000000000001100;
			// PEs: 16 -> 49
			// srcs: (33, 7)(171) -5 --> (171) -5:PUGB2, pass, PENB
			6'd8 : rdata = 41'b11000111000001010000000000000000100000000;
			// PEs: 48 -> 49
			// srcs: (40, 8)(169) 13 --> (169) 13:NI0, pass, PENB
			6'd9 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 24 -> 49
			// srcs: (52, 10)(178) 4 --> (178) 4:PUGB3, pass, PENB
			6'd10 : rdata = 41'b11000111000001110000000000000000100000000;
			// PEs: 40 -> 49
			// srcs: (60, 11)(191) 20 --> (191) 20:PUNB, pass, PENB
			6'd11 : rdata = 41'b11000110111111110000000000000000100000000;
			// PEs: 49 -> 32
			// srcs: (70, 12)(192) 32 --> (192) 32:PEGB1, pass, PUGB4
			6'd12 : rdata = 41'b11000111000000100000000000000000000001100;
			// PEs: 56 -> 51
			// srcs: (133, 13)(225) 0 --> (225) 0:PUGB7, pass, PEGB3
			6'd13 : rdata = 41'b11000111000011110000000000000000010110000;
			// PEs: 56 -> 52
			// srcs: (140, 14)(225) 0 --> (225) 0:PUGB7, pass, PEGB4
			6'd14 : rdata = 41'b11000111000011110000000000000000011000000;
			// PEs: 56 -> 53
			// srcs: (147, 15)(225) 0 --> (225) 0:PUGB7, pass, PEGB5
			6'd15 : rdata = 41'b11000111000011110000000000000000011010000;
			// PEs: 56 -> 54
			// srcs: (150, 16)(225) 0 --> (225) 0:PUGB7, pass, PEGB6
			6'd16 : rdata = 41'b11000111000011110000000000000000011100000;
			// PEs: 56 -> 55
			// srcs: (153, 17)(225) 0 --> (225) 0:PUGB7, pass, PEGB7
			6'd17 : rdata = 41'b11000111000011110000000000000000011110000;
			// PEs: 56 -> 49
			// srcs: (177, 18)(225) 0 --> (225) 0:PUGB7, pass, PENB
			6'd18 : rdata = 41'b11000111000011110000000000000000100000000;
			// PEs: 56 -> 50
			// srcs: (178, 19)(225) 0 --> (225) 0:PUGB7, pass, PEGB2
			6'd19 : rdata = 41'b11000111000011110000000000000000010100000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 49) begin
	always @(*) begin
		case(address)
			// PEs: 49, 49 -> 50
			// srcs: (1, 0)(55) 0, (110) -2 --> (164) 0:ND0, NW0, *, PENB
			6'd0 : rdata = 41'b00011011000000000100000000000000100000000;
			// PEs: 48, 53 -> 48
			// srcs: (17, 1)(183) 9, (133) -2 --> (184) 7:PENB, PEGB5, +, PEGB0
			6'd1 : rdata = 41'b00001110111111101110000101000000010000000;
			// PEs: 48 -> 
			// srcs: (35, 2)(171) -5 --> (171) -5:PENB, pass, 
			6'd2 : rdata = 41'b11000110111111100000000000000000000000000;
			// PEs: 48, 49 -> 
			// srcs: (42, 3)(169) 13, (171) -5 --> (172) 8:PENB, ALU, +, 
			6'd3 : rdata = 41'b00001110111111100011111111100000000000000;
			// PEs: 49, 48 -> 
			// srcs: (55, 4)(172) 8, (178) 4 --> (179) 12:ALU, PENB, +, 
			6'd4 : rdata = 41'b00001001111111111101111111000000000000000;
			// PEs: 49, 48 -> 48
			// srcs: (65, 5)(179) 12, (191) 20 --> (192) 32:ALU, PENB, +, PEGB0
			6'd5 : rdata = 41'b00001001111111111101111111000000010000000;
			// PEs: 48, 49 -> 50
			// srcs: (179, 6)(225) 0, (55) 0 --> (277) 0:PENB, ND0, *, PENB
			6'd6 : rdata = 41'b00011110111111100110000000000000100000000;
			// PEs: 49, 50 -> 49
			// srcs: (188, 7)(110) -2, (331) 0 --> (385) -2:NW0, PEGB2, -, NW0
			6'd7 : rdata = 41'b00010010000000001110000010000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 50) begin
	always @(*) begin
		case(address)
			// PEs: 50, 50 -> 
			// srcs: (1, 0)(56) -2, (111) -2 --> (165) 4:ND0, NW0, *, 
			6'd0 : rdata = 41'b00011011000000000100000000000000000000000;
			// PEs: 49, 50 -> 48
			// srcs: (4, 1)(164) 0, (165) 4 --> (214) 4:PENB, ALU, +, PEGB0
			6'd1 : rdata = 41'b00001110111111100011111111100000010000000;
			// PEs: 50, 49 -> 49
			// srcs: (182, 3)(3) 1, (277) 0 --> (331) 0:NM0, PENB, *, PEGB1
			6'd2 : rdata = 41'b00011100000000001101111111000000010010000;
			// PEs: 48, 50 -> 51
			// srcs: (183, 2)(225) 0, (56) -2 --> (278) 0:PEGB0, ND0, *, PENB
			6'd3 : rdata = 41'b00011111000000000110000000000000100000000;
			// PEs: 50, 51 -> 50
			// srcs: (192, 4)(111) -2, (332) 0 --> (386) -2:NW0, PEGB3, -, NW0
			6'd4 : rdata = 41'b00010010000000001110000011000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 51) begin
	always @(*) begin
		case(address)
			// PEs: 51, 51 -> 48
			// srcs: (1, 0)(10) -1, (65) 2 --> (119) -2:ND0, NW0, *, PEGB0
			6'd0 : rdata = 41'b00011011000000000100000000000000010000000;
			// PEs: 48, 51 -> 
			// srcs: (138, 1)(225) 0, (10) -1 --> (232) 0:PEGB0, ND0, *, 
			6'd1 : rdata = 41'b00011111000000000110000000000000000000000;
			// PEs: 51, 51 -> 
			// srcs: (141, 2)(3) 1, (232) 0 --> (286) 0:NM0, ALU, *, 
			6'd2 : rdata = 41'b00011100000000000011111111100000000000000;
			// PEs: 51, 51 -> 51
			// srcs: (144, 4)(65) 2, (286) 0 --> (340) 2:NW0, ALU, -, NW0
			6'd3 : rdata = 41'b00010010000000000011111111100100000000000;
			// PEs: 51, 50 -> 50
			// srcs: (186, 3)(3) 1, (278) 0 --> (332) 0:NM0, PENB, *, PEGB2
			6'd4 : rdata = 41'b00011100000000001101111111000000010100000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 52) begin
	always @(*) begin
		case(address)
			// PEs: 52, 52 -> 48
			// srcs: (1, 0)(17) -2, (72) -2 --> (126) 4:ND0, NW0, *, PEGB0
			6'd0 : rdata = 41'b00011011000000000100000000000000010000000;
			// PEs: 48, 52 -> 
			// srcs: (145, 1)(225) 0, (17) -2 --> (239) 0:PEGB0, ND0, *, 
			6'd1 : rdata = 41'b00011111000000000110000000000000000000000;
			// PEs: 52, 52 -> 
			// srcs: (148, 2)(3) 1, (239) 0 --> (293) 0:NM0, ALU, *, 
			6'd2 : rdata = 41'b00011100000000000011111111100000000000000;
			// PEs: 52, 52 -> 52
			// srcs: (151, 3)(72) -2, (293) 0 --> (347) -2:NW0, ALU, -, NW0
			6'd3 : rdata = 41'b00010010000000000011111111100100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 53) begin
	always @(*) begin
		case(address)
			// PEs: 53, 53 -> 49
			// srcs: (1, 0)(24) 1, (79) -2 --> (133) -2:ND0, NW0, *, PEGB1
			6'd0 : rdata = 41'b00011011000000000100000000000000010010000;
			// PEs: 48, 53 -> 
			// srcs: (152, 1)(225) 0, (24) 1 --> (246) 0:PEGB0, ND0, *, 
			6'd1 : rdata = 41'b00011111000000000110000000000000000000000;
			// PEs: 53, 53 -> 
			// srcs: (155, 2)(3) 1, (246) 0 --> (300) 0:NM0, ALU, *, 
			6'd2 : rdata = 41'b00011100000000000011111111100000000000000;
			// PEs: 53, 53 -> 53
			// srcs: (158, 3)(79) -2, (300) 0 --> (354) -2:NW0, ALU, -, NW0
			6'd3 : rdata = 41'b00010010000000000011111111100100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 54) begin
	always @(*) begin
		case(address)
			// PEs: 54, 54 -> 48
			// srcs: (1, 0)(27) 2, (82) 2 --> (136) 4:ND0, NW0, *, PEGB0
			6'd0 : rdata = 41'b00011011000000000100000000000000010000000;
			// PEs: 48, 54 -> 
			// srcs: (155, 1)(225) 0, (27) 2 --> (249) 0:PEGB0, ND0, *, 
			6'd1 : rdata = 41'b00011111000000000110000000000000000000000;
			// PEs: 54, 54 -> 
			// srcs: (158, 2)(3) 1, (249) 0 --> (303) 0:NM0, ALU, *, 
			6'd2 : rdata = 41'b00011100000000000011111111100000000000000;
			// PEs: 54, 54 -> 54
			// srcs: (161, 3)(82) 2, (303) 0 --> (357) 2:NW0, ALU, -, NW0
			6'd3 : rdata = 41'b00010010000000000011111111100100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 55) begin
	always @(*) begin
		case(address)
			// PEs: 55, 55 -> 48
			// srcs: (1, 0)(30) 0, (85) -3 --> (139) 0:ND0, NW0, *, PENB
			6'd0 : rdata = 41'b00011011000000000100000000000000100000000;
			// PEs: 48, 55 -> 
			// srcs: (158, 1)(225) 0, (30) 0 --> (252) 0:PEGB0, ND0, *, 
			6'd1 : rdata = 41'b00011111000000000110000000000000000000000;
			// PEs: 55, 55 -> 
			// srcs: (161, 2)(3) 1, (252) 0 --> (306) 0:NM0, ALU, *, 
			6'd2 : rdata = 41'b00011100000000000011111111100000000000000;
			// PEs: 55, 55 -> 55
			// srcs: (164, 3)(85) -3, (306) 0 --> (360) -3:NW0, ALU, -, NW0
			6'd3 : rdata = 41'b00010010000000000011111111100100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 56) begin
	always @(*) begin
		case(address)
			// PEs: 57 -> 0
			// srcs: (6, 3)(146) 6 --> (146) 6:PEGB1, pass, PUNB
			6'd0 : rdata = 41'b11000111000000100000000000000001000000000;
			// PEs: 58 -> 8
			// srcs: (7, 4)(153) 9 --> (153) 9:PEGB2, pass, PUGB1
			6'd1 : rdata = 41'b11000111000001000000000000000000000001001;
			// PEs: 59 -> 40
			// srcs: (8, 5)(160) 2 --> (160) 2:PEGB3, pass, PUGB5
			6'd2 : rdata = 41'b11000111000001100000000000000000000001101;
			// PEs: 48 -> 56
			// srcs: (10, 1)(136) 4 --> (136) 4:PUNB, pass, NI0
			6'd3 : rdata = 41'b11000110111111110000000000010000000000000;
			// PEs: 16 -> 57
			// srcs: (15, 0)(186) 5 --> (186) 5:PUGB2, pass, PENB
			6'd4 : rdata = 41'b11000111000001010000000000000000100000000;
			// PEs: 56 -> 57
			// srcs: (21, 2)(136) 4 --> (136) 4:NI0, pass, PENB
			6'd5 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 40 -> 57
			// srcs: (22, 6)(212) 0 --> (212) 0:PUGB5, pass, PENB
			6'd6 : rdata = 41'b11000111000010110000000000000000100000000;
			// PEs: 48 -> 57
			// srcs: (23, 7)(214) 4 --> (214) 4:PUNB, pass, PENB
			6'd7 : rdata = 41'b11000110111111110000000000000000100000000;
			// PEs: 57 -> 40
			// srcs: (28, 8)(187) 9 --> (187) 9:PEGB1, pass, PUGB5
			6'd8 : rdata = 41'b11000111000000100000000000000000000001101;
			// PEs: 58 -> 0
			// srcs: (39, 9)(216) 0 --> (216) 0:PEGB2, pass, PUNB
			6'd9 : rdata = 41'b11000111000001000000000000000001000000000;
			// PEs: 32 -> 62
			// srcs: (101, 10)(219) 76 --> (219) 76:PUGB4, pass, PEGB6
			6'd10 : rdata = 41'b11000111000010010000000000000000011100000;
			// PEs: 63 -> 0
			// srcs: (119, 11)(225) 0 --> (225) 0:PENB, pass, PUNB
			6'd11 : rdata = 41'b11000110111111100000000000000001000000000;
			// PEs: 63 -> 0
			// srcs: (123, 12)(225) 0 --> (225) 0:PENB, pass, PUNB
			6'd12 : rdata = 41'b11000110111111100000000000000001000000000;
			// PEs: 63 -> 0
			// srcs: (124, 13)(225) 0 --> (225) 0:PENB, pass, PUNB
			6'd13 : rdata = 41'b11000110111111100000000000000001000000000;
			// PEs: 63 -> 0
			// srcs: (125, 14)(225) 0 --> (225) 0:PENB, pass, PUNB
			6'd14 : rdata = 41'b11000110111111100000000000000001000000000;
			// PEs: 63 -> 0
			// srcs: (126, 15)(225) 0 --> (225) 0:PENB, pass, PUNB
			6'd15 : rdata = 41'b11000110111111100000000000000001000000000;
			// PEs: 63 -> 0
			// srcs: (127, 16)(225) 0 --> (225) 0:PENB, pass, PUNB
			6'd16 : rdata = 41'b11000110111111100000000000000001000000000;
			// PEs: 63 -> 48
			// srcs: (128, 17)(225) 0 --> (225) 0:PENB, pass, PUGB6
			6'd17 : rdata = 41'b11000110111111100000000000000000000001110;
			// PEs: 63 -> 0
			// srcs: (129, 18)(225) 0 --> (225) 0:PENB, pass, PUNB
			6'd18 : rdata = 41'b11000110111111100000000000000001000000000;
			// PEs: 63 -> 8
			// srcs: (130, 19)(225) 0 --> (225) 0:PENB, pass, PUGB1
			6'd19 : rdata = 41'b11000110111111100000000000000000000001001;
			// PEs: 63 -> 8
			// srcs: (131, 20)(225) 0 --> (225) 0:PENB, pass, PUGB1
			6'd20 : rdata = 41'b11000110111111100000000000000000000001001;
			// PEs: 63 -> 8
			// srcs: (132, 21)(225) 0 --> (225) 0:PENB, pass, PUGB1
			6'd21 : rdata = 41'b11000110111111100000000000000000000001001;
			// PEs: 63 -> 8
			// srcs: (133, 22)(225) 0 --> (225) 0:PENB, pass, PUGB1
			6'd22 : rdata = 41'b11000110111111100000000000000000000001001;
			// PEs: 63 -> 8
			// srcs: (134, 23)(225) 0 --> (225) 0:PENB, pass, PUGB1
			6'd23 : rdata = 41'b11000110111111100000000000000000000001001;
			// PEs: 63 -> 48
			// srcs: (135, 24)(225) 0 --> (225) 0:PENB, pass, PUGB6
			6'd24 : rdata = 41'b11000110111111100000000000000000000001110;
			// PEs: 63 -> 8
			// srcs: (136, 25)(225) 0 --> (225) 0:PENB, pass, PUGB1
			6'd25 : rdata = 41'b11000110111111100000000000000000000001001;
			// PEs: 63 -> 8
			// srcs: (137, 26)(225) 0 --> (225) 0:PENB, pass, PUGB1
			6'd26 : rdata = 41'b11000110111111100000000000000000000001001;
			// PEs: 63 -> 16
			// srcs: (138, 27)(225) 0 --> (225) 0:PENB, pass, PUGB2
			6'd27 : rdata = 41'b11000110111111100000000000000000000001010;
			// PEs: 63 -> 16
			// srcs: (139, 28)(225) 0 --> (225) 0:PENB, pass, PUGB2
			6'd28 : rdata = 41'b11000110111111100000000000000000000001010;
			// PEs: 63 -> 16
			// srcs: (140, 29)(225) 0 --> (225) 0:PENB, pass, PUGB2
			6'd29 : rdata = 41'b11000110111111100000000000000000000001010;
			// PEs: 63 -> 16
			// srcs: (141, 30)(225) 0 --> (225) 0:PENB, pass, PUGB2
			6'd30 : rdata = 41'b11000110111111100000000000000000000001010;
			// PEs: 63 -> 48
			// srcs: (142, 31)(225) 0 --> (225) 0:PENB, pass, PUGB6
			6'd31 : rdata = 41'b11000110111111100000000000000000000001110;
			// PEs: 63 -> 16
			// srcs: (143, 32)(225) 0 --> (225) 0:PENB, pass, PUGB2
			6'd32 : rdata = 41'b11000110111111100000000000000000000001010;
			// PEs: 63 -> 16
			// srcs: (144, 33)(225) 0 --> (225) 0:PENB, pass, PUGB2
			6'd33 : rdata = 41'b11000110111111100000000000000000000001010;
			// PEs: 63 -> 48
			// srcs: (145, 34)(225) 0 --> (225) 0:PENB, pass, PUGB6
			6'd34 : rdata = 41'b11000110111111100000000000000000000001110;
			// PEs: 63 -> 16
			// srcs: (146, 35)(225) 0 --> (225) 0:PENB, pass, PUGB2
			6'd35 : rdata = 41'b11000110111111100000000000000000000001010;
			// PEs: 63 -> 24
			// srcs: (147, 36)(225) 0 --> (225) 0:PENB, pass, PUGB3
			6'd36 : rdata = 41'b11000110111111100000000000000000000001011;
			// PEs: 63 -> 48
			// srcs: (148, 37)(225) 0 --> (225) 0:PENB, pass, PUGB6
			6'd37 : rdata = 41'b11000110111111100000000000000000000001110;
			// PEs: 63 -> 24
			// srcs: (149, 38)(225) 0 --> (225) 0:PENB, pass, PUGB3
			6'd38 : rdata = 41'b11000110111111100000000000000000000001011;
			// PEs: 63 -> 24
			// srcs: (150, 39)(225) 0 --> (225) 0:PENB, pass, PUGB3
			6'd39 : rdata = 41'b11000110111111100000000000000000000001011;
			// PEs: 63 -> 24
			// srcs: (151, 40)(225) 0 --> (225) 0:PENB, pass, PUGB3
			6'd40 : rdata = 41'b11000110111111100000000000000000000001011;
			// PEs: 63 -> 24
			// srcs: (152, 41)(225) 0 --> (225) 0:PENB, pass, PUGB3
			6'd41 : rdata = 41'b11000110111111100000000000000000000001011;
			// PEs: 63 -> 24
			// srcs: (153, 42)(225) 0 --> (225) 0:PENB, pass, PUGB3
			6'd42 : rdata = 41'b11000110111111100000000000000000000001011;
			// PEs: 63 -> 24
			// srcs: (154, 43)(225) 0 --> (225) 0:PENB, pass, PUGB3
			6'd43 : rdata = 41'b11000110111111100000000000000000000001011;
			// PEs: 63 -> 32
			// srcs: (155, 44)(225) 0 --> (225) 0:PENB, pass, PUGB4
			6'd44 : rdata = 41'b11000110111111100000000000000000000001100;
			// PEs: 63 -> 32
			// srcs: (156, 45)(225) 0 --> (225) 0:PENB, pass, PUGB4
			6'd45 : rdata = 41'b11000110111111100000000000000000000001100;
			// PEs: 63 -> 32
			// srcs: (157, 46)(225) 0 --> (225) 0:PENB, pass, PUGB4
			6'd46 : rdata = 41'b11000110111111100000000000000000000001100;
			// PEs: 63 -> 32
			// srcs: (158, 47)(225) 0 --> (225) 0:PENB, pass, PUGB4
			6'd47 : rdata = 41'b11000110111111100000000000000000000001100;
			// PEs: 63 -> 32
			// srcs: (159, 48)(225) 0 --> (225) 0:PENB, pass, PUGB4
			6'd48 : rdata = 41'b11000110111111100000000000000000000001100;
			// PEs: 63 -> 32
			// srcs: (160, 49)(225) 0 --> (225) 0:PENB, pass, PUGB4
			6'd49 : rdata = 41'b11000110111111100000000000000000000001100;
			// PEs: 63 -> 32
			// srcs: (162, 50)(225) 0 --> (225) 0:PENB, pass, PUGB4
			6'd50 : rdata = 41'b11000110111111100000000000000000000001100;
			// PEs: 63 -> 40
			// srcs: (163, 51)(225) 0 --> (225) 0:PENB, pass, PUGB5
			6'd51 : rdata = 41'b11000110111111100000000000000000000001101;
			// PEs: 63 -> 40
			// srcs: (164, 52)(225) 0 --> (225) 0:PENB, pass, PUGB5
			6'd52 : rdata = 41'b11000110111111100000000000000000000001101;
			// PEs: 63 -> 40
			// srcs: (165, 53)(225) 0 --> (225) 0:PENB, pass, PUGB5
			6'd53 : rdata = 41'b11000110111111100000000000000000000001101;
			// PEs: 63 -> 40
			// srcs: (166, 54)(225) 0 --> (225) 0:PENB, pass, PUGB5
			6'd54 : rdata = 41'b11000110111111100000000000000000000001101;
			// PEs: 63 -> 40
			// srcs: (167, 55)(225) 0 --> (225) 0:PENB, pass, PUGB5
			6'd55 : rdata = 41'b11000110111111100000000000000000000001101;
			// PEs: 63 -> 40
			// srcs: (169, 56)(225) 0 --> (225) 0:PENB, pass, PUGB5
			6'd56 : rdata = 41'b11000110111111100000000000000000000001101;
			// PEs: 63 -> 40
			// srcs: (170, 57)(225) 0 --> (225) 0:PENB, pass, PUGB5
			6'd57 : rdata = 41'b11000110111111100000000000000000000001101;
			// PEs: 63 -> 48
			// srcs: (172, 58)(225) 0 --> (225) 0:PENB, pass, PUGB6
			6'd58 : rdata = 41'b11000110111111100000000000000000000001110;
			// PEs: 63 -> 48
			// srcs: (173, 59)(225) 0 --> (225) 0:PENB, pass, PUGB6
			6'd59 : rdata = 41'b11000110111111100000000000000000000001110;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 57) begin
	always @(*) begin
		case(address)
			// PEs: 57, 57 -> 56
			// srcs: (1, 0)(37) -2, (92) -3 --> (146) 6:ND0, NW0, *, PEGB0
			6'd0 : rdata = 41'b00011011000000000100000000000000010000000;
			// PEs: 56 -> 
			// srcs: (17, 1)(186) 5 --> (186) 5:PENB, pass, 
			6'd1 : rdata = 41'b11000110111111100000000000000000000000000;
			// PEs: 57, 56 -> 56
			// srcs: (23, 2)(186) 5, (136) 4 --> (187) 9:ALU, PENB, +, PEGB0
			6'd2 : rdata = 41'b00001001111111111101111111000000010000000;
			// PEs: 56, 60 -> 57
			// srcs: (24, 3)(212) 0, (163) -4 --> (213) -4:PENB, PEGB4, +, NI0
			6'd3 : rdata = 41'b00001110111111101110000100010000000000000;
			// PEs: 56, 61 -> 58
			// srcs: (25, 4)(214) 4, (166) 0 --> (215) 4:PENB, PEGB5, +, PENB
			6'd4 : rdata = 41'b00001110111111101110000101000000100000000;
			// PEs: 57 -> 58
			// srcs: (32, 5)(213) -4 --> (213) -4:NI0, pass, PENB
			6'd5 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 63, 57 -> 58
			// srcs: (123, 6)(225) 0, (37) -2 --> (259) 0:PEGB7, ND0, *, PENB
			6'd6 : rdata = 41'b00011111000011100110000000000000100000000;
			// PEs: 57, 58 -> 57
			// srcs: (132, 7)(92) -3, (313) 0 --> (367) -3:NW0, PEGB2, -, NW0
			6'd7 : rdata = 41'b00010010000000001110000010000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 58) begin
	always @(*) begin
		case(address)
			// PEs: 58, 58 -> 56
			// srcs: (1, 0)(44) -3, (99) -3 --> (153) 9:ND0, NW0, *, PEGB0
			6'd0 : rdata = 41'b00011011000000000100000000000000010000000;
			// PEs: 57 -> 
			// srcs: (27, 1)(215) 4 --> (215) 4:PENB, pass, 
			6'd1 : rdata = 41'b11000110111111100000000000000000000000000;
			// PEs: 57, 58 -> 56
			// srcs: (34, 2)(213) -4, (215) 4 --> (216) 0:PENB, ALU, +, PEGB0
			6'd2 : rdata = 41'b00001110111111100011111111100000010000000;
			// PEs: 58, 57 -> 57
			// srcs: (126, 4)(3) 1, (259) 0 --> (313) 0:NM0, PENB, *, PEGB1
			6'd3 : rdata = 41'b00011100000000001101111111000000010010000;
			// PEs: 63, 58 -> 59
			// srcs: (164, 3)(225) 0, (44) -3 --> (266) 0:PEGB7, ND0, *, PENB
			6'd4 : rdata = 41'b00011111000011100110000000000000100000000;
			// PEs: 58, 59 -> 58
			// srcs: (173, 5)(99) -3, (320) 0 --> (374) -3:NW0, PEGB3, -, NW0
			6'd5 : rdata = 41'b00010010000000001110000011000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 59) begin
	always @(*) begin
		case(address)
			// PEs: 59, 59 -> 56
			// srcs: (1, 0)(51) 1, (106) 2 --> (160) 2:ND0, NW0, *, PEGB0
			6'd0 : rdata = 41'b00011011000000000100000000000000010000000;
			// PEs: 59, 58 -> 58
			// srcs: (167, 2)(3) 1, (266) 0 --> (320) 0:NM0, PENB, *, PEGB2
			6'd1 : rdata = 41'b00011100000000001101111111000000010100000;
			// PEs: 63, 59 -> 
			// srcs: (171, 1)(225) 0, (51) 1 --> (273) 0:PEGB7, ND0, *, 
			6'd2 : rdata = 41'b00011111000011100110000000000000000000000;
			// PEs: 59, 59 -> 
			// srcs: (174, 3)(3) 1, (273) 0 --> (327) 0:NM0, ALU, *, 
			6'd3 : rdata = 41'b00011100000000000011111111100000000000000;
			// PEs: 59, 59 -> 59
			// srcs: (177, 4)(106) 2, (327) 0 --> (381) 2:NW0, ALU, -, NW0
			6'd4 : rdata = 41'b00010010000000000011111111100100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 60) begin
	always @(*) begin
		case(address)
			// PEs: 60, 60 -> 57
			// srcs: (1, 0)(54) 2, (109) -2 --> (163) -4:ND0, NW0, *, PEGB1
			6'd0 : rdata = 41'b00011011000000000100000000000000010010000;
			// PEs: 63, 60 -> 
			// srcs: (174, 1)(225) 0, (54) 2 --> (276) 0:PEGB7, ND0, *, 
			6'd1 : rdata = 41'b00011111000011100110000000000000000000000;
			// PEs: 60, 60 -> 
			// srcs: (177, 2)(3) 1, (276) 0 --> (330) 0:NM0, ALU, *, 
			6'd2 : rdata = 41'b00011100000000000011111111100000000000000;
			// PEs: 60, 60 -> 60
			// srcs: (180, 3)(109) -2, (330) 0 --> (384) -2:NW0, ALU, -, NW0
			6'd3 : rdata = 41'b00010010000000000011111111100100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 61) begin
	always @(*) begin
		case(address)
			// PEs: 61, 61 -> 57
			// srcs: (1, 0)(57) 0, (112) 0 --> (166) 0:ND0, NW0, *, PEGB1
			6'd0 : rdata = 41'b00011011000000000100000000000000010010000;
			// PEs: 63, 61 -> 
			// srcs: (177, 1)(225) 0, (57) 0 --> (279) 0:PEGB7, ND0, *, 
			6'd1 : rdata = 41'b00011111000011100110000000000000000000000;
			// PEs: 61, 61 -> 
			// srcs: (180, 2)(3) 1, (279) 0 --> (333) 0:NM0, ALU, *, 
			6'd2 : rdata = 41'b00011100000000000011111111100000000000000;
			// PEs: 61, 61 -> 61
			// srcs: (183, 3)(112) 0, (333) 0 --> (387) 0:NW0, ALU, -, NW0
			6'd3 : rdata = 41'b00010010000000000011111111100100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 62) begin
	always @(*) begin
		case(address)
			// PEs: 62, 62 -> 62
			// srcs: (1, 0)(221) 0, (58) 0 --> (222) 0:NM0, ND0, -, NI0
			6'd0 : rdata = 41'b00010100000000000110000000010000000000000;
			// PEs: 62, 56 -> 63
			// srcs: (107, 1)(58) 0, (219) 76 --> (220) 0:ND0, PEGB0, *, PENB
			6'd1 : rdata = 41'b00011011000000001110000000000000100000000;
			// PEs: 62 -> 63
			// srcs: (115, 2)(222) 0 --> (222) 0:NI0, pass, PENB
			6'd2 : rdata = 41'b11000101000000000000000000000000100000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 63) begin
	always @(*) begin
		case(address)
			// PEs: 62, 63 -> 
			// srcs: (110, 0)(220) 0, (223) 1 --> (224) 0:PENB, NM0, >, 
			6'd0 : rdata = 41'b00111110111111101000000000000000000000000;
			// PEs: 63, 62 -> 56, 57, 63
			// srcs: (117, 1)(224) 0, (222) 0 --> (225) 0:ALU, PENB, *, NI0, PENB, PEGB1
			6'd1 : rdata = 41'b00011001111111111101111111010000110010000;
			// PEs: 63 -> 56
			// srcs: (119, 2)(225) 0 --> (225) 0:ALU, pass, PENB
			6'd2 : rdata = 41'b11000001111111110000000000000000100000000;
			// PEs: 63 -> 56
			// srcs: (120, 3)(225) 0 --> (225) 0:NI0, pass, PENB
			6'd3 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 63 -> 56
			// srcs: (121, 4)(225) 0 --> (225) 0:NI0, pass, PENB
			6'd4 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 63 -> 56
			// srcs: (122, 5)(225) 0 --> (225) 0:NI0, pass, PENB
			6'd5 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 63 -> 56
			// srcs: (123, 6)(225) 0 --> (225) 0:NI0, pass, PENB
			6'd6 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 63 -> 56
			// srcs: (124, 7)(225) 0 --> (225) 0:NI0, pass, PENB
			6'd7 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 63 -> 56
			// srcs: (125, 8)(225) 0 --> (225) 0:NI0, pass, PENB
			6'd8 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 63 -> 56
			// srcs: (126, 9)(225) 0 --> (225) 0:NI0, pass, PENB
			6'd9 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 63 -> 56
			// srcs: (127, 10)(225) 0 --> (225) 0:NI0, pass, PENB
			6'd10 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 63 -> 56
			// srcs: (128, 11)(225) 0 --> (225) 0:NI0, pass, PENB
			6'd11 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 63 -> 56
			// srcs: (129, 12)(225) 0 --> (225) 0:NI0, pass, PENB
			6'd12 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 63 -> 56
			// srcs: (130, 13)(225) 0 --> (225) 0:NI0, pass, PENB
			6'd13 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 63 -> 56
			// srcs: (131, 14)(225) 0 --> (225) 0:NI0, pass, PENB
			6'd14 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 63 -> 56
			// srcs: (132, 15)(225) 0 --> (225) 0:NI0, pass, PENB
			6'd15 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 63 -> 56
			// srcs: (133, 16)(225) 0 --> (225) 0:NI0, pass, PENB
			6'd16 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 63 -> 56
			// srcs: (134, 17)(225) 0 --> (225) 0:NI0, pass, PENB
			6'd17 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 63 -> 56
			// srcs: (135, 18)(225) 0 --> (225) 0:NI0, pass, PENB
			6'd18 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 63 -> 56
			// srcs: (136, 19)(225) 0 --> (225) 0:NI0, pass, PENB
			6'd19 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 63 -> 56
			// srcs: (137, 20)(225) 0 --> (225) 0:NI0, pass, PENB
			6'd20 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 63 -> 56
			// srcs: (138, 21)(225) 0 --> (225) 0:NI0, pass, PENB
			6'd21 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 63 -> 56
			// srcs: (139, 22)(225) 0 --> (225) 0:NI0, pass, PENB
			6'd22 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 63 -> 56
			// srcs: (140, 23)(225) 0 --> (225) 0:NI0, pass, PENB
			6'd23 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 63 -> 56
			// srcs: (141, 24)(225) 0 --> (225) 0:NI0, pass, PENB
			6'd24 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 63 -> 56
			// srcs: (142, 25)(225) 0 --> (225) 0:NI0, pass, PENB
			6'd25 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 63 -> 56
			// srcs: (143, 26)(225) 0 --> (225) 0:NI0, pass, PENB
			6'd26 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 63 -> 56
			// srcs: (144, 27)(225) 0 --> (225) 0:NI0, pass, PENB
			6'd27 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 63 -> 56
			// srcs: (145, 28)(225) 0 --> (225) 0:NI0, pass, PENB
			6'd28 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 63 -> 56
			// srcs: (146, 29)(225) 0 --> (225) 0:NI0, pass, PENB
			6'd29 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 63 -> 56
			// srcs: (147, 30)(225) 0 --> (225) 0:NI0, pass, PENB
			6'd30 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 63 -> 56
			// srcs: (148, 31)(225) 0 --> (225) 0:NI0, pass, PENB
			6'd31 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 63 -> 56
			// srcs: (149, 32)(225) 0 --> (225) 0:NI0, pass, PENB
			6'd32 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 63 -> 56
			// srcs: (150, 33)(225) 0 --> (225) 0:NI0, pass, PENB
			6'd33 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 63 -> 56
			// srcs: (151, 34)(225) 0 --> (225) 0:NI0, pass, PENB
			6'd34 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 63 -> 56
			// srcs: (152, 35)(225) 0 --> (225) 0:NI0, pass, PENB
			6'd35 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 63 -> 56
			// srcs: (153, 36)(225) 0 --> (225) 0:NI0, pass, PENB
			6'd36 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 63 -> 56
			// srcs: (154, 37)(225) 0 --> (225) 0:NI0, pass, PENB
			6'd37 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 63 -> 56
			// srcs: (155, 38)(225) 0 --> (225) 0:NI0, pass, PENB
			6'd38 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 63 -> 56
			// srcs: (156, 39)(225) 0 --> (225) 0:NI0, pass, PENB
			6'd39 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 63 -> 58
			// srcs: (157, 40)(225) 0 --> (225) 0:NI0, pass, PEGB2
			6'd40 : rdata = 41'b11000101000000000000000000000000010100000;
			// PEs: 63 -> 56
			// srcs: (158, 41)(225) 0 --> (225) 0:NI0, pass, PENB
			6'd41 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 63 -> 56
			// srcs: (159, 42)(225) 0 --> (225) 0:NI0, pass, PENB
			6'd42 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 63 -> 56
			// srcs: (160, 43)(225) 0 --> (225) 0:NI0, pass, PENB
			6'd43 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 63 -> 56
			// srcs: (161, 44)(225) 0 --> (225) 0:NI0, pass, PENB
			6'd44 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 63 -> 56
			// srcs: (162, 45)(225) 0 --> (225) 0:NI0, pass, PENB
			6'd45 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 63 -> 56
			// srcs: (163, 46)(225) 0 --> (225) 0:NI0, pass, PENB
			6'd46 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 63 -> 59
			// srcs: (164, 47)(225) 0 --> (225) 0:NI0, pass, PEGB3
			6'd47 : rdata = 41'b11000101000000000000000000000000010110000;
			// PEs: 63 -> 56
			// srcs: (165, 48)(225) 0 --> (225) 0:NI0, pass, PENB
			6'd48 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 63 -> 56
			// srcs: (166, 49)(225) 0 --> (225) 0:NI0, pass, PENB
			6'd49 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 63 -> 60
			// srcs: (167, 50)(225) 0 --> (225) 0:NI0, pass, PEGB4
			6'd50 : rdata = 41'b11000101000000000000000000000000011000000;
			// PEs: 63 -> 56
			// srcs: (168, 51)(225) 0 --> (225) 0:NI0, pass, PENB
			6'd51 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 63 -> 56
			// srcs: (169, 52)(225) 0 --> (225) 0:NI0, pass, PENB
			6'd52 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 63 -> 61
			// srcs: (170, 53)(225) 0 --> (225) 0:NI0, pass, PEGB5
			6'd53 : rdata = 41'b11000101000000000000000000000000011010000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

endgenerate
/*****************************************************************************/
endmodule
