`timescale 1ns/1ps
module gaussian(
	in,
	out
);

	parameter dataLen = 16;
	parameter indexLen = 9;
	parameter fracLen = 7;

	input signed [dataLen - 1 : 0] in;
	output reg [dataLen - 1 : 0] out;
	reg [indexLen - 1 :0] index;

	always @(in)
	begin
		out = 0;
		if (in < -(8 << 7)) begin
			out = 0;
		end else if (in > (8 << 7)) begin
			out = 0;
		end else begin
		index[8]	= in[15];
		index[7:5]	= in[9:7];
		index[4:0]	= in[6:2];
		case(index)
			9'd256: out = 16'b0000000000000000; // input=-8.0, output=2.05232614558e-56
			9'd257: out = 16'b0000000000000000; // input=-7.96875, output=5.56791540596e-56
			9'd258: out = 16'b0000000000000000; // input=-7.9375, output=1.50467399787e-55
			9'd259: out = 16'b0000000000000000; // input=-7.90625, output=4.05037972923e-55
			9'd260: out = 16'b0000000000000000; // input=-7.875, output=1.0860569595e-54
			9'd261: out = 16'b0000000000000000; // input=-7.84375, output=2.90076804211e-54
			9'd262: out = 16'b0000000000000000; // input=-7.8125, output=7.71750533773e-54
			9'd263: out = 16'b0000000000000000; // input=-7.78125, output=2.04524063202e-53
			9'd264: out = 16'b0000000000000000; // input=-7.75, output=5.39902604918e-53
			9'd265: out = 16'b0000000000000000; // input=-7.71875, output=1.41967838716e-52
			9'd266: out = 16'b0000000000000000; // input=-7.6875, output=3.71850231248e-52
			9'd267: out = 16'b0000000000000000; // input=-7.65625, output=9.70174103983e-52
			9'd268: out = 16'b0000000000000000; // input=-7.625, output=2.52135987788e-51
			9'd269: out = 16'b0000000000000000; // input=-7.59375, output=6.52714911362e-51
			9'd270: out = 16'b0000000000000000; // input=-7.5625, output=1.68312266462e-50
			9'd271: out = 16'b0000000000000000; // input=-7.53125, output=4.32326183636e-50
			9'd272: out = 16'b0000000000000000; // input=-7.5, output=1.10614190997e-49
			9'd273: out = 16'b0000000000000000; // input=-7.46875, output=2.81912084447e-49
			9'd274: out = 16'b0000000000000000; // input=-7.4375, output=7.15681968385e-49
			9'd275: out = 16'b0000000000000000; // input=-7.40625, output=1.80979754616e-48
			9'd276: out = 16'b0000000000000000; // input=-7.375, output=4.55872560131e-48
			9'd277: out = 16'b0000000000000000; // input=-7.34375, output=1.14382726918e-47
			9'd278: out = 16'b0000000000000000; // input=-7.3125, output=2.85878159428e-47
			9'd279: out = 16'b0000000000000000; // input=-7.28125, output=7.1171324113e-47
			9'd280: out = 16'b0000000000000000; // input=-7.25, output=1.76495099492e-46
			9'd281: out = 16'b0000000000000000; // input=-7.21875, output=4.35977216421e-46
			9'd282: out = 16'b0000000000000000; // input=-7.1875, output=1.07274987899e-45
			9'd283: out = 16'b0000000000000000; // input=-7.15625, output=2.62927911298e-45
			9'd284: out = 16'b0000000000000000; // input=-7.125, output=6.41916362084e-45
			9'd285: out = 16'b0000000000000000; // input=-7.09375, output=1.56107488696e-44
			9'd286: out = 16'b0000000000000000; // input=-7.0625, output=3.78157367485e-44
			9'd287: out = 16'b0000000000000000; // input=-7.03125, output=9.12483314748e-44
			9'd288: out = 16'b0000000000000000; // input=-7.0, output=2.19321311878e-43
			9'd289: out = 16'b0000000000000000; // input=-6.96875, output=5.25097892486e-43
			9'd290: out = 16'b0000000000000000; // input=-6.9375, output=1.25228521358e-42
			9'd291: out = 16'b0000000000000000; // input=-6.90625, output=2.97488215993e-42
			9'd292: out = 16'b0000000000000000; // input=-6.875, output=7.03946767599e-42
			9'd293: out = 16'b0000000000000000; // input=-6.84375, output=1.65925604311e-41
			9'd294: out = 16'b0000000000000000; // input=-6.8125, output=3.89574510993e-41
			9'd295: out = 16'b0000000000000000; // input=-6.78125, output=9.11110806056e-41
			9'd296: out = 16'b0000000000000000; // input=-6.75, output=2.12253762783e-40
			9'd297: out = 16'b0000000000000000; // input=-6.71875, output=4.92541848268e-40
			9'd298: out = 16'b0000000000000000; // input=-6.6875, output=1.13850360632e-39
			9'd299: out = 16'b0000000000000000; // input=-6.65625, output=2.62137541904e-39
			9'd300: out = 16'b0000000000000000; // input=-6.625, output=6.0121190522e-39
			9'd301: out = 16'b0000000000000000; // input=-6.59375, output=1.37350251292e-38
			9'd302: out = 16'b0000000000000000; // input=-6.5625, output=3.12561067823e-38
			9'd303: out = 16'b0000000000000000; // input=-6.53125, output=7.08506506176e-38
			9'd304: out = 16'b0000000000000000; // input=-6.5, output=1.5997655514e-37
			9'd305: out = 16'b0000000000000000; // input=-6.46875, output=3.59809292893e-37
			9'd306: out = 16'b0000000000000000; // input=-6.4375, output=8.06105618402e-37
			9'd307: out = 16'b0000000000000000; // input=-6.40625, output=1.79893328563e-36
			9'd308: out = 16'b0000000000000000; // input=-6.375, output=3.99891068444e-36
			9'd309: out = 16'b0000000000000000; // input=-6.34375, output=8.85465996484e-36
			9'd310: out = 16'b0000000000000000; // input=-6.3125, output=1.9530151363e-35
			9'd311: out = 16'b0000000000000000; // input=-6.28125, output=4.29084540294e-35
			9'd312: out = 16'b0000000000000000; // input=-6.25, output=9.39039071595e-35
			9'd313: out = 16'b0000000000000000; // input=-6.21875, output=2.04704785425e-34
			9'd314: out = 16'b0000000000000000; // input=-6.1875, output=4.44504196183e-34
			9'd315: out = 16'b0000000000000000; // input=-6.15625, output=9.61451258101e-34
			9'd316: out = 16'b0000000000000000; // input=-6.125, output=2.07148701924e-33
			9'd317: out = 16'b0000000000000000; // input=-6.09375, output=4.44570557614e-33
			9'd318: out = 16'b0000000000000000; // input=-6.0625, output=9.50391877478e-33
			9'd319: out = 16'b0000000000000000; // input=-6.03125, output=2.02380316897e-32
			9'd320: out = 16'b0000000000000000; // input=-6.0, output=4.29276747133e-32
			9'd321: out = 16'b0000000000000000; // input=-5.96875, output=9.0700565429e-32
			9'd322: out = 16'b0000000000000000; // input=-5.9375, output=1.90891311466e-31
			9'd323: out = 16'b0000000000000000; // input=-5.90625, output=4.00189662571e-31
			9'd324: out = 16'b0000000000000000; // input=-5.875, output=8.35697508909e-31
			9'd325: out = 16'b0000000000000000; // input=-5.84375, output=1.73834465408e-30
			9'd326: out = 16'b0000000000000000; // input=-5.8125, output=3.60185480783e-30
			9'd327: out = 16'b0000000000000000; // input=-5.78125, output=7.43395718253e-30
			9'd328: out = 16'b0000000000000000; // input=-5.75, output=1.52833108232e-29
			9'd329: out = 16'b0000000000000000; // input=-5.71875, output=3.12981287739e-29
			9'd330: out = 16'b0000000000000000; // input=-5.6875, output=6.38444040927e-29
			9'd331: out = 16'b0000000000000000; // input=-5.65625, output=1.29727138784e-28
			9'd332: out = 16'b0000000000000000; // input=-5.625, output=2.62568352123e-28
			9'd333: out = 16'b0000000000000000; // input=-5.59375, output=5.29367719434e-28
			9'd334: out = 16'b0000000000000000; // input=-5.5625, output=1.0631047732e-27
			9'd335: out = 16'b0000000000000000; // input=-5.53125, output=2.12666076412e-27
			9'd336: out = 16'b0000000000000000; // input=-5.5, output=4.23763850702e-27
			9'd337: out = 16'b0000000000000000; // input=-5.46875, output=8.41110648574e-27
			9'd338: out = 16'b0000000000000000; // input=-5.4375, output=1.66297566216e-26
			9'd339: out = 16'b0000000000000000; // input=-5.40625, output=3.27508210893e-26
			9'd340: out = 16'b0000000000000000; // input=-5.375, output=6.42483574324e-26
			9'd341: out = 16'b0000000000000000; // input=-5.34375, output=1.25546729163e-25
			9'd342: out = 16'b0000000000000000; // input=-5.3125, output=2.4437248966e-25
			9'd343: out = 16'b0000000000000000; // input=-5.28125, output=4.73808405983e-25
			9'd344: out = 16'b0000000000000000; // input=-5.25, output=9.15075118104e-25
			9'd345: out = 16'b0000000000000000; // input=-5.21875, output=1.76041179165e-24
			9'd346: out = 16'b0000000000000000; // input=-5.1875, output=3.37345816254e-24
			9'd347: out = 16'b0000000000000000; // input=-5.15625, output=6.43931877481e-24
			9'd348: out = 16'b0000000000000000; // input=-5.125, output=1.22435697305e-23
			9'd349: out = 16'b0000000000000000; // input=-5.09375, output=2.31888776995e-23
			9'd350: out = 16'b0000000000000000; // input=-5.0625, output=4.37476710924e-23
			9'd351: out = 16'b0000000000000000; // input=-5.03125, output=8.22117104008e-23
			9'd352: out = 16'b0000000000000000; // input=-5.0, output=1.53891972534e-22
			9'd353: out = 16'b0000000000000000; // input=-4.96875, output=2.86947064418e-22
			9'd354: out = 16'b0000000000000000; // input=-4.9375, output=5.32955738878e-22
			9'd355: out = 16'b0000000000000000; // input=-4.90625, output=9.86016170148e-22
			9'd356: out = 16'b0000000000000000; // input=-4.875, output=1.8171068624e-21
			9'd357: out = 16'b0000000000000000; // input=-4.84375, output=3.33564970748e-21
			9'd358: out = 16'b0000000000000000; // input=-4.8125, output=6.09935544127e-21
			9'd359: out = 16'b0000000000000000; // input=-4.78125, output=1.11094097589e-20
			9'd360: out = 16'b0000000000000000; // input=-4.75, output=2.01558707886e-20
			9'd361: out = 16'b0000000000000000; // input=-4.71875, output=3.64263522358e-20
			9'd362: out = 16'b0000000000000000; // input=-4.6875, output=6.55742507756e-20
			9'd363: out = 16'b0000000000000000; // input=-4.65625, output=1.17585705385e-19
			9'd364: out = 16'b0000000000000000; // input=-4.625, output=2.10028996599e-19
			9'd365: out = 16'b0000000000000000; // input=-4.59375, output=3.73686598887e-19
			9'd366: out = 16'b0000000000000000; // input=-4.5625, output=6.62276472038e-19
			9'd367: out = 16'b0000000000000000; // input=-4.53125, output=1.1691619338e-18
			9'd368: out = 16'b0000000000000000; // input=-4.5, output=2.05595471433e-18
			9'd369: out = 16'b0000000000000000; // input=-4.46875, output=3.6012722876e-18
			9'd370: out = 16'b0000000000000000; // input=-4.4375, output=6.28350421733e-18
			9'd371: out = 16'b0000000000000000; // input=-4.40625, output=1.09207232111e-17
			9'd372: out = 16'b0000000000000000; // input=-4.375, output=1.89062077638e-17
			9'd373: out = 16'b0000000000000000; // input=-4.34375, output=3.26032571594e-17
			9'd374: out = 16'b0000000000000000; // input=-4.3125, output=5.6004263471e-17
			9'd375: out = 16'b0000000000000000; // input=-4.28125, output=9.58263017897e-17
			9'd376: out = 16'b0000000000000000; // input=-4.25, output=1.63324712633e-16
			9'd377: out = 16'b0000000000000000; // input=-4.21875, output=2.77282598204e-16
			9'd378: out = 16'b0000000000000000; // input=-4.1875, output=4.68917956941e-16
			9'd379: out = 16'b0000000000000000; // input=-4.15625, output=7.89904613881e-16
			9'd380: out = 16'b0000000000000000; // input=-4.125, output=1.32542749119e-15
			9'd381: out = 16'b0000000000000000; // input=-4.09375, output=2.21534227444e-15
			9'd382: out = 16'b0000000000000000; // input=-4.0625, output=3.68832543083e-15
			9'd383: out = 16'b0000000000000000; // input=-4.03125, output=6.11675616292e-15
			9'd384: out = 16'b0000000000000000; // input=-4.0, output=1.01045421671e-14
			9'd385: out = 16'b0000000000000000; // input=-3.96875, output=1.66270671268e-14
			9'd386: out = 16'b0000000000000000; // input=-3.9375, output=2.72532435195e-14
			9'd387: out = 16'b0000000000000000; // input=-3.90625, output=4.44963390508e-14
			9'd388: out = 16'b0000000000000000; // input=-3.875, output=7.23658890223e-14
			9'd389: out = 16'b0000000000000000; // input=-3.84375, output=1.17232239136e-13
			9'd390: out = 16'b0000000000000000; // input=-3.8125, output=1.89175005616e-13
			9'd391: out = 16'b0000000000000000; // input=-3.78125, output=3.04077291445e-13
			9'd392: out = 16'b0000000000000000; // input=-3.75, output=4.86864106606e-13
			9'd393: out = 16'b0000000000000000; // input=-3.71875, output=7.76488565871e-13
			9'd394: out = 16'b0000000000000000; // input=-3.6875, output=1.23357599371e-12
			9'd395: out = 16'b0000000000000000; // input=-3.65625, output=1.95209203954e-12
			9'd396: out = 16'b0000000000000000; // input=-3.625, output=3.07707590112e-12
			9'd397: out = 16'b0000000000000000; // input=-3.59375, output=4.83147419902e-12
			9'd398: out = 16'b0000000000000000; // input=-3.5625, output=7.55656909133e-12
			9'd399: out = 16'b0000000000000000; // input=-3.53125, output=1.17726216712e-11
			9'd400: out = 16'b0000000000000000; // input=-3.5, output=1.82694408167e-11
			9'd401: out = 16'b0000000000000000; // input=-3.46875, output=2.82410512722e-11
			9'd402: out = 16'b0000000000000000; // input=-3.4375, output=4.34850527144e-11
			9'd403: out = 16'b0000000000000000; // input=-3.40625, output=6.66964440085e-11
			9'd404: out = 16'b0000000000000000; // input=-3.375, output=1.01898759177e-10
			9'd405: out = 16'b0000000000000000; // input=-3.34375, output=1.55073878412e-10
			9'd406: out = 16'b0000000000000000; // input=-3.3125, output=2.35077973981e-10
			9'd407: out = 16'b0000000000000000; // input=-3.28125, output=3.54967642802e-10
			9'd408: out = 16'b0000000000000000; // input=-3.25, output=5.33911322953e-10
			9'd409: out = 16'b0000000000000000; // input=-3.21875, output=7.99931931389e-10
			9'd410: out = 16'b0000000000000000; // input=-3.1875, output=1.19382445829e-09
			9'd411: out = 16'b0000000000000000; // input=-3.15625, output=1.77472655813e-09
			9'd412: out = 16'b0000000000000000; // input=-3.125, output=2.62800363631e-09
			9'd413: out = 16'b0000000000000000; // input=-3.09375, output=3.87635918724e-09
			9'd414: out = 16'b0000000000000000; // input=-3.0625, output=5.69541795659e-09
			9'd415: out = 16'b0000000000000000; // input=-3.03125, output=8.33548213617e-09
			9'd416: out = 16'b0000000000000000; // input=-3.0, output=1.21517656996e-08
			9'd417: out = 16'b0000000000000000; // input=-2.96875, output=1.76462158208e-08
			9'd418: out = 16'b0000000000000000; // input=-2.9375, output=2.55250924071e-08
			9'd419: out = 16'b0000000000000000; // input=-2.90625, output=3.67778719754e-08
			9'd420: out = 16'b0000000000000000; // input=-2.875, output=5.27848640714e-08
			9'd421: out = 16'b0000000000000000; // input=-2.84375, output=7.54632935059e-08
			9'd422: out = 16'b0000000000000000; // input=-2.8125, output=1.07464653011e-07
			9'd423: out = 16'b0000000000000000; // input=-2.78125, output=1.52440043186e-07
			9'd424: out = 16'b0000000000000000; // input=-2.75, output=2.15395200851e-07
			9'd425: out = 16'b0000000000000000; // input=-2.71875, output=3.03163225748e-07
			9'd426: out = 16'b0000000000000000; // input=-2.6875, output=4.25030947662e-07
			9'd427: out = 16'b0000000000000000; // input=-2.65625, output=5.93564781242e-07
			9'd428: out = 16'b0000000000000000; // input=-2.625, output=8.25694197726e-07
			9'd429: out = 16'b0000000000000000; // input=-2.59375, output=1.14412606129e-06
			9'd430: out = 16'b0000000000000000; // input=-2.5625, output=1.57918154814e-06
			9'd431: out = 16'b0000000000000000; // input=-2.53125, output=2.17116975587e-06
			9'd432: out = 16'b0000000000000000; // input=-2.5, output=2.97343902947e-06
			9'd433: out = 16'b0000000000000000; // input=-2.46875, output=4.05627911931e-06
			9'd434: out = 16'b0000000000000000; // input=-2.4375, output=5.5118851951e-06
			9'd435: out = 16'b0000000000000000; // input=-2.40625, output=7.46063909651e-06
			9'd436: out = 16'b0000000000000000; // input=-2.375, output=1.00590145772e-05
			9'd437: out = 16'b0000000000000000; // input=-2.34375, output=1.35094721523e-05
			9'd438: out = 16'b0000000000000000; // input=-2.3125, output=1.80727757781e-05
			9'd439: out = 16'b0000000000000000; // input=-2.28125, output=2.40832380116e-05
			9'd440: out = 16'b0000000000000000; // input=-2.25, output=3.19674822138e-05
			9'd441: out = 16'b0000000000000000; // input=-2.21875, output=4.22673990269e-05
			9'd442: out = 16'b0000000000000000; // input=-2.1875, output=5.56680684584e-05
			9'd443: out = 16'b0000000000000000; // input=-2.15625, output=7.30315164609e-05
			9'd444: out = 16'b0000000000000000; // input=-2.125, output=9.54372730824e-05
			9'd445: out = 16'b0000000000000000; // input=-2.09375, output=0.000124230794341
			9'd446: out = 16'b0000000000000000; // input=-2.0625, output=0.000161080897111
			9'd447: out = 16'b0000000000000000; // input=-2.03125, output=0.000208047429535
			9'd448: out = 16'b0000000000000000; // input=-2.0, output=0.00026766045153
			9'd449: out = 16'b0000000000000000; // input=-1.96875, output=0.000343012222389
			9'd450: out = 16'b0000000000000000; // input=-1.9375, output=0.000437863275529
			9'd451: out = 16'b0000000000000000; // input=-1.90625, output=0.000556763793197
			9'd452: out = 16'b0000000000000000; // input=-1.875, output=0.000705191364735
			9'd453: out = 16'b0000000000000000; // input=-1.84375, output=0.000889706008226
			9'd454: out = 16'b0000000000000000; // input=-1.8125, output=0.00111812304446
			9'd455: out = 16'b0000000000000000; // input=-1.78125, output=0.00139970402189
			9'd456: out = 16'b0000000000000000; // input=-1.75, output=0.00174536539009
			9'd457: out = 16'b0000000000000000; // input=-1.71875, output=0.00216790399823
			9'd458: out = 16'b0000000000000000; // input=-1.6875, output=0.00268223774698
			9'd459: out = 16'b0000000000000000; // input=-1.65625, output=0.00330565884481
			9'd460: out = 16'b0000000000000001; // input=-1.625, output=0.0040580961146
			9'd461: out = 16'b0000000000000001; // input=-1.59375, output=0.00496238167221
			9'd462: out = 16'b0000000000000001; // input=-1.5625, output=0.0060445160704
			9'd463: out = 16'b0000000000000001; // input=-1.53125, output=0.00733392469259
			9'd464: out = 16'b0000000000000001; // input=-1.5, output=0.00886369682388
			9'd465: out = 16'b0000000000000001; // input=-1.46875, output=0.0106707974632
			9'd466: out = 16'b0000000000000010; // input=-1.4375, output=0.0127962406214
			9'd467: out = 16'b0000000000000010; // input=-1.40625, output=0.0152852116375
			9'd468: out = 16'b0000000000000010; // input=-1.375, output=0.0181871250032
			9'd469: out = 16'b0000000000000011; // input=-1.34375, output=0.0215556034005
			9'd470: out = 16'b0000000000000011; // input=-1.3125, output=0.0254483631937
			9'd471: out = 16'b0000000000000100; // input=-1.28125, output=0.0299269915718
			9'd472: out = 16'b0000000000000100; // input=-1.25, output=0.0350566009871
			9'd473: out = 16'b0000000000000101; // input=-1.21875, output=0.0409053475456
			9'd474: out = 16'b0000000000000110; // input=-1.1875, output=0.0475438016598
			9'd475: out = 16'b0000000000000111; // input=-1.15625, output=0.0550441616058
			9'd476: out = 16'b0000000000001000; // input=-1.125, output=0.0634793036713
			9'd477: out = 16'b0000000000001001; // input=-1.09375, output=0.0729216663524
			9'd478: out = 16'b0000000000001011; // input=-1.0625, output=0.0834419705127
			9'd479: out = 16'b0000000000001100; // input=-1.03125, output=0.0951077825213
			9'd480: out = 16'b0000000000001110; // input=-1.0, output=0.107981933026
			9'd481: out = 16'b0000000000010000; // input=-0.96875, output=0.122120810082
			9'd482: out = 16'b0000000000010010; // input=-0.9375, output=0.137572551653
			9'd483: out = 16'b0000000000010100; // input=-0.90625, output=0.154375168879
			9'd484: out = 16'b0000000000010110; // input=-0.875, output=0.172554637653
			9'd485: out = 16'b0000000000011001; // input=-0.84375, output=0.19212300181
			9'd486: out = 16'b0000000000011011; // input=-0.8125, output=0.213076536261
			9'd487: out = 16'b0000000000011110; // input=-0.78125, output=0.235394022449
			9'd488: out = 16'b0000000000100001; // input=-0.75, output=0.259035191332
			9'd489: out = 16'b0000000000100100; // input=-0.71875, output=0.28393939041
			9'd490: out = 16'b0000000000101000; // input=-0.6875, output=0.310024530917
			9'd491: out = 16'b0000000000101011; // input=-0.65625, output=0.337186369036
			9'd492: out = 16'b0000000000101111; // input=-0.625, output=0.365298170778
			9'd493: out = 16'b0000000000110010; // input=-0.59375, output=0.394210803837
			9'd494: out = 16'b0000000000110110; // input=-0.5625, output=0.423753291551
			9'd495: out = 16'b0000000000111010; // input=-0.53125, output=0.453733853938
			9'd496: out = 16'b0000000000111110; // input=-0.5, output=0.483941449038
			9'd497: out = 16'b0000000001000010; // input=-0.46875, output=0.514147814693
			9'd498: out = 16'b0000000001000110; // input=-0.4375, output=0.544109996757
			9'd499: out = 16'b0000000001001001; // input=-0.40625, output=0.573573335133
			9'd500: out = 16'b0000000001001101; // input=-0.375, output=0.60227486431
			9'd501: out = 16'b0000000001010001; // input=-0.34375, output=0.629947070853
			9'd502: out = 16'b0000000001010100; // input=-0.3125, output=0.656321937101
			9'd503: out = 16'b0000000001010111; // input=-0.28125, output=0.68113518864
			9'd504: out = 16'b0000000001011010; // input=-0.25, output=0.704130653529
			9'd505: out = 16'b0000000001011101; // input=-0.21875, output=0.725064634081
			9'd506: out = 16'b0000000001011111; // input=-0.1875, output=0.74371018774
			9'd507: out = 16'b0000000001100001; // input=-0.15625, output=0.759861212397
			9'd508: out = 16'b0000000001100011; // input=-0.125, output=0.773336233606
			9'd509: out = 16'b0000000001100100; // input=-0.09375, output=0.783981796505
			9'd510: out = 16'b0000000001100101; // input=-0.0625, output=0.791675373889
			9'd511: out = 16'b0000000001100110; // input=-0.03125, output=0.796327713374
			9'd0: out = 16'b0000000001100110; // input=0.0, output=0.797884560803
			9'd1: out = 16'b0000000001100110; // input=0.03125, output=0.796327713374
			9'd2: out = 16'b0000000001100101; // input=0.0625, output=0.791675373889
			9'd3: out = 16'b0000000001100100; // input=0.09375, output=0.783981796505
			9'd4: out = 16'b0000000001100011; // input=0.125, output=0.773336233606
			9'd5: out = 16'b0000000001100001; // input=0.15625, output=0.759861212397
			9'd6: out = 16'b0000000001011111; // input=0.1875, output=0.74371018774
			9'd7: out = 16'b0000000001011101; // input=0.21875, output=0.725064634081
			9'd8: out = 16'b0000000001011010; // input=0.25, output=0.704130653529
			9'd9: out = 16'b0000000001010111; // input=0.28125, output=0.68113518864
			9'd10: out = 16'b0000000001010100; // input=0.3125, output=0.656321937101
			9'd11: out = 16'b0000000001010001; // input=0.34375, output=0.629947070853
			9'd12: out = 16'b0000000001001101; // input=0.375, output=0.60227486431
			9'd13: out = 16'b0000000001001001; // input=0.40625, output=0.573573335133
			9'd14: out = 16'b0000000001000110; // input=0.4375, output=0.544109996757
			9'd15: out = 16'b0000000001000010; // input=0.46875, output=0.514147814693
			9'd16: out = 16'b0000000000111110; // input=0.5, output=0.483941449038
			9'd17: out = 16'b0000000000111010; // input=0.53125, output=0.453733853938
			9'd18: out = 16'b0000000000110110; // input=0.5625, output=0.423753291551
			9'd19: out = 16'b0000000000110010; // input=0.59375, output=0.394210803837
			9'd20: out = 16'b0000000000101111; // input=0.625, output=0.365298170778
			9'd21: out = 16'b0000000000101011; // input=0.65625, output=0.337186369036
			9'd22: out = 16'b0000000000101000; // input=0.6875, output=0.310024530917
			9'd23: out = 16'b0000000000100100; // input=0.71875, output=0.28393939041
			9'd24: out = 16'b0000000000100001; // input=0.75, output=0.259035191332
			9'd25: out = 16'b0000000000011110; // input=0.78125, output=0.235394022449
			9'd26: out = 16'b0000000000011011; // input=0.8125, output=0.213076536261
			9'd27: out = 16'b0000000000011001; // input=0.84375, output=0.19212300181
			9'd28: out = 16'b0000000000010110; // input=0.875, output=0.172554637653
			9'd29: out = 16'b0000000000010100; // input=0.90625, output=0.154375168879
			9'd30: out = 16'b0000000000010010; // input=0.9375, output=0.137572551653
			9'd31: out = 16'b0000000000010000; // input=0.96875, output=0.122120810082
			9'd32: out = 16'b0000000000001110; // input=1.0, output=0.107981933026
			9'd33: out = 16'b0000000000001100; // input=1.03125, output=0.0951077825213
			9'd34: out = 16'b0000000000001011; // input=1.0625, output=0.0834419705127
			9'd35: out = 16'b0000000000001001; // input=1.09375, output=0.0729216663524
			9'd36: out = 16'b0000000000001000; // input=1.125, output=0.0634793036713
			9'd37: out = 16'b0000000000000111; // input=1.15625, output=0.0550441616058
			9'd38: out = 16'b0000000000000110; // input=1.1875, output=0.0475438016598
			9'd39: out = 16'b0000000000000101; // input=1.21875, output=0.0409053475456
			9'd40: out = 16'b0000000000000100; // input=1.25, output=0.0350566009871
			9'd41: out = 16'b0000000000000100; // input=1.28125, output=0.0299269915718
			9'd42: out = 16'b0000000000000011; // input=1.3125, output=0.0254483631937
			9'd43: out = 16'b0000000000000011; // input=1.34375, output=0.0215556034005
			9'd44: out = 16'b0000000000000010; // input=1.375, output=0.0181871250032
			9'd45: out = 16'b0000000000000010; // input=1.40625, output=0.0152852116375
			9'd46: out = 16'b0000000000000010; // input=1.4375, output=0.0127962406214
			9'd47: out = 16'b0000000000000001; // input=1.46875, output=0.0106707974632
			9'd48: out = 16'b0000000000000001; // input=1.5, output=0.00886369682388
			9'd49: out = 16'b0000000000000001; // input=1.53125, output=0.00733392469259
			9'd50: out = 16'b0000000000000001; // input=1.5625, output=0.0060445160704
			9'd51: out = 16'b0000000000000001; // input=1.59375, output=0.00496238167221
			9'd52: out = 16'b0000000000000001; // input=1.625, output=0.0040580961146
			9'd53: out = 16'b0000000000000000; // input=1.65625, output=0.00330565884481
			9'd54: out = 16'b0000000000000000; // input=1.6875, output=0.00268223774698
			9'd55: out = 16'b0000000000000000; // input=1.71875, output=0.00216790399823
			9'd56: out = 16'b0000000000000000; // input=1.75, output=0.00174536539009
			9'd57: out = 16'b0000000000000000; // input=1.78125, output=0.00139970402189
			9'd58: out = 16'b0000000000000000; // input=1.8125, output=0.00111812304446
			9'd59: out = 16'b0000000000000000; // input=1.84375, output=0.000889706008226
			9'd60: out = 16'b0000000000000000; // input=1.875, output=0.000705191364735
			9'd61: out = 16'b0000000000000000; // input=1.90625, output=0.000556763793197
			9'd62: out = 16'b0000000000000000; // input=1.9375, output=0.000437863275529
			9'd63: out = 16'b0000000000000000; // input=1.96875, output=0.000343012222389
			9'd64: out = 16'b0000000000000000; // input=2.0, output=0.00026766045153
			9'd65: out = 16'b0000000000000000; // input=2.03125, output=0.000208047429535
			9'd66: out = 16'b0000000000000000; // input=2.0625, output=0.000161080897111
			9'd67: out = 16'b0000000000000000; // input=2.09375, output=0.000124230794341
			9'd68: out = 16'b0000000000000000; // input=2.125, output=9.54372730824e-05
			9'd69: out = 16'b0000000000000000; // input=2.15625, output=7.30315164609e-05
			9'd70: out = 16'b0000000000000000; // input=2.1875, output=5.56680684584e-05
			9'd71: out = 16'b0000000000000000; // input=2.21875, output=4.22673990269e-05
			9'd72: out = 16'b0000000000000000; // input=2.25, output=3.19674822138e-05
			9'd73: out = 16'b0000000000000000; // input=2.28125, output=2.40832380116e-05
			9'd74: out = 16'b0000000000000000; // input=2.3125, output=1.80727757781e-05
			9'd75: out = 16'b0000000000000000; // input=2.34375, output=1.35094721523e-05
			9'd76: out = 16'b0000000000000000; // input=2.375, output=1.00590145772e-05
			9'd77: out = 16'b0000000000000000; // input=2.40625, output=7.46063909651e-06
			9'd78: out = 16'b0000000000000000; // input=2.4375, output=5.5118851951e-06
			9'd79: out = 16'b0000000000000000; // input=2.46875, output=4.05627911931e-06
			9'd80: out = 16'b0000000000000000; // input=2.5, output=2.97343902947e-06
			9'd81: out = 16'b0000000000000000; // input=2.53125, output=2.17116975587e-06
			9'd82: out = 16'b0000000000000000; // input=2.5625, output=1.57918154814e-06
			9'd83: out = 16'b0000000000000000; // input=2.59375, output=1.14412606129e-06
			9'd84: out = 16'b0000000000000000; // input=2.625, output=8.25694197726e-07
			9'd85: out = 16'b0000000000000000; // input=2.65625, output=5.93564781242e-07
			9'd86: out = 16'b0000000000000000; // input=2.6875, output=4.25030947662e-07
			9'd87: out = 16'b0000000000000000; // input=2.71875, output=3.03163225748e-07
			9'd88: out = 16'b0000000000000000; // input=2.75, output=2.15395200851e-07
			9'd89: out = 16'b0000000000000000; // input=2.78125, output=1.52440043186e-07
			9'd90: out = 16'b0000000000000000; // input=2.8125, output=1.07464653011e-07
			9'd91: out = 16'b0000000000000000; // input=2.84375, output=7.54632935059e-08
			9'd92: out = 16'b0000000000000000; // input=2.875, output=5.27848640714e-08
			9'd93: out = 16'b0000000000000000; // input=2.90625, output=3.67778719754e-08
			9'd94: out = 16'b0000000000000000; // input=2.9375, output=2.55250924071e-08
			9'd95: out = 16'b0000000000000000; // input=2.96875, output=1.76462158208e-08
			9'd96: out = 16'b0000000000000000; // input=3.0, output=1.21517656996e-08
			9'd97: out = 16'b0000000000000000; // input=3.03125, output=8.33548213617e-09
			9'd98: out = 16'b0000000000000000; // input=3.0625, output=5.69541795659e-09
			9'd99: out = 16'b0000000000000000; // input=3.09375, output=3.87635918724e-09
			9'd100: out = 16'b0000000000000000; // input=3.125, output=2.62800363631e-09
			9'd101: out = 16'b0000000000000000; // input=3.15625, output=1.77472655813e-09
			9'd102: out = 16'b0000000000000000; // input=3.1875, output=1.19382445829e-09
			9'd103: out = 16'b0000000000000000; // input=3.21875, output=7.99931931389e-10
			9'd104: out = 16'b0000000000000000; // input=3.25, output=5.33911322953e-10
			9'd105: out = 16'b0000000000000000; // input=3.28125, output=3.54967642802e-10
			9'd106: out = 16'b0000000000000000; // input=3.3125, output=2.35077973981e-10
			9'd107: out = 16'b0000000000000000; // input=3.34375, output=1.55073878412e-10
			9'd108: out = 16'b0000000000000000; // input=3.375, output=1.01898759177e-10
			9'd109: out = 16'b0000000000000000; // input=3.40625, output=6.66964440085e-11
			9'd110: out = 16'b0000000000000000; // input=3.4375, output=4.34850527144e-11
			9'd111: out = 16'b0000000000000000; // input=3.46875, output=2.82410512722e-11
			9'd112: out = 16'b0000000000000000; // input=3.5, output=1.82694408167e-11
			9'd113: out = 16'b0000000000000000; // input=3.53125, output=1.17726216712e-11
			9'd114: out = 16'b0000000000000000; // input=3.5625, output=7.55656909133e-12
			9'd115: out = 16'b0000000000000000; // input=3.59375, output=4.83147419902e-12
			9'd116: out = 16'b0000000000000000; // input=3.625, output=3.07707590112e-12
			9'd117: out = 16'b0000000000000000; // input=3.65625, output=1.95209203954e-12
			9'd118: out = 16'b0000000000000000; // input=3.6875, output=1.23357599371e-12
			9'd119: out = 16'b0000000000000000; // input=3.71875, output=7.76488565871e-13
			9'd120: out = 16'b0000000000000000; // input=3.75, output=4.86864106606e-13
			9'd121: out = 16'b0000000000000000; // input=3.78125, output=3.04077291445e-13
			9'd122: out = 16'b0000000000000000; // input=3.8125, output=1.89175005616e-13
			9'd123: out = 16'b0000000000000000; // input=3.84375, output=1.17232239136e-13
			9'd124: out = 16'b0000000000000000; // input=3.875, output=7.23658890223e-14
			9'd125: out = 16'b0000000000000000; // input=3.90625, output=4.44963390508e-14
			9'd126: out = 16'b0000000000000000; // input=3.9375, output=2.72532435195e-14
			9'd127: out = 16'b0000000000000000; // input=3.96875, output=1.66270671268e-14
			9'd128: out = 16'b0000000000000000; // input=4.0, output=1.01045421671e-14
			9'd129: out = 16'b0000000000000000; // input=4.03125, output=6.11675616292e-15
			9'd130: out = 16'b0000000000000000; // input=4.0625, output=3.68832543083e-15
			9'd131: out = 16'b0000000000000000; // input=4.09375, output=2.21534227444e-15
			9'd132: out = 16'b0000000000000000; // input=4.125, output=1.32542749119e-15
			9'd133: out = 16'b0000000000000000; // input=4.15625, output=7.89904613881e-16
			9'd134: out = 16'b0000000000000000; // input=4.1875, output=4.68917956941e-16
			9'd135: out = 16'b0000000000000000; // input=4.21875, output=2.77282598204e-16
			9'd136: out = 16'b0000000000000000; // input=4.25, output=1.63324712633e-16
			9'd137: out = 16'b0000000000000000; // input=4.28125, output=9.58263017897e-17
			9'd138: out = 16'b0000000000000000; // input=4.3125, output=5.6004263471e-17
			9'd139: out = 16'b0000000000000000; // input=4.34375, output=3.26032571594e-17
			9'd140: out = 16'b0000000000000000; // input=4.375, output=1.89062077638e-17
			9'd141: out = 16'b0000000000000000; // input=4.40625, output=1.09207232111e-17
			9'd142: out = 16'b0000000000000000; // input=4.4375, output=6.28350421733e-18
			9'd143: out = 16'b0000000000000000; // input=4.46875, output=3.6012722876e-18
			9'd144: out = 16'b0000000000000000; // input=4.5, output=2.05595471433e-18
			9'd145: out = 16'b0000000000000000; // input=4.53125, output=1.1691619338e-18
			9'd146: out = 16'b0000000000000000; // input=4.5625, output=6.62276472038e-19
			9'd147: out = 16'b0000000000000000; // input=4.59375, output=3.73686598887e-19
			9'd148: out = 16'b0000000000000000; // input=4.625, output=2.10028996599e-19
			9'd149: out = 16'b0000000000000000; // input=4.65625, output=1.17585705385e-19
			9'd150: out = 16'b0000000000000000; // input=4.6875, output=6.55742507756e-20
			9'd151: out = 16'b0000000000000000; // input=4.71875, output=3.64263522358e-20
			9'd152: out = 16'b0000000000000000; // input=4.75, output=2.01558707886e-20
			9'd153: out = 16'b0000000000000000; // input=4.78125, output=1.11094097589e-20
			9'd154: out = 16'b0000000000000000; // input=4.8125, output=6.09935544127e-21
			9'd155: out = 16'b0000000000000000; // input=4.84375, output=3.33564970748e-21
			9'd156: out = 16'b0000000000000000; // input=4.875, output=1.8171068624e-21
			9'd157: out = 16'b0000000000000000; // input=4.90625, output=9.86016170148e-22
			9'd158: out = 16'b0000000000000000; // input=4.9375, output=5.32955738878e-22
			9'd159: out = 16'b0000000000000000; // input=4.96875, output=2.86947064418e-22
			9'd160: out = 16'b0000000000000000; // input=5.0, output=1.53891972534e-22
			9'd161: out = 16'b0000000000000000; // input=5.03125, output=8.22117104008e-23
			9'd162: out = 16'b0000000000000000; // input=5.0625, output=4.37476710924e-23
			9'd163: out = 16'b0000000000000000; // input=5.09375, output=2.31888776995e-23
			9'd164: out = 16'b0000000000000000; // input=5.125, output=1.22435697305e-23
			9'd165: out = 16'b0000000000000000; // input=5.15625, output=6.43931877481e-24
			9'd166: out = 16'b0000000000000000; // input=5.1875, output=3.37345816254e-24
			9'd167: out = 16'b0000000000000000; // input=5.21875, output=1.76041179165e-24
			9'd168: out = 16'b0000000000000000; // input=5.25, output=9.15075118104e-25
			9'd169: out = 16'b0000000000000000; // input=5.28125, output=4.73808405983e-25
			9'd170: out = 16'b0000000000000000; // input=5.3125, output=2.4437248966e-25
			9'd171: out = 16'b0000000000000000; // input=5.34375, output=1.25546729163e-25
			9'd172: out = 16'b0000000000000000; // input=5.375, output=6.42483574324e-26
			9'd173: out = 16'b0000000000000000; // input=5.40625, output=3.27508210893e-26
			9'd174: out = 16'b0000000000000000; // input=5.4375, output=1.66297566216e-26
			9'd175: out = 16'b0000000000000000; // input=5.46875, output=8.41110648574e-27
			9'd176: out = 16'b0000000000000000; // input=5.5, output=4.23763850702e-27
			9'd177: out = 16'b0000000000000000; // input=5.53125, output=2.12666076412e-27
			9'd178: out = 16'b0000000000000000; // input=5.5625, output=1.0631047732e-27
			9'd179: out = 16'b0000000000000000; // input=5.59375, output=5.29367719434e-28
			9'd180: out = 16'b0000000000000000; // input=5.625, output=2.62568352123e-28
			9'd181: out = 16'b0000000000000000; // input=5.65625, output=1.29727138784e-28
			9'd182: out = 16'b0000000000000000; // input=5.6875, output=6.38444040927e-29
			9'd183: out = 16'b0000000000000000; // input=5.71875, output=3.12981287739e-29
			9'd184: out = 16'b0000000000000000; // input=5.75, output=1.52833108232e-29
			9'd185: out = 16'b0000000000000000; // input=5.78125, output=7.43395718253e-30
			9'd186: out = 16'b0000000000000000; // input=5.8125, output=3.60185480783e-30
			9'd187: out = 16'b0000000000000000; // input=5.84375, output=1.73834465408e-30
			9'd188: out = 16'b0000000000000000; // input=5.875, output=8.35697508909e-31
			9'd189: out = 16'b0000000000000000; // input=5.90625, output=4.00189662571e-31
			9'd190: out = 16'b0000000000000000; // input=5.9375, output=1.90891311466e-31
			9'd191: out = 16'b0000000000000000; // input=5.96875, output=9.0700565429e-32
			9'd192: out = 16'b0000000000000000; // input=6.0, output=4.29276747133e-32
			9'd193: out = 16'b0000000000000000; // input=6.03125, output=2.02380316897e-32
			9'd194: out = 16'b0000000000000000; // input=6.0625, output=9.50391877478e-33
			9'd195: out = 16'b0000000000000000; // input=6.09375, output=4.44570557614e-33
			9'd196: out = 16'b0000000000000000; // input=6.125, output=2.07148701924e-33
			9'd197: out = 16'b0000000000000000; // input=6.15625, output=9.61451258101e-34
			9'd198: out = 16'b0000000000000000; // input=6.1875, output=4.44504196183e-34
			9'd199: out = 16'b0000000000000000; // input=6.21875, output=2.04704785425e-34
			9'd200: out = 16'b0000000000000000; // input=6.25, output=9.39039071595e-35
			9'd201: out = 16'b0000000000000000; // input=6.28125, output=4.29084540294e-35
			9'd202: out = 16'b0000000000000000; // input=6.3125, output=1.9530151363e-35
			9'd203: out = 16'b0000000000000000; // input=6.34375, output=8.85465996484e-36
			9'd204: out = 16'b0000000000000000; // input=6.375, output=3.99891068444e-36
			9'd205: out = 16'b0000000000000000; // input=6.40625, output=1.79893328563e-36
			9'd206: out = 16'b0000000000000000; // input=6.4375, output=8.06105618402e-37
			9'd207: out = 16'b0000000000000000; // input=6.46875, output=3.59809292893e-37
			9'd208: out = 16'b0000000000000000; // input=6.5, output=1.5997655514e-37
			9'd209: out = 16'b0000000000000000; // input=6.53125, output=7.08506506176e-38
			9'd210: out = 16'b0000000000000000; // input=6.5625, output=3.12561067823e-38
			9'd211: out = 16'b0000000000000000; // input=6.59375, output=1.37350251292e-38
			9'd212: out = 16'b0000000000000000; // input=6.625, output=6.0121190522e-39
			9'd213: out = 16'b0000000000000000; // input=6.65625, output=2.62137541904e-39
			9'd214: out = 16'b0000000000000000; // input=6.6875, output=1.13850360632e-39
			9'd215: out = 16'b0000000000000000; // input=6.71875, output=4.92541848268e-40
			9'd216: out = 16'b0000000000000000; // input=6.75, output=2.12253762783e-40
			9'd217: out = 16'b0000000000000000; // input=6.78125, output=9.11110806056e-41
			9'd218: out = 16'b0000000000000000; // input=6.8125, output=3.89574510993e-41
			9'd219: out = 16'b0000000000000000; // input=6.84375, output=1.65925604311e-41
			9'd220: out = 16'b0000000000000000; // input=6.875, output=7.03946767599e-42
			9'd221: out = 16'b0000000000000000; // input=6.90625, output=2.97488215993e-42
			9'd222: out = 16'b0000000000000000; // input=6.9375, output=1.25228521358e-42
			9'd223: out = 16'b0000000000000000; // input=6.96875, output=5.25097892486e-43
			9'd224: out = 16'b0000000000000000; // input=7.0, output=2.19321311878e-43
			9'd225: out = 16'b0000000000000000; // input=7.03125, output=9.12483314748e-44
			9'd226: out = 16'b0000000000000000; // input=7.0625, output=3.78157367485e-44
			9'd227: out = 16'b0000000000000000; // input=7.09375, output=1.56107488696e-44
			9'd228: out = 16'b0000000000000000; // input=7.125, output=6.41916362084e-45
			9'd229: out = 16'b0000000000000000; // input=7.15625, output=2.62927911298e-45
			9'd230: out = 16'b0000000000000000; // input=7.1875, output=1.07274987899e-45
			9'd231: out = 16'b0000000000000000; // input=7.21875, output=4.35977216421e-46
			9'd232: out = 16'b0000000000000000; // input=7.25, output=1.76495099492e-46
			9'd233: out = 16'b0000000000000000; // input=7.28125, output=7.1171324113e-47
			9'd234: out = 16'b0000000000000000; // input=7.3125, output=2.85878159428e-47
			9'd235: out = 16'b0000000000000000; // input=7.34375, output=1.14382726918e-47
			9'd236: out = 16'b0000000000000000; // input=7.375, output=4.55872560131e-48
			9'd237: out = 16'b0000000000000000; // input=7.40625, output=1.80979754616e-48
			9'd238: out = 16'b0000000000000000; // input=7.4375, output=7.15681968385e-49
			9'd239: out = 16'b0000000000000000; // input=7.46875, output=2.81912084447e-49
			9'd240: out = 16'b0000000000000000; // input=7.5, output=1.10614190997e-49
			9'd241: out = 16'b0000000000000000; // input=7.53125, output=4.32326183636e-50
			9'd242: out = 16'b0000000000000000; // input=7.5625, output=1.68312266462e-50
			9'd243: out = 16'b0000000000000000; // input=7.59375, output=6.52714911362e-51
			9'd244: out = 16'b0000000000000000; // input=7.625, output=2.52135987788e-51
			9'd245: out = 16'b0000000000000000; // input=7.65625, output=9.70174103983e-52
			9'd246: out = 16'b0000000000000000; // input=7.6875, output=3.71850231248e-52
			9'd247: out = 16'b0000000000000000; // input=7.71875, output=1.41967838716e-52
			9'd248: out = 16'b0000000000000000; // input=7.75, output=5.39902604918e-53
			9'd249: out = 16'b0000000000000000; // input=7.78125, output=2.04524063202e-53
			9'd250: out = 16'b0000000000000000; // input=7.8125, output=7.71750533773e-54
			9'd251: out = 16'b0000000000000000; // input=7.84375, output=2.90076804211e-54
			9'd252: out = 16'b0000000000000000; // input=7.875, output=1.0860569595e-54
			9'd253: out = 16'b0000000000000000; // input=7.90625, output=4.05037972923e-55
			9'd254: out = 16'b0000000000000000; // input=7.9375, output=1.50467399787e-55
			9'd255: out = 16'b0000000000000000; // input=7.96875, output=5.56791540596e-56
		endcase
		end
	end
endmodule
