
`timescale 1ns/1ps
module instruction_memory #(
    parameter integer addrLen = 5,
    parameter integer dataLen = 32,
    parameter integer peId  = 1
)(
    input clk,
    input rstn,
    
    input stall,
    input start,
    input restart,
    
    output reg [dataLen - 1: 0] data_out
);
//--------------------------------------------------------------------------------------
//reg [dataLen - 1: 0] mem  [0: (1 << addrLen) - 1];
reg [addrLen-1:0]        address;
reg enable;
reg [dataLen - 1: 0] rdata;
wire end_of_instruction;
always @(posedge clk or negedge rstn)
    if(~rstn)
        enable <= 1'b0;
    else if(start)
        enable <= 1'b1;
    else if(end_of_instruction)
       enable <= 1'b0;
always @(posedge clk or negedge rstn) begin
    if(~rstn)
        address <= {addrLen{1'b0}};
    else begin
        if(end_of_instruction)
            address <= {addrLen{1'b0}};
        else if(~stall && enable )
            address <= address + {{addrLen-1{1'b0}},1'b1};   
    end     
end
always @(posedge clk or negedge rstn) begin
    if(~rstn)
        data_out <= {1'b1,{dataLen-1{1'b0}}};
    else if((~stall && enable && ~end_of_instruction)||(end_of_instruction && start))
       data_out <= rdata;
end
    
assign end_of_instruction = (data_out[dataLen-1:dataLen-5] == 5'b0);
/****************************************************************************/
generate
if(peId == 0) begin
	always @(*) begin
		case(address)
			// PEs: 5 -> 16
			// srcs: (6, 0)(1577) -4 --> (1577) -4:PEGB5, pass, PUGB2
			10'd0 : rdata = 48'b110001110000101000000000000000000000000000001010;
			// PEs: 6 -> 16
			// srcs: (7, 1)(1578) -6 --> (1578) -6:PEGB6, pass, PUGB2
			10'd1 : rdata = 48'b110001110000110000000000000000000000000000001010;
			// PEs: 1 -> 16
			// srcs: (8, 18)(1653) 0 --> (1653) 0:PEGB1, pass, PUGB2
			10'd2 : rdata = 48'b110001110000001000000000000000000000000000001010;
			// PEs: 2 -> 16
			// srcs: (9, 19)(1654) -4 --> (1654) -4:PEGB2, pass, PUGB2
			10'd3 : rdata = 48'b110001110000010000000000000000000000000000001010;
			// PEs: 3 -> 24
			// srcs: (10, 20)(1656) 0 --> (1656) 0:PEGB3, pass, PUGB3
			10'd4 : rdata = 48'b110001110000011000000000000000000000000000001011;
			// PEs: 8 -> 2
			// srcs: (11, 2)(1581) 1 --> (1581) 1:PUGB1, pass, PEGB2
			10'd5 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 0
			// srcs: (12, 3)(1583) -4 --> (1583) -4:PUGB1, pass, NI0
			10'd6 : rdata = 48'b110001110000001100000000000100000000000000000000;
			// PEs: 8 -> 3
			// srcs: (13, 4)(1584) -4 --> (1584) -4:PUGB1, pass, PEGB3
			10'd7 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 0
			// srcs: (14, 6)(1586) -4 --> (1586) -4:PUGB1, pass, NI1
			10'd8 : rdata = 48'b110001110000001100000000000100001000000000000000;
			// PEs: 8 -> 4
			// srcs: (15, 7)(1587) 3 --> (1587) 3:PUGB1, pass, PEGB4
			10'd9 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 0
			// srcs: (16, 9)(1589) 6 --> (1589) 6:PUGB1, pass, NI2
			10'd10 : rdata = 48'b110001110000001100000000000100010000000000000000;
			// PEs: 8 -> 5
			// srcs: (17, 10)(1590) 3 --> (1590) 3:PUGB1, pass, PEGB5
			10'd11 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 16 -> 0
			// srcs: (18, 12)(1592) 9 --> (1592) 9:PUGB2, pass, NI3
			10'd12 : rdata = 48'b110001110000010100000000000100011000000000000000;
			// PEs: 16 -> 6
			// srcs: (19, 13)(1593) -3 --> (1593) -3:PUGB2, pass, PEGB6
			10'd13 : rdata = 48'b110001110000010100000000000000000000000011100000;
			// PEs: 16 -> 0
			// srcs: (20, 15)(1595) 0 --> (1595) 0:PUGB2, pass, NI4
			10'd14 : rdata = 48'b110001110000010100000000000100100000000000000000;
			// PEs: 16 -> 7
			// srcs: (21, 16)(1596) -6 --> (1596) -6:PUGB2, pass, PEGB7
			10'd15 : rdata = 48'b110001110000010100000000000000000000000011110000;
			// PEs: 0 -> 3
			// srcs: (22, 5)(1583) -4 --> (1583) -4:NI0, pass, PEGB3
			10'd16 : rdata = 48'b110001010000000000000000000000000000000010110000;
			// PEs: 4 -> 24
			// srcs: (23, 21)(1657) 1 --> (1657) 1:PEGB4, pass, PUGB3
			10'd17 : rdata = 48'b110001110000100000000000000000000000000000001011;
			// PEs: 0 -> 4
			// srcs: (24, 8)(1586) -4 --> (1586) -4:NI1, pass, PEGB4
			10'd18 : rdata = 48'b110001010000000100000000000000000000000011000000;
			// PEs: 5 -> 32
			// srcs: (25, 22)(1659) 2 --> (1659) 2:PEGB5, pass, PUGB4
			10'd19 : rdata = 48'b110001110000101000000000000000000000000000001100;
			// PEs: 0 -> 5
			// srcs: (26, 11)(1589) 6 --> (1589) 6:NI2, pass, PEGB5
			10'd20 : rdata = 48'b110001010000001000000000000000000000000011010000;
			// PEs: 6 -> 32
			// srcs: (27, 23)(1660) 0 --> (1660) 0:PEGB6, pass, PUGB4
			10'd21 : rdata = 48'b110001110000110000000000000000000000000000001100;
			// PEs: 0 -> 6
			// srcs: (28, 14)(1592) 9 --> (1592) 9:NI3, pass, PEGB6
			10'd22 : rdata = 48'b110001010000001100000000000000000000000011100000;
			// PEs: 56 -> 0
			// srcs: (29, 25)(1724) 2 --> (1724) 2:PUNB, pass, NI0
			10'd23 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 0 -> 7
			// srcs: (30, 17)(1595) 0 --> (1595) 0:NI4, pass, PEGB7
			10'd24 : rdata = 48'b110001010000010000000000000000000000000011110000;
			// PEs: 8 -> 1
			// srcs: (31, 24)(1663) -3 --> (1663) -3:PUGB1, pass, PENB
			10'd25 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 56 -> 2
			// srcs: (32, 26)(1725) 6 --> (1725) 6:PUNB, pass, PEGB2
			10'd26 : rdata = 48'b110001101111111100000000000000000000000010100000;
			// PEs: 56 -> 0
			// srcs: (33, 28)(1727) 0 --> (1727) 0:PUNB, pass, NI1
			10'd27 : rdata = 48'b110001101111111100000000000100001000000000000000;
			// PEs: 56 -> 3
			// srcs: (34, 29)(1728) 6 --> (1728) 6:PUNB, pass, PEGB3
			10'd28 : rdata = 48'b110001101111111100000000000000000000000010110000;
			// PEs: 56 -> 0
			// srcs: (35, 31)(1730) 0 --> (1730) 0:PUNB, pass, NI2
			10'd29 : rdata = 48'b110001101111111100000000000100010000000000000000;
			// PEs: 56 -> 4
			// srcs: (36, 32)(1731) -2 --> (1731) -2:PUNB, pass, PEGB4
			10'd30 : rdata = 48'b110001101111111100000000000000000000000011000000;
			// PEs: 1 -> 8
			// srcs: (37, 34)(1733) 4 --> (1733) 4:PEGB1, pass, PUNB
			10'd31 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 2 -> 8
			// srcs: (38, 35)(1734) -1 --> (1734) -1:PEGB2, pass, PUNB
			10'd32 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 3 -> 8
			// srcs: (39, 36)(1736) -2 --> (1736) -2:PEGB3, pass, PUNB
			10'd33 : rdata = 48'b110001110000011000000000000000000000001000000000;
			// PEs: 4 -> 8
			// srcs: (40, 37)(1737) 0 --> (1737) 0:PEGB4, pass, PUNB
			10'd34 : rdata = 48'b110001110000100000000000000000000000001000000000;
			// PEs: 0 -> 2
			// srcs: (41, 27)(1724) 2 --> (1724) 2:NI0, pass, PEGB2
			10'd35 : rdata = 48'b110001010000000000000000000000000000000010100000;
			// PEs: 5 -> 8
			// srcs: (42, 38)(1739) -1 --> (1739) -1:PEGB5, pass, PUNB
			10'd36 : rdata = 48'b110001110000101000000000000000000000001000000000;
			// PEs: 0 -> 3
			// srcs: (43, 30)(1727) 0 --> (1727) 0:NI1, pass, PEGB3
			10'd37 : rdata = 48'b110001010000000100000000000000000000000010110000;
			// PEs: 6 -> 8
			// srcs: (44, 39)(1740) 0 --> (1740) 0:PEGB6, pass, PUNB
			10'd38 : rdata = 48'b110001110000110000000000000000000000001000000000;
			// PEs: 0 -> 4
			// srcs: (45, 33)(1730) 0 --> (1730) 0:NI2, pass, PEGB4
			10'd39 : rdata = 48'b110001010000001000000000000000000000000011000000;
			// PEs: 8 -> 1
			// srcs: (46, 40)(1743) 1 --> (1743) 1:PUGB1, pass, PENB
			10'd40 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 48 -> 0
			// srcs: (47, 44)(1803) 0 --> (1803) 0:PUGB6, pass, NI0
			10'd41 : rdata = 48'b110001110000110100000000000100000000000000000000;
			// PEs: 8 -> 0
			// srcs: (48, 41)(1745) 2 --> (1745) 2:PUGB1, pass, NI1
			10'd42 : rdata = 48'b110001110000001100000000000100001000000000000000;
			// PEs: 56 -> 5
			// srcs: (49, 45)(1804) -4 --> (1804) -4:PUNB, pass, PEGB5
			10'd43 : rdata = 48'b110001101111111100000000000000000000000011010000;
			// PEs: 56 -> 0
			// srcs: (50, 47)(1806) 4 --> (1806) 4:PUNB, pass, NI2
			10'd44 : rdata = 48'b110001101111111100000000000100010000000000000000;
			// PEs: 56 -> 6
			// srcs: (51, 48)(1807) 4 --> (1807) 4:PUNB, pass, PEGB6
			10'd45 : rdata = 48'b110001101111111100000000000000000000000011100000;
			// PEs: 8 -> 1
			// srcs: (52, 42)(1746) -2 --> (1746) -2:PUGB1, pass, PENB
			10'd46 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 56 -> 0
			// srcs: (53, 50)(1809) 3 --> (1809) 3:PUNB, pass, NI3
			10'd47 : rdata = 48'b110001101111111100000000000100011000000000000000;
			// PEs: 56 -> 7
			// srcs: (54, 51)(1810) 3 --> (1810) 3:PUNB, pass, PEGB7
			10'd48 : rdata = 48'b110001101111111100000000000000000000000011110000;
			// PEs: 1 -> 8
			// srcs: (55, 53)(1815) -3 --> (1815) -3:PEGB1, pass, PUNB
			10'd49 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 2 -> 8
			// srcs: (56, 54)(1816) 0 --> (1816) 0:PEGB2, pass, PUNB
			10'd50 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 7 -> 16
			// srcs: (57, 55)(1822) 0 --> (1822) 0:PENB, pass, PUGB2
			10'd51 : rdata = 48'b110001101111111000000000000000000000000000001010;
			// PEs: 0 -> 1
			// srcs: (58, 43)(1745) 2 --> (1745) 2:NI1, pass, PENB
			10'd52 : rdata = 48'b110001010000000100000000000000000000000100000000;
			// PEs: 0 -> 5
			// srcs: (59, 46)(1803) 0 --> (1803) 0:NI0, pass, PEGB5
			10'd53 : rdata = 48'b110001010000000000000000000000000000000011010000;
			// PEs: 0 -> 6
			// srcs: (60, 49)(1806) 4 --> (1806) 4:NI2, pass, PEGB6
			10'd54 : rdata = 48'b110001010000001000000000000000000000000011100000;
			// PEs: 56 -> 0
			// srcs: (61, 56)(1889) 0 --> (1889) 0:PUNB, pass, NI0
			10'd55 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 56 -> 2
			// srcs: (62, 57)(1890) -2 --> (1890) -2:PUNB, pass, PEGB2
			10'd56 : rdata = 48'b110001101111111100000000000000000000000010100000;
			// PEs: 0 -> 7
			// srcs: (63, 52)(1809) 3 --> (1809) 3:NI3, pass, PEGB7
			10'd57 : rdata = 48'b110001010000001100000000000000000000000011110000;
			// PEs: 56 -> 0
			// srcs: (64, 59)(1892) 2 --> (1892) 2:PUNB, pass, NI1
			10'd58 : rdata = 48'b110001101111111100000000000100001000000000000000;
			// PEs: 56 -> 3
			// srcs: (65, 60)(1893) 0 --> (1893) 0:PUNB, pass, PEGB3
			10'd59 : rdata = 48'b110001101111111100000000000000000000000010110000;
			// PEs: 1 -> 8
			// srcs: (66, 62)(1895) -4 --> (1895) -4:PEGB1, pass, PUNB
			10'd60 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 2 -> 8
			// srcs: (67, 63)(1896) -3 --> (1896) -3:PEGB2, pass, PUNB
			10'd61 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 3 -> 8
			// srcs: (68, 64)(1898) 4 --> (1898) 4:PEGB3, pass, PUNB
			10'd62 : rdata = 48'b110001110000011000000000000000000000001000000000;
			// PEs: 4 -> 8
			// srcs: (69, 65)(1899) 0 --> (1899) 0:PEGB4, pass, PUNB
			10'd63 : rdata = 48'b110001110000100000000000000000000000001000000000;
			// PEs: 5 -> 8
			// srcs: (70, 66)(1901) -2 --> (1901) -2:PEGB5, pass, PUNB
			10'd64 : rdata = 48'b110001110000101000000000000000000000001000000000;
			// PEs: 0 -> 2
			// srcs: (71, 58)(1889) 0 --> (1889) 0:NI0, pass, PEGB2
			10'd65 : rdata = 48'b110001010000000000000000000000000000000010100000;
			// PEs: 6 -> 8
			// srcs: (72, 67)(1902) -6 --> (1902) -6:PEGB6, pass, PUNB
			10'd66 : rdata = 48'b110001110000110000000000000000000000001000000000;
			// PEs: 7 -> 8
			// srcs: (73, 68)(1904) -2 --> (1904) -2:PENB, pass, PUNB
			10'd67 : rdata = 48'b110001101111111000000000000000000000001000000000;
			// PEs: 0 -> 3
			// srcs: (74, 61)(1892) 2 --> (1892) 2:NI1, pass, PEGB3
			10'd68 : rdata = 48'b110001010000000100000000000000000000000010110000;
			// PEs: 56 -> 0
			// srcs: (75, 69)(1969) -6 --> (1969) -6:PUNB, pass, NI0
			10'd69 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 56 -> 1
			// srcs: (76, 70)(1970) 2 --> (1970) 2:PUNB, pass, PENB
			10'd70 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 1 -> 8
			// srcs: (77, 75)(1975) -2 --> (1975) -2:PEGB1, pass, PUNB
			10'd71 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 2 -> 8
			// srcs: (78, 76)(1976) -3 --> (1976) -3:PEGB2, pass, PUNB
			10'd72 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 3 -> 8
			// srcs: (79, 77)(1978) 0 --> (1978) 0:PEGB3, pass, PUNB
			10'd73 : rdata = 48'b110001110000011000000000000000000000001000000000;
			// PEs: 4 -> 8
			// srcs: (80, 78)(1979) 0 --> (1979) 0:PEGB4, pass, PUNB
			10'd74 : rdata = 48'b110001110000100000000000000000000000001000000000;
			// PEs: 5 -> 8
			// srcs: (81, 79)(1981) -6 --> (1981) -6:PEGB5, pass, PUNB
			10'd75 : rdata = 48'b110001110000101000000000000000000000001000000000;
			// PEs: 0 -> 1
			// srcs: (82, 71)(1969) -6 --> (1969) -6:NI0, pass, PENB
			10'd76 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 56 -> 0
			// srcs: (83, 72)(1972) -2 --> (1972) -2:PUNB, pass, NI0
			10'd77 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 56 -> 1
			// srcs: (84, 73)(1973) -6 --> (1973) -6:PUNB, pass, PENB
			10'd78 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 6 -> 8
			// srcs: (85, 80)(1982) 0 --> (1982) 0:PEGB6, pass, PUNB
			10'd79 : rdata = 48'b110001110000110000000000000000000000001000000000;
			// PEs: 7 -> 8
			// srcs: (86, 81)(1984) -3 --> (1984) -3:PENB, pass, PUNB
			10'd80 : rdata = 48'b110001101111111000000000000000000000001000000000;
			// PEs: 1 -> 8
			// srcs: (87, 91)(2057) 0 --> (2057) 0:PEGB1, pass, PUNB
			10'd81 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 2 -> 8
			// srcs: (88, 92)(2058) 0 --> (2058) 0:PEGB2, pass, PUNB
			10'd82 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 3 -> 8
			// srcs: (89, 93)(2060) -6 --> (2060) -6:PEGB3, pass, PUNB
			10'd83 : rdata = 48'b110001110000011000000000000000000000001000000000;
			// PEs: 0 -> 1
			// srcs: (90, 74)(1972) -2 --> (1972) -2:NI0, pass, PENB
			10'd84 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 56 -> 0
			// srcs: (91, 82)(2048) 1 --> (2048) 1:PUNB, pass, NI0
			10'd85 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 56 -> 1
			// srcs: (92, 83)(2049) 0 --> (2049) 0:PUNB, pass, PENB
			10'd86 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 4 -> 8
			// srcs: (93, 94)(2061) -2 --> (2061) -2:PEGB4, pass, PUNB
			10'd87 : rdata = 48'b110001110000100000000000000000000000001000000000;
			// PEs: 1 -> 8
			// srcs: (94, 104)(2137) 0 --> (2137) 0:PEGB1, pass, PUNB
			10'd88 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 2 -> 8
			// srcs: (95, 105)(2138) 0 --> (2138) 0:PEGB2, pass, PUNB
			10'd89 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 3 -> 8
			// srcs: (96, 106)(2140) 2 --> (2140) 2:PEGB3, pass, PUNB
			10'd90 : rdata = 48'b110001110000011000000000000000000000001000000000;
			// PEs: 4 -> 8
			// srcs: (97, 107)(2141) -2 --> (2141) -2:PEGB4, pass, PUNB
			10'd91 : rdata = 48'b110001110000100000000000000000000000001000000000;
			// PEs: 0 -> 1
			// srcs: (98, 84)(2048) 1 --> (2048) 1:NI0, pass, PENB
			10'd92 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 56 -> 0
			// srcs: (99, 85)(2051) -4 --> (2051) -4:PUNB, pass, NI0
			10'd93 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 56 -> 1
			// srcs: (100, 86)(2052) 0 --> (2052) 0:PUNB, pass, PENB
			10'd94 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 5 -> 8
			// srcs: (101, 108)(2143) 0 --> (2143) 0:PEGB5, pass, PUNB
			10'd95 : rdata = 48'b110001110000101000000000000000000000001000000000;
			// PEs: 6 -> 8
			// srcs: (102, 109)(2144) 0 --> (2144) 0:PEGB6, pass, PUNB
			10'd96 : rdata = 48'b110001110000110000000000000000000000001000000000;
			// PEs: 7 -> 8
			// srcs: (103, 110)(2146) -4 --> (2146) -4:PENB, pass, PUNB
			10'd97 : rdata = 48'b110001101111111000000000000000000000001000000000;
			// PEs: 7 -> 8
			// srcs: (104, 114)(2226) 0 --> (2226) 0:PENB, pass, PUNB
			10'd98 : rdata = 48'b110001101111111000000000000000000000001000000000;
			// PEs: 3 -> 16
			// srcs: (105, 143)(2365) -8 --> (2365) -8:PEGB3, pass, PUGB2
			10'd99 : rdata = 48'b110001110000011000000000000000000000000000001010;
			// PEs: 0 -> 1
			// srcs: (106, 87)(2051) -4 --> (2051) -4:NI0, pass, PENB
			10'd100 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 56 -> 0
			// srcs: (107, 88)(2054) -6 --> (2054) -6:PUNB, pass, NI0
			10'd101 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 56 -> 1
			// srcs: (108, 89)(2055) 0 --> (2055) 0:PUNB, pass, PENB
			10'd102 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 4 -> 32
			// srcs: (109, 144)(2369) -1 --> (2369) -1:PEGB4, pass, PUGB4
			10'd103 : rdata = 48'b110001110000100000000000000000000000000000001100;
			// PEs: 1 -> 40
			// srcs: (110, 151)(1631) 0 --> (1631) 0:PEGB1, pass, PUGB5
			10'd104 : rdata = 48'b110001110000001000000000000000000000000000001101;
			// PEs: 6 -> 16
			// srcs: (111, 156)(1646) 0 --> (1646) 0:PEGB6, pass, PUGB2
			10'd105 : rdata = 48'b110001110000110000000000000000000000000000001010;
			// PEs: 1 -> 48
			// srcs: (112, 115)(1573) 6 --> (1573) 6:PEGB1, pass, PUGB6
			10'd106 : rdata = 48'b110001110000001000000000000000000000000000001110;
			// PEs: 3 -> 56
			// srcs: (113, 117)(1575) 0 --> (1575) 0:PEGB3, pass, PUGB7
			10'd107 : rdata = 48'b110001110000011000000000000000000000000000001111;
			// PEs: 0 -> 1
			// srcs: (114, 90)(2054) -6 --> (2054) -6:NI0, pass, PENB
			10'd108 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 56 -> 0
			// srcs: (115, 95)(2128) -4 --> (2128) -4:PUNB, pass, NI0
			10'd109 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 56 -> 1
			// srcs: (116, 96)(2129) 6 --> (2129) 6:PUNB, pass, PENB
			10'd110 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 3 -> 8
			// srcs: (117, 122)(1818) 2 --> (1818) 2:PEGB3, pass, PUNB
			10'd111 : rdata = 48'b110001110000011000000000000000000000001000000000;
			// PEs: 3 -> 24
			// srcs: (118, 153)(1637) 0 --> (1637) 0:PEGB3, pass, PUGB3
			10'd112 : rdata = 48'b110001110000011000000000000000000000000000001011;
			// PEs: 4 -> 32
			// srcs: (119, 154)(1640) -1 --> (1640) -1:PEGB4, pass, PUGB4
			10'd113 : rdata = 48'b110001110000100000000000000000000000000000001100;
			// PEs: 2 -> 48
			// srcs: (120, 116)(1574) 3 --> (1574) 3:PEGB2, pass, PUGB6
			10'd114 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 5 -> 48
			// srcs: (121, 145)(2371) 9 --> (2371) 9:PEGB5, pass, PUGB6
			10'd115 : rdata = 48'b110001110000101000000000000000000000000000001110;
			// PEs: 0 -> 1
			// srcs: (122, 97)(2128) -4 --> (2128) -4:NI0, pass, PENB
			10'd116 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 56 -> 0
			// srcs: (123, 98)(2131) 2 --> (2131) 2:PUNB, pass, NI0
			10'd117 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 56 -> 1
			// srcs: (124, 99)(2132) -2 --> (2132) -2:PUNB, pass, PENB
			10'd118 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 4 -> 56
			// srcs: (125, 118)(1576) 0 --> (1576) 0:PEGB4, pass, PUGB7
			10'd119 : rdata = 48'b110001110000100000000000000000000000000000001111;
			// PEs: 4 -> 8
			// srcs: (126, 123)(1819) 9 --> (1819) 9:PEGB4, pass, PUNB
			10'd120 : rdata = 48'b110001110000100000000000000000000000001000000000;
			// PEs: 6 -> 56
			// srcs: (127, 146)(2374) 6 --> (2374) 6:PEGB6, pass, PUGB7
			10'd121 : rdata = 48'b110001110000110000000000000000000000000000001111;
			// PEs: 7 -> 48
			// srcs: (128, 147)(2376) -6 --> (2376) -6:PENB, pass, PUGB6
			10'd122 : rdata = 48'b110001101111111000000000000000000000000000001110;
			// PEs: 0 -> 1
			// srcs: (130, 100)(2131) 2 --> (2131) 2:NI0, pass, PENB
			10'd123 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 56 -> 0
			// srcs: (131, 101)(2134) 2 --> (2134) 2:PUNB, pass, NI0
			10'd124 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 56 -> 1
			// srcs: (132, 102)(2135) -3 --> (2135) -3:PUNB, pass, PENB
			10'd125 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 7 -> 24
			// srcs: (133, 157)(1649) 0 --> (1649) 0:PENB, pass, PUGB3
			10'd126 : rdata = 48'b110001101111111000000000000000000000000000001011;
			// PEs: 5 -> 8
			// srcs: (134, 124)(1820) 2 --> (1820) 2:PEGB5, pass, PUNB
			10'd127 : rdata = 48'b110001110000101000000000000000000000001000000000;
			// PEs: 3 -> 48
			// srcs: (136, 170)(2508) 6 --> (2508) 6:PEGB3, pass, PUGB6
			10'd128 : rdata = 48'b110001110000011000000000000000000000000000001110;
			// PEs: 4 -> 16
			// srcs: (137, 171)(2510) -2 --> (2510) -2:PEGB4, pass, PUGB2
			10'd129 : rdata = 48'b110001110000100000000000000000000000000000001010;
			// PEs: 0 -> 1
			// srcs: (138, 103)(2134) 2 --> (2134) 2:NI0, pass, PENB
			10'd130 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 56 -> 0
			// srcs: (139, 111)(2214) -3 --> (2214) -3:PUNB, pass, NI0
			10'd131 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 56 -> 1
			// srcs: (140, 112)(2215) 2 --> (2215) 2:PUNB, pass, PENB
			10'd132 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 1 -> 56
			// srcs: (141, 172)(2521) 4 --> (2521) 4:PEGB1, pass, PUGB7
			10'd133 : rdata = 48'b110001110000001000000000000000000000000000001111;
			// PEs: 6 -> 8
			// srcs: (142, 125)(1821) 0 --> (1821) 0:PEGB6, pass, PUNB
			10'd134 : rdata = 48'b110001110000110000000000000000000000001000000000;
			// PEs: 2 -> 24
			// srcs: (143, 169)(2505) 8 --> (2505) 8:PEGB2, pass, PUGB3
			10'd135 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 6 -> 32
			// srcs: (144, 180)(1830) 0 --> (1830) 0:PEGB6, pass, PUGB4
			10'd136 : rdata = 48'b110001110000110000000000000000000000000000001100;
			// PEs: 6 -> 40
			// srcs: (145, 204)(2010) -2 --> (2010) -2:PEGB6, pass, PUGB5
			10'd137 : rdata = 48'b110001110000110000000000000000000000000000001101;
			// PEs: 0 -> 1
			// srcs: (146, 113)(2214) -3 --> (2214) -3:NI0, pass, PENB
			10'd138 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 5 -> 8
			// srcs: (150, 129)(2063) 0 --> (2063) 0:PEGB5, pass, PUNB
			10'd139 : rdata = 48'b110001110000101000000000000000000000001000000000;
			// PEs: 1 -> 24
			// srcs: (151, 173)(2526) 0 --> (2526) 0:PEGB1, pass, PUGB3
			10'd140 : rdata = 48'b110001110000001000000000000000000000000000001011;
			// PEs: 4 -> 56
			// srcs: (152, 178)(1824) 3 --> (1824) 3:PEGB4, pass, PUGB7
			10'd141 : rdata = 48'b110001110000100000000000000000000000000000001111;
			// PEs: 5 -> 16
			// srcs: (153, 179)(1827) 3 --> (1827) 3:PEGB5, pass, PUGB2
			10'd142 : rdata = 48'b110001110000101000000000000000000000000000001010;
			// PEs: 2 -> 48
			// srcs: (154, 188)(2668) -2 --> (2668) -2:PEGB2, pass, PUGB6
			10'd143 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 1 -> 32
			// srcs: (155, 199)(1995) 4 --> (1995) 4:PEGB1, pass, PUGB4
			10'd144 : rdata = 48'b110001110000001000000000000000000000000000001100;
			// PEs: 7 -> 40
			// srcs: (156, 205)(2013) 2 --> (2013) 2:PENB, pass, PUGB5
			10'd145 : rdata = 48'b110001101111111000000000000000000000000000001101;
			// PEs: 6 -> 8
			// srcs: (158, 130)(2064) -3 --> (2064) -3:PEGB6, pass, PUNB
			10'd146 : rdata = 48'b110001110000110000000000000000000000001000000000;
			// PEs: 7 -> 24
			// srcs: (159, 181)(1833) 0 --> (1833) 0:PENB, pass, PUGB3
			10'd147 : rdata = 48'b110001101111111000000000000000000000000000001011;
			// PEs: 3 -> 56
			// srcs: (162, 189)(2673) 2 --> (2673) 2:PEGB3, pass, PUGB7
			10'd148 : rdata = 48'b110001110000011000000000000000000000000000001111;
			// PEs: 7 -> 8
			// srcs: (163, 131)(2065) 0 --> (2065) 0:PENB, pass, PUNB
			10'd149 : rdata = 48'b110001101111111000000000000000000000001000000000;
			// PEs: 5 -> 48
			// srcs: (164, 203)(2007) 0 --> (2007) 0:PEGB5, pass, PUGB6
			10'd150 : rdata = 48'b110001110000101000000000000000000000000000001110;
			// PEs: 2 -> 32
			// srcs: (165, 222)(2182) -3 --> (2182) -3:PEGB2, pass, PUGB4
			10'd151 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 6 -> 16
			// srcs: (166, 226)(2194) -1 --> (2194) -1:PEGB6, pass, PUGB2
			10'd152 : rdata = 48'b110001110000110000000000000000000000000000001010;
			// PEs: 1 -> 24
			// srcs: (167, 216)(2831) -4 --> (2831) -4:PEGB1, pass, PUGB3
			10'd153 : rdata = 48'b110001110000001000000000000000000000000000001011;
			// PEs: 7 -> 8
			// srcs: (168, 138)(2308) 6 --> (2308) 6:PENB, pass, PUNB
			10'd154 : rdata = 48'b110001101111111000000000000000000000001000000000;
			// PEs: 3 -> 56
			// srcs: (171, 201)(2001) 0 --> (2001) 0:PEGB3, pass, PUGB7
			10'd155 : rdata = 48'b110001110000011000000000000000000000000000001111;
			// PEs: 1 -> 48
			// srcs: (172, 219)(2910) 0 --> (2910) 0:PEGB1, pass, PUGB6
			10'd156 : rdata = 48'b110001110000001000000000000000000000000000001110;
			// PEs: 7 -> 16
			// srcs: (173, 234)(3003) 0 --> (3003) 0:PENB, pass, PUGB2
			10'd157 : rdata = 48'b110001101111111000000000000000000000000000001010;
			// PEs: 2 -> 8
			// srcs: (176, 152)(1634) 3 --> (1634) 3:PEGB2, pass, PUNB
			10'd158 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 5 -> 24
			// srcs: (177, 236)(3080) 0 --> (3080) 0:PEGB5, pass, PUGB3
			10'd159 : rdata = 48'b110001110000101000000000000000000000000000001011;
			// PEs: 1 -> 56
			// srcs: (179, 217)(2833) -6 --> (2833) -6:PEGB1, pass, PUGB7
			10'd160 : rdata = 48'b110001110000001000000000000000000000000000001111;
			// PEs: 1 -> 48
			// srcs: (180, 220)(2912) -1 --> (2912) -1:PEGB1, pass, PUGB6
			10'd161 : rdata = 48'b110001110000001000000000000000000000000000001110;
			// PEs: 1 -> 8
			// srcs: (184, 158)(2442) -6 --> (2442) -6:PEGB1, pass, PUNB
			10'd162 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 1 -> 48
			// srcs: (188, 221)(2179) -3 --> (2179) -3:PEGB1, pass, PUGB6
			10'd163 : rdata = 48'b110001110000001000000000000000000000000000001110;
			// PEs: 3 -> 56
			// srcs: (189, 223)(2185) -2 --> (2185) -2:PEGB3, pass, PUGB7
			10'd164 : rdata = 48'b110001110000011000000000000000000000000000001111;
			// PEs: 2 -> 8
			// srcs: (192, 176)(1814) -6 --> (1814) -6:PEGB2, pass, PUNB
			10'd165 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 4 -> 56
			// srcs: (197, 224)(2188) 0 --> (2188) 0:PEGB4, pass, PUGB7
			10'd166 : rdata = 48'b110001110000100000000000000000000000000000001111;
			// PEs: 5 -> 48
			// srcs: (198, 225)(2191) 6 --> (2191) 6:PEGB5, pass, PUGB6
			10'd167 : rdata = 48'b110001110000101000000000000000000000000000001110;
			// PEs: 3 -> 8
			// srcs: (200, 177)(1817) -1 --> (1817) -1:PEGB3, pass, PUNB
			10'd168 : rdata = 48'b110001110000011000000000000000000000001000000000;
			// PEs: 7 -> 48
			// srcs: (203, 227)(2197) 0 --> (2197) 0:PENB, pass, PUGB6
			10'd169 : rdata = 48'b110001101111111000000000000000000000000000001110;
			// PEs: 1 -> 8
			// srcs: (208, 194)(2751) -4 --> (2751) -4:PEGB1, pass, PUNB
			10'd170 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 7 -> 48
			// srcs: (209, 237)(3082) -4 --> (3082) -4:PENB, pass, PUGB6
			10'd171 : rdata = 48'b110001101111111000000000000000000000000000001110;
			// PEs: 48 -> 0
			// srcs: (213, 119)(1722) -6 --> (1722) -6:PUGB6, pass, NI0
			10'd172 : rdata = 48'b110001110000110100000000000100000000000000000000;
			// PEs: 56 -> 2
			// srcs: (214, 120)(1723) 0 --> (1723) 0:PUNB, pass, PEGB2
			10'd173 : rdata = 48'b110001101111111100000000000000000000000010100000;
			// PEs: 56 -> 0
			// srcs: (215, 126)(1967) 0 --> (1967) 0:PUNB, pass, NI1
			10'd174 : rdata = 48'b110001101111111100000000000100001000000000000000;
			// PEs: 56 -> 1
			// srcs: (216, 127)(1968) 0 --> (1968) 0:PUNB, pass, PENB
			10'd175 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 2 -> 8
			// srcs: (217, 200)(1998) 0 --> (1998) 0:PEGB2, pass, PUNB
			10'd176 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 0 -> 1
			// srcs: (222, 128)(1967) 0 --> (1967) 0:NI1, pass, PENB
			10'd177 : rdata = 48'b110001010000000100000000000000000000000100000000;
			// PEs: 0 -> 2
			// srcs: (223, 121)(1722) -6 --> (1722) -6:NI0, pass, PEGB2
			10'd178 : rdata = 48'b110001010000000000000000000000000000000010100000;
			// PEs: 56 -> 0
			// srcs: (225, 132)(2210) -1 --> (2210) -1:PUNB, pass, NI0
			10'd179 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 4 -> 8
			// srcs: (226, 202)(2004) -2 --> (2004) -2:PEGB4, pass, PUNB
			10'd180 : rdata = 48'b110001110000100000000000000000000000001000000000;
			// PEs: 1 -> 8
			// srcs: (234, 215)(2827) 1 --> (2827) 1:PEGB1, pass, PUNB
			10'd181 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 56 -> 1
			// srcs: (241, 133)(2211) -1 --> (2211) -1:PUNB, pass, PENB
			10'd182 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 1 -> 8
			// srcs: (242, 218)(2907) 2 --> (2907) 2:PEGB1, pass, PUNB
			10'd183 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 0 -> 1
			// srcs: (247, 134)(2210) -1 --> (2210) -1:NI0, pass, PENB
			10'd184 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 56 -> 0
			// srcs: (248, 135)(2212) 0 --> (2212) 0:PUNB, pass, NI0
			10'd185 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 56 -> 1
			// srcs: (249, 136)(2213) 0 --> (2213) 0:PUNB, pass, PENB
			10'd186 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 1 -> 8
			// srcs: (250, 231)(2994) -1 --> (2994) -1:PEGB1, pass, PUNB
			10'd187 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 0 -> 1
			// srcs: (255, 137)(2212) 0 --> (2212) 0:NI0, pass, PENB
			10'd188 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 16 -> 0
			// srcs: (256, 139)(2360) -10 --> (2360) -10:PUGB2, pass, NI0
			10'd189 : rdata = 48'b110001110000010100000000000100000000000000000000;
			// PEs: 40 -> 1
			// srcs: (257, 140)(1579) -6 --> (1579) -6:PUGB5, pass, PENB
			10'd190 : rdata = 48'b110001110000101100000000000000000000000100000000;
			// PEs: 4 -> 8
			// srcs: (258, 232)(2997) 1 --> (2997) 1:PEGB4, pass, PUNB
			10'd191 : rdata = 48'b110001110000100000000000000000000000001000000000;
			// PEs: 0 -> 1
			// srcs: (263, 141)(2360) -10 --> (2360) -10:NI0, pass, PENB
			10'd192 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 40 -> 1
			// srcs: (264, 142)(1582) -6 --> (1582) -6:PUGB5, pass, PENB
			10'd193 : rdata = 48'b110001110000101100000000000000000000000100000000;
			// PEs: 8 -> 0
			// srcs: (265, 148)(2392) -8 --> (2392) -8:PUGB1, pass, NI0
			10'd194 : rdata = 48'b110001110000001100000000000100000000000000000000;
			// PEs: 56 -> 1
			// srcs: (266, 149)(1612) 0 --> (1612) 0:PUNB, pass, PENB
			10'd195 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 5 -> 8
			// srcs: (267, 233)(2999) 0 --> (2999) 0:PEGB5, pass, PUNB
			10'd196 : rdata = 48'b110001110000101000000000000000000000001000000000;
			// PEs: 1 -> 16
			// srcs: (270, 244)(2361) -16 --> (2361) -16:PEGB1, pass, PUGB2
			10'd197 : rdata = 48'b110001110000001000000000000000000000000000001010;
			// PEs: 1 -> 48
			// srcs: (271, 245)(2364) -11 --> (2364) -11:PEGB1, pass, PUGB6
			10'd198 : rdata = 48'b110001110000001000000000000000000000000000001110;
			// PEs: 0 -> 1
			// srcs: (272, 150)(2392) -8 --> (2392) -8:NI0, pass, PENB
			10'd199 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 24 -> 1
			// srcs: (273, 155)(2422) -5 --> (2422) -5:PUGB3, pass, PENB
			10'd200 : rdata = 48'b110001110000011100000000000000000000000100000000;
			// PEs: 32 -> 0
			// srcs: (274, 159)(2462) 1 --> (2462) 1:PUGB4, pass, NI0
			10'd201 : rdata = 48'b110001110000100100000000000100000000000000000000;
			// PEs: 16 -> 1
			// srcs: (275, 160)(1683) 1 --> (1683) 1:PUGB2, pass, PENB
			10'd202 : rdata = 48'b110001110000010100000000000000000000000100000000;
			// PEs: 1 -> 8
			// srcs: (280, 250)(2423) -3 --> (2423) -3:PEGB1, pass, PUNB
			10'd203 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 0 -> 1
			// srcs: (281, 161)(2462) 1 --> (2462) 1:NI0, pass, PENB
			10'd204 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 48 -> 0
			// srcs: (282, 162)(2483) -1 --> (2483) -1:PUGB6, pass, NI0
			10'd205 : rdata = 48'b110001110000110100000000000100000000000000000000;
			// PEs: 24 -> 1
			// srcs: (283, 163)(1704) -2 --> (1704) -2:PUGB3, pass, PENB
			10'd206 : rdata = 48'b110001110000011100000000000000000000000100000000;
			// PEs: 1 -> 56
			// srcs: (288, 251)(2463) 2 --> (2463) 2:PEGB1, pass, PUGB7
			10'd207 : rdata = 48'b110001110000001000000000000000000000000000001111;
			// PEs: 0 -> 1
			// srcs: (289, 164)(2483) -1 --> (2483) -1:NI0, pass, PENB
			10'd208 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 56 -> 0
			// srcs: (290, 165)(2494) 7 --> (2494) 7:PUNB, pass, NI0
			10'd209 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 24 -> 1
			// srcs: (291, 166)(1716) -2 --> (1716) -2:PUGB3, pass, PENB
			10'd210 : rdata = 48'b110001110000011100000000000000000000000100000000;
			// PEs: 1 -> 8
			// srcs: (296, 255)(2484) -3 --> (2484) -3:PEGB1, pass, PUNB
			10'd211 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 0 -> 1
			// srcs: (297, 167)(2494) 7 --> (2494) 7:NI0, pass, PENB
			10'd212 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 56 -> 1
			// srcs: (298, 168)(2502) 7 --> (2502) 7:PUNB, pass, PENB
			10'd213 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 56 -> 1
			// srcs: (299, 174)(1805) 0 --> (1805) 0:PUNB, pass, PENB
			10'd214 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 1 -> 8
			// srcs: (304, 256)(2495) 5 --> (2495) 5:PEGB1, pass, PUNB
			10'd215 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 1 -> 32
			// srcs: (305, 257)(2504) 1 --> (2504) 1:PEGB1, pass, PUGB4
			10'd216 : rdata = 48'b110001110000001000000000000000000000000000001100;
			// PEs: 56 -> 1
			// srcs: (525, 175)(1808) 0 --> (1808) 0:PUNB, pass, PENB
			10'd217 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 32 -> 0
			// srcs: (526, 182)(2629) 3 --> (2629) 3:PUGB4, pass, NI0
			10'd218 : rdata = 48'b110001110000100100000000000100000000000000000000;
			// PEs: 8 -> 1
			// srcs: (527, 183)(1851) 0 --> (1851) 0:PUGB1, pass, PENB
			10'd219 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 0 -> 1
			// srcs: (533, 184)(2629) 3 --> (2629) 3:NI0, pass, PENB
			10'd220 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 48 -> 0
			// srcs: (534, 185)(2663) -2 --> (2663) -2:PUGB6, pass, NI0
			10'd221 : rdata = 48'b110001110000110100000000000100000000000000000000;
			// PEs: 24 -> 1
			// srcs: (535, 186)(1885) -2 --> (1885) -2:PUGB3, pass, PENB
			10'd222 : rdata = 48'b110001110000011100000000000000000000000100000000;
			// PEs: 1 -> 8
			// srcs: (540, 265)(2630) 3 --> (2630) 3:PEGB1, pass, PUNB
			10'd223 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 0 -> 1
			// srcs: (541, 187)(2663) -2 --> (2663) -2:NI0, pass, PENB
			10'd224 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 8 -> 0
			// srcs: (542, 190)(2680) -8 --> (2680) -8:PUGB1, pass, NI0
			10'd225 : rdata = 48'b110001110000001100000000000100000000000000000000;
			// PEs: 32 -> 1
			// srcs: (543, 191)(1903) 3 --> (1903) 3:PUGB4, pass, PENB
			10'd226 : rdata = 48'b110001110000100100000000000000000000000100000000;
			// PEs: 1 -> 24
			// srcs: (548, 266)(2664) -4 --> (2664) -4:PEGB1, pass, PUGB3
			10'd227 : rdata = 48'b110001110000001000000000000000000000000000001011;
			// PEs: 0 -> 1
			// srcs: (549, 192)(2680) -8 --> (2680) -8:NI0, pass, PENB
			10'd228 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 56 -> 1
			// srcs: (550, 193)(2748) -1 --> (2748) -1:PUNB, pass, PENB
			10'd229 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 56 -> 6
			// srcs: (551, 195)(1974) 6 --> (1974) 6:PUNB, pass, PEGB6
			10'd230 : rdata = 48'b110001101111111100000000000000000000000011100000;
			// PEs: 8 -> 0
			// srcs: (552, 196)(2765) -4 --> (2765) -4:PUGB1, pass, NI0
			10'd231 : rdata = 48'b110001110000001100000000000100000000000000000000;
			// PEs: 56 -> 1
			// srcs: (553, 197)(1986) 0 --> (1986) 0:PUNB, pass, PENB
			10'd232 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 1 -> 48
			// srcs: (556, 267)(2681) -5 --> (2681) -5:PEGB1, pass, PUGB6
			10'd233 : rdata = 48'b110001110000001000000000000000000000000000001110;
			// PEs: 1 -> 8
			// srcs: (557, 271)(2750) -1 --> (2750) -1:PEGB1, pass, PUNB
			10'd234 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 2 -> 8
			// srcs: (558, 284)(2993) -2 --> (2993) -2:PEGB2, pass, PUNB
			10'd235 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 0 -> 1
			// srcs: (559, 198)(2765) -4 --> (2765) -4:NI0, pass, PENB
			10'd236 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 40 -> 0
			// srcs: (560, 206)(2799) -2 --> (2799) -2:PUGB5, pass, NI0
			10'd237 : rdata = 48'b110001110000101100000000000100000000000000000000;
			// PEs: 8 -> 1
			// srcs: (561, 207)(2020) 1 --> (2020) 1:PUGB1, pass, PENB
			10'd238 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 1 -> 16
			// srcs: (566, 273)(2766) -4 --> (2766) -4:PEGB1, pass, PUGB2
			10'd239 : rdata = 48'b110001110000001000000000000000000000000000001010;
			// PEs: 0 -> 1
			// srcs: (567, 208)(2799) -2 --> (2799) -2:NI0, pass, PENB
			10'd240 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 48 -> 0
			// srcs: (568, 209)(2808) -6 --> (2808) -6:PUGB6, pass, NI0
			10'd241 : rdata = 48'b110001110000110100000000000100000000000000000000;
			// PEs: 8 -> 1
			// srcs: (569, 210)(2029) 0 --> (2029) 0:PUGB1, pass, PENB
			10'd242 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 1 -> 16
			// srcs: (574, 274)(2800) -1 --> (2800) -1:PEGB1, pass, PUGB2
			10'd243 : rdata = 48'b110001110000001000000000000000000000000000001010;
			// PEs: 0 -> 1
			// srcs: (575, 211)(2808) -6 --> (2808) -6:NI0, pass, PENB
			10'd244 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 56 -> 0
			// srcs: (576, 212)(2815) -1 --> (2815) -1:PUNB, pass, NI0
			10'd245 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 8 -> 1
			// srcs: (577, 213)(2038) -2 --> (2038) -2:PUGB1, pass, PENB
			10'd246 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 1 -> 40
			// srcs: (582, 275)(2809) -6 --> (2809) -6:PEGB1, pass, PUGB5
			10'd247 : rdata = 48'b110001110000001000000000000000000000000000001101;
			// PEs: 0 -> 1
			// srcs: (583, 214)(2815) -1 --> (2815) -1:NI0, pass, PENB
			10'd248 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 56 -> 0
			// srcs: (584, 228)(2985) -2 --> (2985) -2:PUNB, pass, NI0
			10'd249 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 8 -> 1
			// srcs: (585, 229)(2209) 0 --> (2209) 0:PUGB1, pass, PENB
			10'd250 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 1 -> 48
			// srcs: (590, 276)(2816) -3 --> (2816) -3:PEGB1, pass, PUGB6
			10'd251 : rdata = 48'b110001110000001000000000000000000000000000001110;
			// PEs: 0 -> 1
			// srcs: (591, 230)(2985) -2 --> (2985) -2:NI0, pass, PENB
			10'd252 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 40 -> 1
			// srcs: (592, 235)(2301) 0 --> (2301) 0:PUGB5, pass, PENB
			10'd253 : rdata = 48'b110001110000101100000000000000000000000100000000;
			// PEs: 16 -> 0
			// srcs: (593, 238)(3096) 2 --> (3096) 2:PUGB2, pass, NI0
			10'd254 : rdata = 48'b110001110000010100000000000100000000000000000000;
			// PEs: 48 -> 1
			// srcs: (594, 239)(2320) 0 --> (2320) 0:PUGB6, pass, PENB
			10'd255 : rdata = 48'b110001110000110100000000000000000000000100000000;
			// PEs: 1 -> 16
			// srcs: (598, 283)(2986) -2 --> (2986) -2:PEGB1, pass, PUGB2
			10'd256 : rdata = 48'b110001110000001000000000000000000000000000001010;
			// PEs: 0 -> 1
			// srcs: (605, 240)(3096) 2 --> (3096) 2:NI0, pass, PENB
			10'd257 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 32 -> 0
			// srcs: (606, 241)(3119) -4 --> (3119) -4:PUGB4, pass, NI0
			10'd258 : rdata = 48'b110001110000100100000000000100000000000000000000;
			// PEs: 56 -> 1
			// srcs: (607, 242)(2344) 0 --> (2344) 0:PUNB, pass, PENB
			10'd259 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 1 -> 24
			// srcs: (608, 288)(3078) -2 --> (3078) -2:PEGB1, pass, PUGB3
			10'd260 : rdata = 48'b110001110000001000000000000000000000000000001011;
			// PEs: 0 -> 1
			// srcs: (613, 243)(3119) -4 --> (3119) -4:NI0, pass, PENB
			10'd261 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 32 -> 0
			// srcs: (614, 246)(2370) 1 --> (2370) 1:PUGB4, pass, NI0
			10'd262 : rdata = 48'b110001110000100100000000000100000000000000000000;
			// PEs: 48 -> 1
			// srcs: (615, 247)(2372) 11 --> (2372) 11:PUGB6, pass, PENB
			10'd263 : rdata = 48'b110001110000110100000000000000000000000100000000;
			// PEs: 1 -> 8
			// srcs: (620, 293)(3120) -4 --> (3120) -4:PEGB1, pass, PUNB
			10'd264 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 0 -> 1
			// srcs: (621, 248)(2370) 1 --> (2370) 1:NI0, pass, PENB
			10'd265 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 56 -> 1
			// srcs: (622, 249)(2395) 6 --> (2395) 6:PUNB, pass, PENB
			10'd266 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 8 -> 0
			// srcs: (623, 252)(2472) 15 --> (2472) 15:PUGB1, pass, NI0
			10'd267 : rdata = 48'b110001110000001100000000000100000000000000000000;
			// PEs: 48 -> 1
			// srcs: (624, 253)(2474) -3 --> (2474) -3:PUGB6, pass, PENB
			10'd268 : rdata = 48'b110001110000110100000000000000000000000100000000;
			// PEs: 3 -> 8
			// srcs: (625, 302)(2591) 14 --> (2591) 14:PEGB3, pass, PUNB
			10'd269 : rdata = 48'b110001110000011000000000000000000000001000000000;
			// PEs: 1 -> 16
			// srcs: (629, 295)(2396) -2 --> (2396) -2:PEGB1, pass, PUGB2
			10'd270 : rdata = 48'b110001110000001000000000000000000000000000001010;
			// PEs: 0 -> 1
			// srcs: (630, 254)(2472) 15 --> (2472) 15:NI0, pass, PENB
			10'd271 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 8 -> 0
			// srcs: (631, 258)(2520) -1 --> (2520) -1:PUGB1, pass, NI0
			10'd272 : rdata = 48'b110001110000001100000000000100000000000000000000;
			// PEs: 56 -> 1
			// srcs: (632, 259)(2522) 5 --> (2522) 5:PUNB, pass, PENB
			10'd273 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 1 -> 48
			// srcs: (637, 296)(2475) 12 --> (2475) 12:PEGB1, pass, PUGB6
			10'd274 : rdata = 48'b110001110000001000000000000000000000000000001110;
			// PEs: 0 -> 1
			// srcs: (638, 260)(2520) -1 --> (2520) -1:NI0, pass, PENB
			10'd275 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 1 -> 40
			// srcs: (645, 300)(2523) 4 --> (2523) 4:PEGB1, pass, PUGB5
			10'd276 : rdata = 48'b110001110000001000000000000000000000000000001101;
			// PEs: 56 -> 1
			// srcs: (950, 261)(2582) 1 --> (2582) 1:PUNB, pass, PENB
			10'd277 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 24 -> 0
			// srcs: (951, 262)(2625) 10 --> (2625) 10:PUGB3, pass, NI0
			10'd278 : rdata = 48'b110001110000011100000000000100000000000000000000;
			// PEs: 8 -> 1
			// srcs: (952, 263)(2627) 6 --> (2627) 6:PUGB1, pass, PENB
			10'd279 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 0 -> 1
			// srcs: (958, 264)(2625) 10 --> (2625) 10:NI0, pass, PENB
			10'd280 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 8 -> 0
			// srcs: (959, 268)(2685) 4 --> (2685) 4:PUGB1, pass, NI0
			10'd281 : rdata = 48'b110001110000001100000000000100000000000000000000;
			// PEs: 32 -> 1
			// srcs: (960, 269)(2687) -7 --> (2687) -7:PUGB4, pass, PENB
			10'd282 : rdata = 48'b110001110000100100000000000000000000000100000000;
			// PEs: 1 -> 8
			// srcs: (965, 303)(2628) 16 --> (2628) 16:PEGB1, pass, PUNB
			10'd283 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 0 -> 1
			// srcs: (966, 270)(2685) 4 --> (2685) 4:NI0, pass, PENB
			10'd284 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 56 -> 1
			// srcs: (967, 272)(2757) -5 --> (2757) -5:PUNB, pass, PENB
			10'd285 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 24 -> 0
			// srcs: (968, 277)(2832) 0 --> (2832) 0:PUGB3, pass, NI0
			10'd286 : rdata = 48'b110001110000011100000000000100000000000000000000;
			// PEs: 56 -> 1
			// srcs: (969, 278)(2834) -6 --> (2834) -6:PUNB, pass, PENB
			10'd287 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 1 -> 16
			// srcs: (973, 307)(2688) -3 --> (2688) -3:PEGB1, pass, PUGB2
			10'd288 : rdata = 48'b110001110000001000000000000000000000000000001010;
			// PEs: 0 -> 1
			// srcs: (980, 279)(2832) 0 --> (2832) 0:NI0, pass, PENB
			10'd289 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 40 -> 0
			// srcs: (981, 280)(2950) -8 --> (2950) -8:PUGB5, pass, NI0
			10'd290 : rdata = 48'b110001110000101100000000000100000000000000000000;
			// PEs: 56 -> 1
			// srcs: (982, 281)(2952) 4 --> (2952) 4:PUNB, pass, PENB
			10'd291 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 1 -> 8
			// srcs: (983, 308)(2758) -7 --> (2758) -7:PEGB1, pass, PUNB
			10'd292 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 1 -> 56
			// srcs: (987, 309)(2835) -6 --> (2835) -6:PEGB1, pass, PUGB7
			10'd293 : rdata = 48'b110001110000001000000000000000000000000000001111;
			// PEs: 0 -> 1
			// srcs: (988, 282)(2950) -8 --> (2950) -8:NI0, pass, PENB
			10'd294 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 32 -> 0
			// srcs: (989, 285)(3065) -3 --> (3065) -3:PUGB4, pass, NI0
			10'd295 : rdata = 48'b110001110000100100000000000100000000000000000000;
			// PEs: 56 -> 1
			// srcs: (990, 286)(3067) -2 --> (3067) -2:PUNB, pass, PENB
			10'd296 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 56 -> 4
			// srcs: (991, 289)(3095) -3 --> (3095) -3:PUNB, pass, PEGB4
			10'd297 : rdata = 48'b110001101111111100000000000000000000000011000000;
			// PEs: 1 -> 8
			// srcs: (995, 313)(2953) -4 --> (2953) -4:PEGB1, pass, PUNB
			10'd298 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 0 -> 1
			// srcs: (996, 287)(3065) -3 --> (3065) -3:NI0, pass, PENB
			10'd299 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 24 -> 0
			// srcs: (997, 290)(3113) -6 --> (3113) -6:PUGB3, pass, NI0
			10'd300 : rdata = 48'b110001110000011100000000000100000000000000000000;
			// PEs: 8 -> 1
			// srcs: (998, 291)(3115) 4 --> (3115) 4:PUGB1, pass, PENB
			10'd301 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 1 -> 32
			// srcs: (1003, 317)(3068) -5 --> (3068) -5:PEGB1, pass, PUGB4
			10'd302 : rdata = 48'b110001110000001000000000000000000000000000001100;
			// PEs: 0 -> 1
			// srcs: (1004, 292)(3113) -6 --> (3113) -6:NI0, pass, PENB
			10'd303 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 56 -> 1
			// srcs: (1005, 294)(2378) -1 --> (2378) -1:PUNB, pass, PENB
			10'd304 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 24 -> 0
			// srcs: (1006, 297)(2493) -6 --> (2493) -6:PUGB3, pass, NI0
			10'd305 : rdata = 48'b110001110000011100000000000100000000000000000000;
			// PEs: 8 -> 1
			// srcs: (1007, 298)(2498) 13 --> (2498) 13:PUGB1, pass, PENB
			10'd306 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 4 -> 8
			// srcs: (1008, 318)(3098) -1 --> (3098) -1:PEGB4, pass, PUNB
			10'd307 : rdata = 48'b110001110000100000000000000000000000001000000000;
			// PEs: 1 -> 8
			// srcs: (1011, 319)(3116) -2 --> (3116) -2:PEGB1, pass, PUNB
			10'd308 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 1 -> 16
			// srcs: (1012, 320)(2379) 11 --> (2379) 11:PEGB1, pass, PUGB2
			10'd309 : rdata = 48'b110001110000001000000000000000000000000000001010;
			// PEs: 0 -> 1
			// srcs: (1013, 299)(2493) -6 --> (2493) -6:NI0, pass, PENB
			10'd310 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 24 -> 0
			// srcs: (1014, 304)(2665) -4 --> (2665) -4:PUGB3, pass, NI0
			10'd311 : rdata = 48'b110001110000011100000000000100000000000000000000;
			// PEs: 48 -> 1
			// srcs: (1015, 305)(2670) -10 --> (2670) -10:PUGB6, pass, PENB
			10'd312 : rdata = 48'b110001110000110100000000000000000000000100000000;
			// PEs: 0 -> 1
			// srcs: (1021, 306)(2665) -4 --> (2665) -4:NI0, pass, PENB
			10'd313 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 8 -> 0
			// srcs: (1022, 310)(2850) -4 --> (2850) -4:PUGB1, pass, NI0
			10'd314 : rdata = 48'b110001110000001100000000000100000000000000000000;
			// PEs: 24 -> 1
			// srcs: (1023, 311)(2855) 13 --> (2855) 13:PUGB3, pass, PENB
			10'd315 : rdata = 48'b110001110000011100000000000000000000000100000000;
			// PEs: 1 -> 40
			// srcs: (1028, 326)(2671) -14 --> (2671) -14:PEGB1, pass, PUGB5
			10'd316 : rdata = 48'b110001110000001000000000000000000000000000001101;
			// PEs: 0 -> 1
			// srcs: (1029, 312)(2850) -4 --> (2850) -4:NI0, pass, PENB
			10'd317 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 40 -> 0
			// srcs: (1030, 314)(2982) -2 --> (2982) -2:PUGB5, pass, NI0
			10'd318 : rdata = 48'b110001110000101100000000000100000000000000000000;
			// PEs: 16 -> 1
			// srcs: (1031, 315)(2987) -5 --> (2987) -5:PUGB2, pass, PENB
			10'd319 : rdata = 48'b110001110000010100000000000000000000000100000000;
			// PEs: 1 -> 40
			// srcs: (1036, 327)(2856) 9 --> (2856) 9:PEGB1, pass, PUGB5
			10'd320 : rdata = 48'b110001110000001000000000000000000000000000001101;
			// PEs: 0 -> 1
			// srcs: (1037, 316)(2982) -2 --> (2982) -2:NI0, pass, PENB
			10'd321 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 40 -> 1
			// srcs: (1038, 321)(2488) 11 --> (2488) 11:PUGB5, pass, PENB
			10'd322 : rdata = 48'b110001110000101100000000000000000000000100000000;
			// PEs: 24 -> 0
			// srcs: (1039, 322)(2536) -9 --> (2536) -9:PUGB3, pass, NI0
			10'd323 : rdata = 48'b110001110000011100000000000100000000000000000000;
			// PEs: 48 -> 1
			// srcs: (1040, 323)(2547) -12 --> (2547) -12:PUGB6, pass, PENB
			10'd324 : rdata = 48'b110001110000110100000000000000000000000100000000;
			// PEs: 0 -> 1
			// srcs: (1046, 324)(2536) -9 --> (2536) -9:NI0, pass, PENB
			10'd325 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 1 -> 32
			// srcs: (1053, 333)(2548) -21 --> (2548) -21:PEGB1, pass, PUGB4
			10'd326 : rdata = 48'b110001110000001000000000000000000000000000001100;
			// PEs: 32 -> 1
			// srcs: (1130, 328)(2977) -3 --> (2977) -3:PUGB4, pass, PENB
			10'd327 : rdata = 48'b110001110000100100000000000000000000000100000000;
			// PEs: 1 -> 56
			// srcs: (1138, 334)(2989) -10 --> (2989) -10:PEGB1, pass, PUGB7
			10'd328 : rdata = 48'b110001110000001000000000000000000000000000001111;
			// PEs: 8 -> 0
			// srcs: (1139, 329)(3099) 15 --> (3099) 15:PUGB1, pass, NI0
			10'd329 : rdata = 48'b110001110000001100000000000100000000000000000000;
			// PEs: 56 -> 7
			// srcs: (1162, 301)(2580) -21 --> (2580) -21:PUNB, pass, PEGB7
			10'd330 : rdata = 48'b110001101111111100000000000000000000000011110000;
			// PEs: 56 -> 1
			// srcs: (1163, 330)(3110) -12 --> (3110) -12:PUNB, pass, PENB
			10'd331 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 0 -> 1
			// srcs: (1169, 331)(3099) 15 --> (3099) 15:NI0, pass, PENB
			10'd332 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 7 -> 8
			// srcs: (1171, 325)(2586) -24 --> (2586) -24:PENB, pass, PUNB
			10'd333 : rdata = 48'b110001101111111000000000000000000000001000000000;
			// PEs: 56 -> 1
			// srcs: (1173, 332)(2477) 8 --> (2477) 8:PUNB, pass, PENB
			10'd334 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 1 -> 8
			// srcs: (1176, 338)(3111) 3 --> (3111) 3:PEGB1, pass, PUNB
			10'd335 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 1 -> 40
			// srcs: (1181, 339)(2501) 26 --> (2501) 26:PEGB1, pass, PUGB5
			10'd336 : rdata = 48'b110001110000001000000000000000000000000000001101;
			// PEs: 56 -> 0
			// srcs: (1415, 335)(3063) -28 --> (3063) -28:PUNB, pass, NI0
			10'd337 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 40 -> 1
			// srcs: (1416, 336)(3086) 0 --> (3086) 0:PUGB5, pass, PENB
			10'd338 : rdata = 48'b110001110000101100000000000000000000000100000000;
			// PEs: 0 -> 1
			// srcs: (1425, 337)(3063) -28 --> (3063) -28:NI0, pass, PENB
			10'd339 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 24 -> 0
			// srcs: (1430, 341)(2453) -10 --> (2453) -10:PUGB3, pass, NI0
			10'd340 : rdata = 48'b110001110000011100000000000100000000000000000000;
			// PEs: 40 -> 1
			// srcs: (1431, 342)(2550) 24 --> (2550) 24:PUGB5, pass, PENB
			10'd341 : rdata = 48'b110001110000101100000000000000000000000100000000;
			// PEs: 1 -> 8
			// srcs: (1432, 340)(3087) -28 --> (3087) -28:PEGB1, pass, PUNB
			10'd342 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 0 -> 1
			// srcs: (1437, 343)(2453) -10 --> (2453) -10:NI0, pass, PENB
			10'd343 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 56 -> 1
			// srcs: (1444, 344)(2746) 74 --> (2746) 74:PUNB, pass, PENB
			10'd344 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 1 -> 8
			// srcs: (1454, 345)(2747) 88 --> (2747) 88:PEGB1, pass, PUNB
			10'd345 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 8 -> 1
			// srcs: (1507, 346)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd346 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 2
			// srcs: (1511, 347)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd347 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 3
			// srcs: (1512, 348)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd348 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 4
			// srcs: (1513, 349)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd349 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 5
			// srcs: (1514, 350)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd350 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 6
			// srcs: (1515, 351)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd351 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 7
			// srcs: (1517, 352)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd352 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 1
			// srcs: (1567, 353)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd353 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 2
			// srcs: (1570, 354)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd354 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 3
			// srcs: (1573, 355)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd355 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 4
			// srcs: (1576, 356)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd356 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 5
			// srcs: (1579, 357)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd357 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 6
			// srcs: (1582, 358)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd358 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 7
			// srcs: (1585, 359)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd359 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 1
			// srcs: (1589, 360)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd360 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 2
			// srcs: (1590, 361)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd361 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 3
			// srcs: (1592, 362)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd362 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 4
			// srcs: (1593, 363)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd363 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 5
			// srcs: (1595, 364)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd364 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 6
			// srcs: (1596, 365)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd365 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 7
			// srcs: (1598, 366)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd366 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 1
			// srcs: (1669, 367)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd367 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 2
			// srcs: (1670, 368)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd368 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 3
			// srcs: (1672, 369)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd369 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 4
			// srcs: (1673, 370)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd370 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 5
			// srcs: (1675, 371)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd371 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 6
			// srcs: (1676, 372)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd372 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 7
			// srcs: (1678, 373)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd373 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 1
			// srcs: (1747, 374)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd374 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 2
			// srcs: (1750, 375)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd375 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 1
			// srcs: (1751, 376)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd376 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 2
			// srcs: (1752, 377)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd377 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 3
			// srcs: (1753, 378)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd378 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 3
			// srcs: (1754, 379)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd379 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 4
			// srcs: (1755, 380)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd380 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 5
			// srcs: (1756, 381)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd381 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 6
			// srcs: (1757, 382)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd382 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 7
			// srcs: (1758, 383)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd383 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 4
			// srcs: (1760, 384)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd384 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 5
			// srcs: (1763, 385)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd385 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 6
			// srcs: (1766, 386)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd386 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 7
			// srcs: (1769, 387)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd387 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 1
			// srcs: (1831, 388)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd388 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 2
			// srcs: (1832, 389)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd389 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 3
			// srcs: (1834, 390)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd390 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 4
			// srcs: (1835, 391)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd391 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 5
			// srcs: (1837, 392)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd392 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 6
			// srcs: (1838, 393)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd393 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 7
			// srcs: (1840, 394)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd394 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 1
			// srcs: (1911, 395)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd395 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 2
			// srcs: (1912, 396)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd396 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 3
			// srcs: (1914, 397)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd397 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 4
			// srcs: (1915, 398)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd398 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 5
			// srcs: (1917, 399)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd399 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 6
			// srcs: (1918, 400)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd400 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 7
			// srcs: (1920, 401)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd401 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 1
			// srcs: (1931, 402)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd402 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 2
			// srcs: (1934, 403)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd403 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 3
			// srcs: (1937, 404)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd404 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 4
			// srcs: (1940, 405)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd405 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 5
			// srcs: (1943, 406)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd406 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 6
			// srcs: (1946, 407)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd407 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 7
			// srcs: (1949, 408)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd408 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 1
			// srcs: (1993, 409)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd409 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 2
			// srcs: (1994, 410)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd410 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 3
			// srcs: (1996, 411)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd411 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 4
			// srcs: (1997, 412)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd412 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 5
			// srcs: (1999, 413)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd413 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 6
			// srcs: (2000, 414)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd414 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 7
			// srcs: (2001, 415)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd415 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 1
			// srcs: (2073, 416)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd416 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 2
			// srcs: (2074, 417)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd417 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 3
			// srcs: (2076, 418)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd418 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 4
			// srcs: (2077, 419)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd419 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 5
			// srcs: (2079, 420)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd420 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 6
			// srcs: (2080, 421)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd421 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 7
			// srcs: (2082, 422)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd422 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 1
			// srcs: (2115, 423)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd423 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 2
			// srcs: (2118, 424)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd424 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 3
			// srcs: (2121, 425)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd425 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 4
			// srcs: (2124, 426)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd426 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 5
			// srcs: (2127, 427)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd427 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 6
			// srcs: (2130, 428)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd428 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 7
			// srcs: (2133, 429)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd429 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 1
			// srcs: (2153, 430)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd430 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 2
			// srcs: (2154, 431)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd431 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 3
			// srcs: (2156, 432)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd432 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 4
			// srcs: (2157, 433)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd433 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 5
			// srcs: (2159, 434)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd434 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 6
			// srcs: (2160, 435)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd435 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 7
			// srcs: (2162, 436)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd436 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 1
			// srcs: (2235, 437)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd437 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 2
			// srcs: (2236, 438)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd438 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 3
			// srcs: (2238, 439)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd439 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 4
			// srcs: (2239, 440)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd440 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 5
			// srcs: (2241, 441)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd441 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 6
			// srcs: (2242, 442)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd442 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 7
			// srcs: (2244, 443)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd443 : rdata = 48'b110001110000001100000000000000000000000011110000;
			default : rdata = 48'b000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 1) begin
	always @(*) begin
		case(address)
			// PEs: 1, 1 -> 1
			// srcs: (1, 0)(4) -3, (789) -2 --> (1573) 6:ND0, NW0, *, NI0
			10'd0 : rdata = 48'b000110110000000001000000000100000000000000000000;
			// PEs: 1, 1 -> 0
			// srcs: (2, 1)(84) -3, (869) 0 --> (1653) 0:ND1, NW1, *, PEGB0
			10'd1 : rdata = 48'b000110110000000101000000001000000000000010000000;
			// PEs: 1, 1 -> 0
			// srcs: (3, 2)(164) -2, (949) -2 --> (1733) 4:ND2, NW2, *, PEGB0
			10'd2 : rdata = 48'b000110110000001001000000010000000000000010000000;
			// PEs: 1, 1 -> 0
			// srcs: (4, 3)(246) -3, (1031) 1 --> (1815) -3:ND3, NW3, *, PEGB0
			10'd3 : rdata = 48'b000110110000001101000000011000000000000010000000;
			// PEs: 1, 1 -> 0
			// srcs: (5, 4)(326) -2, (1111) 2 --> (1895) -4:ND4, NW4, *, PEGB0
			10'd4 : rdata = 48'b000110110000010001000000100000000000000010000000;
			// PEs: 1, 1 -> 0
			// srcs: (6, 5)(406) -2, (1191) 1 --> (1975) -2:ND5, NW5, *, PEGB0
			10'd5 : rdata = 48'b000110110000010101000000101000000000000010000000;
			// PEs: 1, 1 -> 0
			// srcs: (7, 6)(488) -1, (1273) 0 --> (2057) 0:ND6, NW6, *, PEGB0
			10'd6 : rdata = 48'b000110110000011001000000110000000000000010000000;
			// PEs: 1, 1 -> 0
			// srcs: (8, 7)(568) 1, (1353) 0 --> (2137) 0:ND7, NW7, *, PEGB0
			10'd7 : rdata = 48'b000110110000011101000000111000000000000010000000;
			// PEs: 1, 1 -> 4
			// srcs: (9, 8)(648) 2, (1433) 0 --> (2217) 0:ND8, NW8, *, PEGB4
			10'd8 : rdata = 48'b000110110000100001000001000000000000000011000000;
			// PEs: 1, 1 -> 6
			// srcs: (10, 9)(730) 1, (1515) 1 --> (2299) 1:ND9, NW9, *, PEGB6
			10'd9 : rdata = 48'b000110110000100101000001001000000000000011100000;
			// PEs: 1, 1 -> 0
			// srcs: (11, 10)(62) 0, (847) 0 --> (1631) 0:ND10, NW10, *, PEGB0
			10'd10 : rdata = 48'b000110110000101001000001010000000000000010000000;
			// PEs: 1, 1 -> 5
			// srcs: (12, 11)(242) -2, (1027) 0 --> (1811) 0:ND11, NW11, *, PEGB5
			10'd11 : rdata = 48'b000110110000101101000001011000000000000011010000;
			// PEs: 1, 1 -> 1
			// srcs: (13, 12)(426) 2, (1211) 2 --> (1995) 4:ND12, NW12, *, NI1
			10'd12 : rdata = 48'b000110110000110001000001100100001000000000000000;
			// PEs: 1, 1 -> 1
			// srcs: (14, 13)(610) -3, (1395) 1 --> (2179) -3:ND13, NW13, *, NI2
			10'd13 : rdata = 48'b000110110000110101000001101100010000000000000000;
			// PEs: 7, 0 -> 1
			// srcs: (33, 14)(1662) -3, (1663) -3 --> (2442) -6:PEGB7, PENB, +, NI3
			10'd14 : rdata = 48'b000011110000111011011111110100011000000000000000;
			// PEs: 7, 0 -> 1
			// srcs: (48, 15)(1742) 3, (1743) 1 --> (2521) 4:PEGB7, PENB, +, NI4
			10'd15 : rdata = 48'b000011110000111011011111110100100000000000000000;
			// PEs: 0 -> 
			// srcs: (54, 16)(1746) -2 --> (1746) -2:PENB, pass, 
			10'd16 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 0, 1 -> 1
			// srcs: (60, 17)(1745) 2, (1746) -2 --> (2526) 0:PENB, ALU, +, NI5
			10'd17 : rdata = 48'b000011101111111000111111111100101000000000000000;
			// PEs: 0 -> 
			// srcs: (78, 18)(1970) 2 --> (1970) 2:PENB, pass, 
			10'd18 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 0, 1 -> 1
			// srcs: (84, 19)(1969) -6, (1970) 2 --> (2751) -4:PENB, ALU, +, NI6
			10'd19 : rdata = 48'b000011101111111000111111111100110000000000000000;
			// PEs: 0 -> 
			// srcs: (86, 20)(1973) -6 --> (1973) -6:PENB, pass, 
			10'd20 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 0, 1 -> 6
			// srcs: (92, 21)(1972) -2, (1973) -6 --> (2754) -8:PENB, ALU, +, PEGB6
			10'd21 : rdata = 48'b000011101111111000111111111000000000000011100000;
			// PEs: 0 -> 
			// srcs: (94, 22)(2049) 0 --> (2049) 0:PENB, pass, 
			10'd22 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 0, 1 -> 1
			// srcs: (100, 23)(2048) 1, (2049) 0 --> (2827) 1:PENB, ALU, +, NI7
			10'd23 : rdata = 48'b000011101111111000111111111100111000000000000000;
			// PEs: 0 -> 1
			// srcs: (102, 24)(2052) 0 --> (2052) 0:PENB, pass, NI8
			10'd24 : rdata = 48'b110001101111111000000000000101000000000000000000;
			// PEs: 1 -> 0
			// srcs: (107, 36)(1573) 6 --> (1573) 6:NI0, pass, PEGB0
			10'd25 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 0, 1 -> 1
			// srcs: (108, 25)(2051) -4, (2052) 0 --> (2831) -4:PENB, NI8, +, NI0
			10'd26 : rdata = 48'b000011101111111010100001000100000000000000000000;
			// PEs: 0 -> 
			// srcs: (110, 26)(2055) 0 --> (2055) 0:PENB, pass, 
			10'd27 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 0, 1 -> 1
			// srcs: (116, 27)(2054) -6, (2055) 0 --> (2833) -6:PENB, ALU, +, NI8
			10'd28 : rdata = 48'b000011101111111000111111111101000000000000000000;
			// PEs: 0 -> 
			// srcs: (118, 28)(2129) 6 --> (2129) 6:PENB, pass, 
			10'd29 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 0, 1 -> 1
			// srcs: (124, 29)(2128) -4, (2129) 6 --> (2907) 2:PENB, ALU, +, NI9
			10'd30 : rdata = 48'b000011101111111000111111111101001000000000000000;
			// PEs: 0 -> 1
			// srcs: (126, 30)(2132) -2 --> (2132) -2:PENB, pass, NI10
			10'd31 : rdata = 48'b110001101111111000000000000101010000000000000000;
			// PEs: 1 -> 0
			// srcs: (131, 57)(2521) 4 --> (2521) 4:NI4, pass, PEGB0
			10'd32 : rdata = 48'b110001010000010000000000000000000000000010000000;
			// PEs: 0, 1 -> 1
			// srcs: (132, 31)(2131) 2, (2132) -2 --> (2910) 0:PENB, NI10, +, NI4
			10'd33 : rdata = 48'b000011101111111010100001010100100000000000000000;
			// PEs: 0 -> 
			// srcs: (134, 32)(2135) -3 --> (2135) -3:PENB, pass, 
			10'd34 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 0, 1 -> 1
			// srcs: (140, 33)(2134) 2, (2135) -3 --> (2912) -1:PENB, ALU, +, NI10
			10'd35 : rdata = 48'b000011101111111000111111111101010000000000000000;
			// PEs: 0 -> 1
			// srcs: (142, 34)(2215) 2 --> (2215) 2:PENB, pass, NI11
			10'd36 : rdata = 48'b110001101111111000000000000101011000000000000000;
			// PEs: 1 -> 0
			// srcs: (146, 58)(2526) 0 --> (2526) 0:NI5, pass, PEGB0
			10'd37 : rdata = 48'b110001010000010100000000000000000000000010000000;
			// PEs: 1 -> 0
			// srcs: (147, 71)(1995) 4 --> (1995) 4:NI1, pass, PEGB0
			10'd38 : rdata = 48'b110001010000000100000000000000000000000010000000;
			// PEs: 0, 1 -> 1
			// srcs: (148, 35)(2214) -3, (2215) 2 --> (2994) -1:PENB, NI11, +, NI1
			10'd39 : rdata = 48'b000011101111111010100001011100001000000000000000;
			// PEs: 1 -> 0
			// srcs: (162, 79)(2831) -4 --> (2831) -4:NI0, pass, PEGB0
			10'd40 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 1 -> 0
			// srcs: (167, 82)(2910) 0 --> (2910) 0:NI4, pass, PEGB0
			10'd41 : rdata = 48'b110001010000010000000000000000000000000010000000;
			// PEs: 1 -> 0
			// srcs: (174, 80)(2833) -6 --> (2833) -6:NI8, pass, PEGB0
			10'd42 : rdata = 48'b110001010000100000000000000000000000000010000000;
			// PEs: 1 -> 0
			// srcs: (175, 83)(2912) -1 --> (2912) -1:NI10, pass, PEGB0
			10'd43 : rdata = 48'b110001010000101000000000000000000000000010000000;
			// PEs: 1 -> 0
			// srcs: (179, 49)(2442) -6 --> (2442) -6:NI3, pass, PEGB0
			10'd44 : rdata = 48'b110001010000001100000000000000000000000010000000;
			// PEs: 1 -> 0
			// srcs: (183, 84)(2179) -3 --> (2179) -3:NI2, pass, PEGB0
			10'd45 : rdata = 48'b110001010000001000000000000000000000000010000000;
			// PEs: 1 -> 0
			// srcs: (203, 68)(2751) -4 --> (2751) -4:NI6, pass, PEGB0
			10'd46 : rdata = 48'b110001010000011000000000000000000000000010000000;
			// PEs: 0 -> 
			// srcs: (218, 37)(1968) 0 --> (1968) 0:PENB, pass, 
			10'd47 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 0, 1 -> 1
			// srcs: (224, 38)(1967) 0, (1968) 0 --> (2749) 0:PENB, ALU, +, NI0
			10'd48 : rdata = 48'b000011101111111000111111111100000000000000000000;
			// PEs: 1 -> 0
			// srcs: (229, 78)(2827) 1 --> (2827) 1:NI7, pass, PEGB0
			10'd49 : rdata = 48'b110001010000011100000000000000000000000010000000;
			// PEs: 1 -> 0
			// srcs: (237, 81)(2907) 2 --> (2907) 2:NI9, pass, PEGB0
			10'd50 : rdata = 48'b110001010000100100000000000000000000000010000000;
			// PEs: 0 -> 1
			// srcs: (243, 39)(2211) -1 --> (2211) -1:PENB, pass, NI2
			10'd51 : rdata = 48'b110001101111111000000000000100010000000000000000;
			// PEs: 1 -> 0
			// srcs: (245, 88)(2994) -1 --> (2994) -1:NI1, pass, PEGB0
			10'd52 : rdata = 48'b110001010000000100000000000000000000000010000000;
			// PEs: 0, 1 -> 1
			// srcs: (249, 40)(2210) -1, (2211) -1 --> (2991) -2:PENB, NI2, +, NI1
			10'd53 : rdata = 48'b000011101111111010100000010100001000000000000000;
			// PEs: 0 -> 
			// srcs: (251, 41)(2213) 0 --> (2213) 0:PENB, pass, 
			10'd54 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 0, 1 -> 2
			// srcs: (257, 42)(2212) 0, (2213) 0 --> (2992) 0:PENB, ALU, +, PENB
			10'd55 : rdata = 48'b000011101111111000111111111000000000000100000000;
			// PEs: 0 -> 1
			// srcs: (259, 43)(1579) -6 --> (1579) -6:PENB, pass, NI2
			10'd56 : rdata = 48'b110001101111111000000000000100010000000000000000;
			// PEs: 1 -> 2
			// srcs: (264, 87)(2991) -2 --> (2991) -2:NI1, pass, PENB
			10'd57 : rdata = 48'b110001010000000100000000000000000000000100000000;
			// PEs: 0, 1 -> 0
			// srcs: (265, 44)(2360) -10, (1579) -6 --> (2361) -16:PENB, NI2, +, PEGB0
			10'd58 : rdata = 48'b000011101111111010100000010000000000000010000000;
			// PEs: 2, 0 -> 0
			// srcs: (266, 45)(2363) -5, (1582) -6 --> (2364) -11:PEGB2, PENB, +, PEGB0
			10'd59 : rdata = 48'b000011110000010011011111110000000000000010000000;
			// PEs: 0 -> 
			// srcs: (268, 46)(1612) 0 --> (1612) 0:PENB, pass, 
			10'd60 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 0, 1 -> 1
			// srcs: (274, 47)(2392) -8, (1612) 0 --> (2393) -8:PENB, ALU, +, NI1
			10'd61 : rdata = 48'b000011101111111000111111111100001000000000000000;
			// PEs: 0, 5 -> 0
			// srcs: (275, 48)(2422) -5, (1643) 2 --> (2423) -3:PENB, PEGB5, +, PEGB0
			10'd62 : rdata = 48'b000011101111111011100001010000000000000010000000;
			// PEs: 0 -> 
			// srcs: (277, 50)(1683) 1 --> (1683) 1:PENB, pass, 
			10'd63 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 0, 1 -> 0
			// srcs: (283, 51)(2462) 1, (1683) 1 --> (2463) 2:PENB, ALU, +, PEGB0
			10'd64 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 0 -> 
			// srcs: (285, 52)(1704) -2 --> (1704) -2:PENB, pass, 
			10'd65 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 0, 1 -> 0
			// srcs: (291, 53)(2483) -1, (1704) -2 --> (2484) -3:PENB, ALU, +, PEGB0
			10'd66 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 0 -> 
			// srcs: (293, 54)(1716) -2 --> (1716) -2:PENB, pass, 
			10'd67 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 0, 1 -> 0
			// srcs: (299, 55)(2494) 7, (1716) -2 --> (2495) 5:PENB, ALU, +, PEGB0
			10'd68 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 0, 2 -> 0
			// srcs: (300, 56)(2502) 7, (2503) -6 --> (2504) 1:PENB, PEGB2, +, PEGB0
			10'd69 : rdata = 48'b000011101111111011100000100000000000000010000000;
			// PEs: 5, 0 -> 1
			// srcs: (301, 59)(2583) -4, (1805) 0 --> (2584) -4:PEGB5, PENB, +, NI2
			10'd70 : rdata = 48'b000011110000101011011111110100010000000000000000;
			// PEs: 6, 0 -> 3
			// srcs: (527, 60)(2587) 8, (1808) 0 --> (2588) 8:PEGB6, PENB, +, PEGB3
			10'd71 : rdata = 48'b000011110000110011011111110000000000000010110000;
			// PEs: 0 -> 
			// srcs: (529, 61)(1851) 0 --> (1851) 0:PENB, pass, 
			10'd72 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 0, 1 -> 0
			// srcs: (535, 62)(2629) 3, (1851) 0 --> (2630) 3:PENB, ALU, +, PEGB0
			10'd73 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 0 -> 
			// srcs: (537, 63)(1885) -2 --> (1885) -2:PENB, pass, 
			10'd74 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 0, 1 -> 0
			// srcs: (543, 64)(2663) -2, (1885) -2 --> (2664) -4:PENB, ALU, +, PEGB0
			10'd75 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 0 -> 
			// srcs: (545, 65)(1903) 3 --> (1903) 3:PENB, pass, 
			10'd76 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 0, 1 -> 0
			// srcs: (551, 66)(2680) -8, (1903) 3 --> (2681) -5:PENB, ALU, +, PEGB0
			10'd77 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 0, 1 -> 0
			// srcs: (552, 67)(2748) -1, (2749) 0 --> (2750) -1:PENB, NI0, +, PEGB0
			10'd78 : rdata = 48'b000011101111111010100000000000000000000010000000;
			// PEs: 0 -> 
			// srcs: (555, 69)(1986) 0 --> (1986) 0:PENB, pass, 
			10'd79 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 0, 1 -> 0
			// srcs: (561, 70)(2765) -4, (1986) 0 --> (2766) -4:PENB, ALU, +, PEGB0
			10'd80 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 0 -> 
			// srcs: (563, 72)(2020) 1 --> (2020) 1:PENB, pass, 
			10'd81 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 0, 1 -> 0
			// srcs: (569, 73)(2799) -2, (2020) 1 --> (2800) -1:PENB, ALU, +, PEGB0
			10'd82 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 0 -> 
			// srcs: (571, 74)(2029) 0 --> (2029) 0:PENB, pass, 
			10'd83 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 0, 1 -> 0
			// srcs: (577, 75)(2808) -6, (2029) 0 --> (2809) -6:PENB, ALU, +, PEGB0
			10'd84 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 0 -> 
			// srcs: (579, 76)(2038) -2 --> (2038) -2:PENB, pass, 
			10'd85 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 0, 1 -> 0
			// srcs: (585, 77)(2815) -1, (2038) -2 --> (2816) -3:PENB, ALU, +, PEGB0
			10'd86 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 0 -> 
			// srcs: (587, 85)(2209) 0 --> (2209) 0:PENB, pass, 
			10'd87 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 0, 1 -> 0
			// srcs: (593, 86)(2985) -2, (2209) 0 --> (2986) -2:PENB, ALU, +, PEGB0
			10'd88 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 6, 0 -> 0
			// srcs: (601, 89)(3077) -2, (2301) 0 --> (3078) -2:PEGB6, PENB, +, PEGB0
			10'd89 : rdata = 48'b000011110000110011011111110000000000000010000000;
			// PEs: 0 -> 
			// srcs: (602, 90)(2320) 0 --> (2320) 0:PENB, pass, 
			10'd90 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 0, 1 -> 4
			// srcs: (607, 91)(3096) 2, (2320) 0 --> (3097) 2:PENB, ALU, +, PEGB4
			10'd91 : rdata = 48'b000011101111111000111111111000000000000011000000;
			// PEs: 0 -> 
			// srcs: (609, 92)(2344) 0 --> (2344) 0:PENB, pass, 
			10'd92 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 0, 1 -> 0
			// srcs: (615, 93)(3119) -4, (2344) 0 --> (3120) -4:PENB, ALU, +, PEGB0
			10'd93 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 0 -> 
			// srcs: (617, 94)(2372) 11 --> (2372) 11:PENB, pass, 
			10'd94 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 0, 1 -> 1
			// srcs: (623, 95)(2370) 1, (2372) 11 --> (2373) 12:PENB, ALU, +, NI0
			10'd95 : rdata = 48'b000011101111111000111111111100000000000000000000;
			// PEs: 1, 0 -> 0
			// srcs: (624, 96)(2393) -8, (2395) 6 --> (2396) -2:NI1, PENB, +, PEGB0
			10'd96 : rdata = 48'b000011010000000111011111110000000000000010000000;
			// PEs: 0 -> 
			// srcs: (626, 97)(2474) -3 --> (2474) -3:PENB, pass, 
			10'd97 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 0, 1 -> 0
			// srcs: (632, 98)(2472) 15, (2474) -3 --> (2475) 12:PENB, ALU, +, PEGB0
			10'd98 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 0 -> 
			// srcs: (634, 99)(2522) 5 --> (2522) 5:PENB, pass, 
			10'd99 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 0, 1 -> 0
			// srcs: (640, 100)(2520) -1, (2522) 5 --> (2523) 4:PENB, ALU, +, PEGB0
			10'd100 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 0, 1 -> 7
			// srcs: (952, 101)(2582) 1, (2584) -4 --> (2585) -3:PENB, NI2, +, PEGB7
			10'd101 : rdata = 48'b000011101111111010100000010000000000000011110000;
			// PEs: 0 -> 
			// srcs: (954, 102)(2627) 6 --> (2627) 6:PENB, pass, 
			10'd102 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 0, 1 -> 0
			// srcs: (960, 103)(2625) 10, (2627) 6 --> (2628) 16:PENB, ALU, +, PEGB0
			10'd103 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 0 -> 
			// srcs: (962, 104)(2687) -7 --> (2687) -7:PENB, pass, 
			10'd104 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 0, 1 -> 0
			// srcs: (968, 105)(2685) 4, (2687) -7 --> (2688) -3:PENB, ALU, +, PEGB0
			10'd105 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 6, 0 -> 0
			// srcs: (976, 106)(2755) -2, (2757) -5 --> (2758) -7:PEGB6, PENB, +, PEGB0
			10'd106 : rdata = 48'b000011110000110011011111110000000000000010000000;
			// PEs: 0 -> 
			// srcs: (977, 107)(2834) -6 --> (2834) -6:PENB, pass, 
			10'd107 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 0, 1 -> 0
			// srcs: (982, 108)(2832) 0, (2834) -6 --> (2835) -6:PENB, ALU, +, PEGB0
			10'd108 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 0 -> 
			// srcs: (984, 109)(2952) 4 --> (2952) 4:PENB, pass, 
			10'd109 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 0, 1 -> 0
			// srcs: (990, 110)(2950) -8, (2952) 4 --> (2953) -4:PENB, ALU, +, PEGB0
			10'd110 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 0 -> 
			// srcs: (992, 111)(3067) -2 --> (3067) -2:PENB, pass, 
			10'd111 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 0, 1 -> 0
			// srcs: (998, 112)(3065) -3, (3067) -2 --> (3068) -5:PENB, ALU, +, PEGB0
			10'd112 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 0 -> 
			// srcs: (1000, 113)(3115) 4 --> (3115) 4:PENB, pass, 
			10'd113 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 0, 1 -> 0
			// srcs: (1006, 114)(3113) -6, (3115) 4 --> (3116) -2:PENB, ALU, +, PEGB0
			10'd114 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 1, 0 -> 0
			// srcs: (1007, 115)(2373) 12, (2378) -1 --> (2379) 11:NI0, PENB, +, PEGB0
			10'd115 : rdata = 48'b000011010000000011011111110000000000000010000000;
			// PEs: 0 -> 
			// srcs: (1009, 116)(2498) 13 --> (2498) 13:PENB, pass, 
			10'd116 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 0, 1 -> 1
			// srcs: (1015, 117)(2493) -6, (2498) 13 --> (2499) 7:PENB, ALU, +, NI0
			10'd117 : rdata = 48'b000011101111111000111111111100000000000000000000;
			// PEs: 0 -> 
			// srcs: (1017, 118)(2670) -10 --> (2670) -10:PENB, pass, 
			10'd118 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 0, 1 -> 0
			// srcs: (1023, 119)(2665) -4, (2670) -10 --> (2671) -14:PENB, ALU, +, PEGB0
			10'd119 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 0 -> 
			// srcs: (1025, 120)(2855) 13 --> (2855) 13:PENB, pass, 
			10'd120 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 0, 1 -> 0
			// srcs: (1031, 121)(2850) -4, (2855) 13 --> (2856) 9:PENB, ALU, +, PEGB0
			10'd121 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 0 -> 
			// srcs: (1033, 122)(2987) -5 --> (2987) -5:PENB, pass, 
			10'd122 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 0, 1 -> 1
			// srcs: (1039, 123)(2982) -2, (2987) -5 --> (2988) -7:PENB, ALU, +, NI1
			10'd123 : rdata = 48'b000011101111111000111111111100001000000000000000;
			// PEs: 0, 1 -> 1
			// srcs: (1040, 124)(2488) 11, (2499) 7 --> (2500) 18:PENB, NI0, +, NI2
			10'd124 : rdata = 48'b000011101111111010100000000100010000000000000000;
			// PEs: 0 -> 
			// srcs: (1042, 125)(2547) -12 --> (2547) -12:PENB, pass, 
			10'd125 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 0, 1 -> 0
			// srcs: (1048, 126)(2536) -9, (2547) -12 --> (2548) -21:PENB, ALU, +, PEGB0
			10'd126 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 0, 1 -> 0
			// srcs: (1133, 127)(2977) -3, (2988) -7 --> (2989) -10:PENB, NI1, +, PEGB0
			10'd127 : rdata = 48'b000011101111111010100000001000000000000010000000;
			// PEs: 0 -> 
			// srcs: (1165, 128)(3110) -12 --> (3110) -12:PENB, pass, 
			10'd128 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 0, 1 -> 0
			// srcs: (1171, 129)(3099) 15, (3110) -12 --> (3111) 3:PENB, ALU, +, PEGB0
			10'd129 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 0, 1 -> 0
			// srcs: (1176, 130)(2477) 8, (2500) 18 --> (2501) 26:PENB, NI2, +, PEGB0
			10'd130 : rdata = 48'b000011101111111010100000010000000000000010000000;
			// PEs: 0 -> 
			// srcs: (1418, 131)(3086) 0 --> (3086) 0:PENB, pass, 
			10'd131 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 0, 1 -> 0
			// srcs: (1427, 132)(3063) -28, (3086) 0 --> (3087) -28:PENB, ALU, +, PEGB0
			10'd132 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 0 -> 
			// srcs: (1433, 133)(2550) 24 --> (2550) 24:PENB, pass, 
			10'd133 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 0, 1 -> 
			// srcs: (1439, 134)(2453) -10, (2550) 24 --> (2551) 14:PENB, ALU, +, 
			10'd134 : rdata = 48'b000011101111111000111111111000000000000000000000;
			// PEs: 1, 0 -> 0
			// srcs: (1449, 135)(2551) 14, (2746) 74 --> (2747) 88:ALU, PENB, +, PEGB0
			10'd135 : rdata = 48'b000010011111111111011111110000000000000010000000;
			// PEs: 0, 1 -> 2
			// srcs: (1510, 136)(3140) 47, (4) -3 --> (3141) -141:PENB, ND0, *, PENB
			10'd136 : rdata = 48'b000111101111111001100000000000000000000100000000;
			// PEs: 1, 2 -> 1
			// srcs: (1519, 150)(789) -2, (3925) -141 --> (4709) 139:NW0, PEGB2, -, NW0
			10'd137 : rdata = 48'b000100100000000011100000100000000100000000000000;
			// PEs: 0, 1 -> 2
			// srcs: (1569, 137)(3140) 47, (62) 0 --> (3199) 0:PENB, ND10, *, PENB
			10'd138 : rdata = 48'b000111101111111001100001010000000000000100000000;
			// PEs: 1, 2 -> 1
			// srcs: (1578, 151)(847) 0, (3983) 0 --> (4767) 0:NW10, PEGB2, -, NW10
			10'd139 : rdata = 48'b000100100000101011100000100000000110100000000000;
			// PEs: 0, 1 -> 2
			// srcs: (1591, 138)(3140) 47, (84) -3 --> (3221) -141:PENB, ND1, *, PENB
			10'd140 : rdata = 48'b000111101111111001100000001000000000000100000000;
			// PEs: 1, 2 -> 1
			// srcs: (1600, 152)(869) 0, (4005) -141 --> (4789) 141:NW1, PEGB2, -, NW1
			10'd141 : rdata = 48'b000100100000000111100000100000000100010000000000;
			// PEs: 0, 1 -> 2
			// srcs: (1671, 139)(3140) 47, (164) -2 --> (3301) -94:PENB, ND2, *, PENB
			10'd142 : rdata = 48'b000111101111111001100000010000000000000100000000;
			// PEs: 1, 2 -> 1
			// srcs: (1680, 153)(949) -2, (4085) -94 --> (4869) 92:NW2, PEGB2, -, NW2
			10'd143 : rdata = 48'b000100100000001011100000100000000100100000000000;
			// PEs: 0, 1 -> 2
			// srcs: (1749, 140)(3140) 47, (242) -2 --> (3379) -94:PENB, ND11, *, PENB
			10'd144 : rdata = 48'b000111101111111001100001011000000000000100000000;
			// PEs: 0, 1 -> 2
			// srcs: (1753, 141)(3140) 47, (246) -3 --> (3383) -141:PENB, ND3, *, PENB
			10'd145 : rdata = 48'b000111101111111001100000011000000000000100000000;
			// PEs: 1, 2 -> 1
			// srcs: (1758, 154)(1027) 0, (4163) -94 --> (4947) 94:NW11, PEGB2, -, NW11
			10'd146 : rdata = 48'b000100100000101111100000100000000110110000000000;
			// PEs: 1, 2 -> 1
			// srcs: (1762, 155)(1031) 1, (4167) -141 --> (4951) 142:NW3, PEGB2, -, NW3
			10'd147 : rdata = 48'b000100100000001111100000100000000100110000000000;
			// PEs: 0, 1 -> 2
			// srcs: (1833, 142)(3140) 47, (326) -2 --> (3463) -94:PENB, ND4, *, PENB
			10'd148 : rdata = 48'b000111101111111001100000100000000000000100000000;
			// PEs: 1, 2 -> 1
			// srcs: (1842, 156)(1111) 2, (4247) -94 --> (5031) 96:NW4, PEGB2, -, NW4
			10'd149 : rdata = 48'b000100100000010011100000100000000101000000000000;
			// PEs: 0, 1 -> 2
			// srcs: (1913, 143)(3140) 47, (406) -2 --> (3543) -94:PENB, ND5, *, PENB
			10'd150 : rdata = 48'b000111101111111001100000101000000000000100000000;
			// PEs: 1, 2 -> 1
			// srcs: (1922, 157)(1191) 1, (4327) -94 --> (5111) 95:NW5, PEGB2, -, NW5
			10'd151 : rdata = 48'b000100100000010111100000100000000101010000000000;
			// PEs: 0, 1 -> 2
			// srcs: (1933, 144)(3140) 47, (426) 2 --> (3563) 94:PENB, ND12, *, PENB
			10'd152 : rdata = 48'b000111101111111001100001100000000000000100000000;
			// PEs: 1, 2 -> 1
			// srcs: (1942, 158)(1211) 2, (4347) 94 --> (5131) -92:NW12, PEGB2, -, NW12
			10'd153 : rdata = 48'b000100100000110011100000100000000111000000000000;
			// PEs: 0, 1 -> 2
			// srcs: (1995, 145)(3140) 47, (488) -1 --> (3625) -47:PENB, ND6, *, PENB
			10'd154 : rdata = 48'b000111101111111001100000110000000000000100000000;
			// PEs: 1, 2 -> 1
			// srcs: (2004, 159)(1273) 0, (4409) -47 --> (5193) 47:NW6, PEGB2, -, NW6
			10'd155 : rdata = 48'b000100100000011011100000100000000101100000000000;
			// PEs: 0, 1 -> 2
			// srcs: (2075, 146)(3140) 47, (568) 1 --> (3705) 47:PENB, ND7, *, PENB
			10'd156 : rdata = 48'b000111101111111001100000111000000000000100000000;
			// PEs: 1, 2 -> 1
			// srcs: (2084, 160)(1353) 0, (4489) 47 --> (5273) -47:NW7, PEGB2, -, NW7
			10'd157 : rdata = 48'b000100100000011111100000100000000101110000000000;
			// PEs: 0, 1 -> 2
			// srcs: (2117, 147)(3140) 47, (610) -3 --> (3747) -141:PENB, ND13, *, PENB
			10'd158 : rdata = 48'b000111101111111001100001101000000000000100000000;
			// PEs: 1, 2 -> 1
			// srcs: (2126, 161)(1395) 1, (4531) -141 --> (5315) 142:NW13, PEGB2, -, NW13
			10'd159 : rdata = 48'b000100100000110111100000100000000111010000000000;
			// PEs: 0, 1 -> 2
			// srcs: (2155, 148)(3140) 47, (648) 2 --> (3785) 94:PENB, ND8, *, PENB
			10'd160 : rdata = 48'b000111101111111001100001000000000000000100000000;
			// PEs: 1, 2 -> 1
			// srcs: (2164, 162)(1433) 0, (4569) 94 --> (5353) -94:NW8, PEGB2, -, NW8
			10'd161 : rdata = 48'b000100100000100011100000100000000110000000000000;
			// PEs: 0, 1 -> 2
			// srcs: (2237, 149)(3140) 47, (730) 1 --> (3867) 47:PENB, ND9, *, PENB
			10'd162 : rdata = 48'b000111101111111001100001001000000000000100000000;
			// PEs: 1, 2 -> 1
			// srcs: (2246, 163)(1515) 1, (4651) 47 --> (5435) -46:NW9, PEGB2, -, NW9
			10'd163 : rdata = 48'b000100100000100111100000100000000110010000000000;
			default : rdata = 48'b000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 2) begin
	always @(*) begin
		case(address)
			// PEs: 2, 2 -> 2
			// srcs: (1, 0)(5) -1, (790) -3 --> (1574) 3:ND0, NW0, *, NI0
			10'd0 : rdata = 48'b000110110000000001000000000100000000000000000000;
			// PEs: 2, 2 -> 0
			// srcs: (2, 1)(85) 2, (870) -2 --> (1654) -4:ND1, NW1, *, PEGB0
			10'd1 : rdata = 48'b000110110000000101000000001000000000000010000000;
			// PEs: 2, 2 -> 0
			// srcs: (3, 2)(165) -1, (950) 1 --> (1734) -1:ND2, NW2, *, PEGB0
			10'd2 : rdata = 48'b000110110000001001000000010000000000000010000000;
			// PEs: 2, 2 -> 0
			// srcs: (4, 3)(247) 0, (1032) -1 --> (1816) 0:ND3, NW3, *, PEGB0
			10'd3 : rdata = 48'b000110110000001101000000011000000000000010000000;
			// PEs: 2, 2 -> 0
			// srcs: (5, 4)(327) 1, (1112) -3 --> (1896) -3:ND4, NW4, *, PEGB0
			10'd4 : rdata = 48'b000110110000010001000000100000000000000010000000;
			// PEs: 2, 2 -> 0
			// srcs: (6, 5)(407) 1, (1192) -3 --> (1976) -3:ND5, NW5, *, PEGB0
			10'd5 : rdata = 48'b000110110000010101000000101000000000000010000000;
			// PEs: 2, 2 -> 0
			// srcs: (7, 6)(489) 1, (1274) 0 --> (2058) 0:ND6, NW6, *, PEGB0
			10'd6 : rdata = 48'b000110110000011001000000110000000000000010000000;
			// PEs: 2, 2 -> 0
			// srcs: (8, 7)(569) 0, (1354) -1 --> (2138) 0:ND7, NW7, *, PEGB0
			10'd7 : rdata = 48'b000110110000011101000000111000000000000010000000;
			// PEs: 2, 2 -> 4
			// srcs: (9, 8)(649) -1, (1434) -1 --> (2218) 1:ND8, NW8, *, PEGB4
			10'd8 : rdata = 48'b000110110000100001000001000000000000000011000000;
			// PEs: 2, 2 -> 6
			// srcs: (10, 9)(731) 1, (1516) -3 --> (2300) -3:ND9, NW9, *, PEGB6
			10'd9 : rdata = 48'b000110110000100101000001001000000000000011100000;
			// PEs: 2, 2 -> 2
			// srcs: (11, 10)(65) -3, (850) -1 --> (1634) 3:ND10, NW10, *, NI1
			10'd10 : rdata = 48'b000110110000101001000001010100001000000000000000;
			// PEs: 2, 2 -> 2
			// srcs: (12, 11)(245) 2, (1030) -3 --> (1814) -6:ND11, NW11, *, NI2
			10'd11 : rdata = 48'b000110110000101101000001011100010000000000000000;
			// PEs: 2, 2 -> 2
			// srcs: (13, 12)(429) 0, (1214) 2 --> (1998) 0:ND12, NW12, *, NI3
			10'd12 : rdata = 48'b000110110000110001000001100100011000000000000000;
			// PEs: 2, 2 -> 2
			// srcs: (14, 13)(613) -3, (1398) 1 --> (2182) -3:ND13, NW13, *, NI4
			10'd13 : rdata = 48'b000110110000110101000001101100100000000000000000;
			// PEs: 0 -> 
			// srcs: (16, 14)(1581) 1 --> (1581) 1:PEGB0, pass, 
			10'd14 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 7, 2 -> 1
			// srcs: (19, 15)(1580) -6, (1581) 1 --> (2363) -5:PEGB7, ALU, +, PEGB1
			10'd15 : rdata = 48'b000011110000111000111111111000000000000010010000;
			// PEs: 0 -> 
			// srcs: (37, 16)(1725) 6 --> (1725) 6:PEGB0, pass, 
			10'd16 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 0, 2 -> 2
			// srcs: (46, 17)(1724) 2, (1725) 6 --> (2505) 8:PEGB0, ALU, +, NI5
			10'd17 : rdata = 48'b000011110000000000111111111100101000000000000000;
			// PEs: 0 -> 
			// srcs: (67, 18)(1890) -2 --> (1890) -2:PEGB0, pass, 
			10'd18 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 0, 2 -> 2
			// srcs: (76, 19)(1889) 0, (1890) -2 --> (2668) -2:PEGB0, ALU, +, NI6
			10'd19 : rdata = 48'b000011110000000000111111111100110000000000000000;
			// PEs: 2 -> 0
			// srcs: (115, 20)(1574) 3 --> (1574) 3:NI0, pass, PEGB0
			10'd20 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (137, 24)(2505) 8 --> (2505) 8:NI5, pass, PEGB0
			10'd21 : rdata = 48'b110001010000010100000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (147, 26)(2668) -2 --> (2668) -2:NI6, pass, PEGB0
			10'd22 : rdata = 48'b110001010000011000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (159, 28)(2182) -3 --> (2182) -3:NI4, pass, PEGB0
			10'd23 : rdata = 48'b110001010000010000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (171, 23)(1634) 3 --> (1634) 3:NI1, pass, PEGB0
			10'd24 : rdata = 48'b110001010000000100000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (187, 25)(1814) -6 --> (1814) -6:NI2, pass, PEGB0
			10'd25 : rdata = 48'b110001010000001000000000000000000000000010000000;
			// PEs: 2 -> 0
			// srcs: (211, 27)(1998) 0 --> (1998) 0:NI3, pass, PEGB0
			10'd26 : rdata = 48'b110001010000001100000000000000000000000010000000;
			// PEs: 0 -> 
			// srcs: (219, 21)(1723) 0 --> (1723) 0:PEGB0, pass, 
			10'd27 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 0, 2 -> 1
			// srcs: (228, 22)(1722) -6, (1723) 0 --> (2503) -6:PEGB0, ALU, +, PEGB1
			10'd28 : rdata = 48'b000011110000000000111111111000000000000010010000;
			// PEs: 1 -> 
			// srcs: (259, 29)(2992) 0 --> (2992) 0:PENB, pass, 
			10'd29 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 1, 2 -> 0
			// srcs: (266, 30)(2991) -2, (2992) 0 --> (2993) -2:PENB, ALU, +, PEGB0
			10'd30 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 2, 1 -> 1
			// srcs: (1513, 45)(3) 1, (3141) -141 --> (3925) -141:NM0, PENB, *, PEGB1
			10'd31 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 0, 2 -> 3
			// srcs: (1516, 31)(3140) 47, (5) -1 --> (3142) -47:PEGB0, ND0, *, PENB
			10'd32 : rdata = 48'b000111110000000001100000000000000000000100000000;
			// PEs: 2, 3 -> 2
			// srcs: (1525, 63)(790) -3, (3926) -47 --> (4710) 44:NW0, PEGB3, -, NW0
			10'd33 : rdata = 48'b000100100000000011100000110000000100000000000000;
			// PEs: 2, 1 -> 1
			// srcs: (1572, 46)(3) 1, (3199) 0 --> (3983) 0:NM0, PENB, *, PEGB1
			10'd34 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 0, 2 -> 
			// srcs: (1575, 32)(3140) 47, (65) -3 --> (3202) -141:PEGB0, ND10, *, 
			10'd35 : rdata = 48'b000111110000000001100001010000000000000000000000;
			// PEs: 2, 2 -> 
			// srcs: (1578, 47)(3) 1, (3202) -141 --> (3986) -141:NM0, ALU, *, 
			10'd36 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 2, 2 -> 2
			// srcs: (1581, 64)(850) -1, (3986) -141 --> (4770) 140:NW10, ALU, -, NW10
			10'd37 : rdata = 48'b000100100000101000111111111000000110100000000000;
			// PEs: 2, 1 -> 1
			// srcs: (1594, 48)(3) 1, (3221) -141 --> (4005) -141:NM0, PENB, *, PEGB1
			10'd38 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 0, 2 -> 3
			// srcs: (1595, 33)(3140) 47, (85) 2 --> (3222) 94:PEGB0, ND1, *, PENB
			10'd39 : rdata = 48'b000111110000000001100000001000000000000100000000;
			// PEs: 2, 3 -> 2
			// srcs: (1604, 65)(870) -2, (4006) 94 --> (4790) -96:NW1, PEGB3, -, NW1
			10'd40 : rdata = 48'b000100100000000111100000110000000100010000000000;
			// PEs: 2, 1 -> 1
			// srcs: (1674, 49)(3) 1, (3301) -94 --> (4085) -94:NM0, PENB, *, PEGB1
			10'd41 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 0, 2 -> 3
			// srcs: (1675, 34)(3140) 47, (165) -1 --> (3302) -47:PEGB0, ND2, *, PENB
			10'd42 : rdata = 48'b000111110000000001100000010000000000000100000000;
			// PEs: 2, 3 -> 2
			// srcs: (1684, 66)(950) 1, (4086) -47 --> (4870) 48:NW2, PEGB3, -, NW2
			10'd43 : rdata = 48'b000100100000001011100000110000000100100000000000;
			// PEs: 2, 1 -> 1
			// srcs: (1752, 50)(3) 1, (3379) -94 --> (4163) -94:NM0, PENB, *, PEGB1
			10'd44 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 0, 2 -> 2
			// srcs: (1755, 35)(3140) 47, (245) 2 --> (3382) 94:PEGB0, ND11, *, NI0
			10'd45 : rdata = 48'b000111110000000001100001011100000000000000000000;
			// PEs: 2, 1 -> 1
			// srcs: (1756, 52)(3) 1, (3383) -141 --> (4167) -141:NM0, PENB, *, PEGB1
			10'd46 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 0, 2 -> 3
			// srcs: (1757, 36)(3140) 47, (247) 0 --> (3384) 0:PEGB0, ND3, *, PENB
			10'd47 : rdata = 48'b000111110000000001100000011000000000000100000000;
			// PEs: 2, 2 -> 
			// srcs: (1758, 51)(3) 1, (3382) 94 --> (4166) 94:NM0, NI0, *, 
			10'd48 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 2, 2 -> 2
			// srcs: (1761, 67)(1030) -3, (4166) 94 --> (4950) -97:NW11, ALU, -, NW11
			10'd49 : rdata = 48'b000100100000101100111111111000000110110000000000;
			// PEs: 2, 3 -> 2
			// srcs: (1766, 68)(1032) -1, (4168) 0 --> (4952) -1:NW3, PEGB3, -, NW3
			10'd50 : rdata = 48'b000100100000001111100000110000000100110000000000;
			// PEs: 2, 1 -> 1
			// srcs: (1836, 53)(3) 1, (3463) -94 --> (4247) -94:NM0, PENB, *, PEGB1
			10'd51 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 0, 2 -> 3
			// srcs: (1837, 37)(3140) 47, (327) 1 --> (3464) 47:PEGB0, ND4, *, PENB
			10'd52 : rdata = 48'b000111110000000001100000100000000000000100000000;
			// PEs: 2, 3 -> 2
			// srcs: (1846, 69)(1112) -3, (4248) 47 --> (5032) -50:NW4, PEGB3, -, NW4
			10'd53 : rdata = 48'b000100100000010011100000110000000101000000000000;
			// PEs: 2, 1 -> 1
			// srcs: (1916, 54)(3) 1, (3543) -94 --> (4327) -94:NM0, PENB, *, PEGB1
			10'd54 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 0, 2 -> 3
			// srcs: (1917, 38)(3140) 47, (407) 1 --> (3544) 47:PEGB0, ND5, *, PENB
			10'd55 : rdata = 48'b000111110000000001100000101000000000000100000000;
			// PEs: 2, 3 -> 2
			// srcs: (1926, 70)(1192) -3, (4328) 47 --> (5112) -50:NW5, PEGB3, -, NW5
			10'd56 : rdata = 48'b000100100000010111100000110000000101010000000000;
			// PEs: 2, 1 -> 1
			// srcs: (1936, 55)(3) 1, (3563) 94 --> (4347) 94:NM0, PENB, *, PEGB1
			10'd57 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 0, 2 -> 
			// srcs: (1939, 39)(3140) 47, (429) 0 --> (3566) 0:PEGB0, ND12, *, 
			10'd58 : rdata = 48'b000111110000000001100001100000000000000000000000;
			// PEs: 2, 2 -> 
			// srcs: (1942, 56)(3) 1, (3566) 0 --> (4350) 0:NM0, ALU, *, 
			10'd59 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 2, 2 -> 2
			// srcs: (1945, 71)(1214) 2, (4350) 0 --> (5134) 2:NW12, ALU, -, NW12
			10'd60 : rdata = 48'b000100100000110000111111111000000111000000000000;
			// PEs: 2, 1 -> 1
			// srcs: (1998, 57)(3) 1, (3625) -47 --> (4409) -47:NM0, PENB, *, PEGB1
			10'd61 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 0, 2 -> 3
			// srcs: (1999, 40)(3140) 47, (489) 1 --> (3626) 47:PEGB0, ND6, *, PENB
			10'd62 : rdata = 48'b000111110000000001100000110000000000000100000000;
			// PEs: 2, 3 -> 2
			// srcs: (2008, 72)(1274) 0, (4410) 47 --> (5194) -47:NW6, PEGB3, -, NW6
			10'd63 : rdata = 48'b000100100000011011100000110000000101100000000000;
			// PEs: 2, 1 -> 1
			// srcs: (2078, 58)(3) 1, (3705) 47 --> (4489) 47:NM0, PENB, *, PEGB1
			10'd64 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 0, 2 -> 3
			// srcs: (2079, 41)(3140) 47, (569) 0 --> (3706) 0:PEGB0, ND7, *, PENB
			10'd65 : rdata = 48'b000111110000000001100000111000000000000100000000;
			// PEs: 2, 3 -> 2
			// srcs: (2088, 73)(1354) -1, (4490) 0 --> (5274) -1:NW7, PEGB3, -, NW7
			10'd66 : rdata = 48'b000100100000011111100000110000000101110000000000;
			// PEs: 2, 1 -> 1
			// srcs: (2120, 59)(3) 1, (3747) -141 --> (4531) -141:NM0, PENB, *, PEGB1
			10'd67 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 0, 2 -> 
			// srcs: (2123, 42)(3140) 47, (613) -3 --> (3750) -141:PEGB0, ND13, *, 
			10'd68 : rdata = 48'b000111110000000001100001101000000000000000000000;
			// PEs: 2, 2 -> 
			// srcs: (2126, 60)(3) 1, (3750) -141 --> (4534) -141:NM0, ALU, *, 
			10'd69 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 2, 2 -> 2
			// srcs: (2129, 74)(1398) 1, (4534) -141 --> (5318) 142:NW13, ALU, -, NW13
			10'd70 : rdata = 48'b000100100000110100111111111000000111010000000000;
			// PEs: 2, 1 -> 1
			// srcs: (2158, 61)(3) 1, (3785) 94 --> (4569) 94:NM0, PENB, *, PEGB1
			10'd71 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 0, 2 -> 3
			// srcs: (2159, 43)(3140) 47, (649) -1 --> (3786) -47:PEGB0, ND8, *, PENB
			10'd72 : rdata = 48'b000111110000000001100001000000000000000100000000;
			// PEs: 2, 3 -> 2
			// srcs: (2168, 75)(1434) -1, (4570) -47 --> (5354) 46:NW8, PEGB3, -, NW8
			10'd73 : rdata = 48'b000100100000100011100000110000000110000000000000;
			// PEs: 2, 1 -> 1
			// srcs: (2240, 62)(3) 1, (3867) 47 --> (4651) 47:NM0, PENB, *, PEGB1
			10'd74 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 0, 2 -> 3
			// srcs: (2241, 44)(3140) 47, (731) 1 --> (3868) 47:PEGB0, ND9, *, PENB
			10'd75 : rdata = 48'b000111110000000001100001001000000000000100000000;
			// PEs: 2, 3 -> 2
			// srcs: (2250, 76)(1516) -3, (4652) 47 --> (5436) -50:NW9, PEGB3, -, NW9
			10'd76 : rdata = 48'b000100100000100111100000110000000110010000000000;
			default : rdata = 48'b000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 3) begin
	always @(*) begin
		case(address)
			// PEs: 3, 3 -> 3
			// srcs: (1, 0)(6) 0, (791) -2 --> (1575) 0:ND0, NW0, *, NI0
			10'd0 : rdata = 48'b000110110000000001000000000100000000000000000000;
			// PEs: 3, 3 -> 0
			// srcs: (2, 1)(87) 1, (872) 0 --> (1656) 0:ND1, NW1, *, PEGB0
			10'd1 : rdata = 48'b000110110000000101000000001000000000000010000000;
			// PEs: 3, 3 -> 0
			// srcs: (3, 2)(167) 1, (952) -2 --> (1736) -2:ND2, NW2, *, PEGB0
			10'd2 : rdata = 48'b000110110000001001000000010000000000000010000000;
			// PEs: 3, 3 -> 3
			// srcs: (4, 3)(249) 1, (1034) 2 --> (1818) 2:ND3, NW3, *, NI1
			10'd3 : rdata = 48'b000110110000001101000000011100001000000000000000;
			// PEs: 3, 3 -> 0
			// srcs: (5, 4)(329) 2, (1114) 2 --> (1898) 4:ND4, NW4, *, PEGB0
			10'd4 : rdata = 48'b000110110000010001000000100000000000000010000000;
			// PEs: 3, 3 -> 0
			// srcs: (6, 5)(409) 0, (1194) -2 --> (1978) 0:ND5, NW5, *, PEGB0
			10'd5 : rdata = 48'b000110110000010101000000101000000000000010000000;
			// PEs: 3, 3 -> 0
			// srcs: (7, 6)(491) -3, (1276) 2 --> (2060) -6:ND6, NW6, *, PEGB0
			10'd6 : rdata = 48'b000110110000011001000000110000000000000010000000;
			// PEs: 3, 3 -> 0
			// srcs: (8, 7)(571) -2, (1356) -1 --> (2140) 2:ND7, NW7, *, PEGB0
			10'd7 : rdata = 48'b000110110000011101000000111000000000000010000000;
			// PEs: 3, 3 -> 5
			// srcs: (9, 8)(651) 1, (1436) -3 --> (2220) -3:ND8, NW8, *, PEGB5
			10'd8 : rdata = 48'b000110110000100001000001000000000000000011010000;
			// PEs: 3, 3 -> 5
			// srcs: (10, 9)(733) 0, (1518) 0 --> (2302) 0:ND9, NW9, *, PEGB5
			10'd9 : rdata = 48'b000110110000100101000001001000000000000011010000;
			// PEs: 3, 3 -> 3
			// srcs: (11, 10)(68) 0, (853) 2 --> (1637) 0:ND10, NW10, *, NI2
			10'd10 : rdata = 48'b000110110000101001000001010100010000000000000000;
			// PEs: 3, 3 -> 3
			// srcs: (12, 11)(248) 1, (1033) -1 --> (1817) -1:ND11, NW11, *, NI3
			10'd11 : rdata = 48'b000110110000101101000001011100011000000000000000;
			// PEs: 3, 3 -> 3
			// srcs: (13, 12)(432) -2, (1217) 0 --> (2001) 0:ND12, NW12, *, NI4
			10'd12 : rdata = 48'b000110110000110001000001100100100000000000000000;
			// PEs: 3, 3 -> 3
			// srcs: (14, 13)(616) -2, (1401) 1 --> (2185) -2:ND13, NW13, *, NI5
			10'd13 : rdata = 48'b000110110000110101000001101100101000000000000000;
			// PEs: 0 -> 
			// srcs: (18, 14)(1584) -4 --> (1584) -4:PEGB0, pass, 
			10'd14 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 0, 3 -> 0
			// srcs: (27, 15)(1583) -4, (1584) -4 --> (2365) -8:PEGB0, ALU, +, PEGB0
			10'd15 : rdata = 48'b000011110000000000111111111000000000000010000000;
			// PEs: 0 -> 
			// srcs: (39, 16)(1728) 6 --> (1728) 6:PEGB0, pass, 
			10'd16 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 0, 3 -> 3
			// srcs: (48, 17)(1727) 0, (1728) 6 --> (2508) 6:PEGB0, ALU, +, NI6
			10'd17 : rdata = 48'b000011110000000000111111111100110000000000000000;
			// PEs: 0 -> 
			// srcs: (70, 18)(1893) 0 --> (1893) 0:PEGB0, pass, 
			10'd18 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 0, 3 -> 3
			// srcs: (79, 19)(1892) 2, (1893) 0 --> (2673) 2:PEGB0, ALU, +, NI7
			10'd19 : rdata = 48'b000011110000000000111111111100111000000000000000;
			// PEs: 3 -> 0
			// srcs: (107, 20)(1575) 0 --> (1575) 0:NI0, pass, PEGB0
			10'd20 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 3 -> 0
			// srcs: (108, 21)(1818) 2 --> (1818) 2:NI1, pass, PEGB0
			10'd21 : rdata = 48'b110001010000000100000000000000000000000010000000;
			// PEs: 3 -> 0
			// srcs: (113, 22)(1637) 0 --> (1637) 0:NI2, pass, PEGB0
			10'd22 : rdata = 48'b110001010000001000000000000000000000000010000000;
			// PEs: 3 -> 0
			// srcs: (131, 23)(2508) 6 --> (2508) 6:NI6, pass, PEGB0
			10'd23 : rdata = 48'b110001010000011000000000000000000000000010000000;
			// PEs: 3 -> 0
			// srcs: (157, 25)(2673) 2 --> (2673) 2:NI7, pass, PEGB0
			10'd24 : rdata = 48'b110001010000011100000000000000000000000010000000;
			// PEs: 3 -> 0
			// srcs: (166, 26)(2001) 0 --> (2001) 0:NI4, pass, PEGB0
			10'd25 : rdata = 48'b110001010000010000000000000000000000000010000000;
			// PEs: 3 -> 0
			// srcs: (183, 27)(2185) -2 --> (2185) -2:NI5, pass, PEGB0
			10'd26 : rdata = 48'b110001010000010100000000000000000000000010000000;
			// PEs: 3 -> 0
			// srcs: (195, 24)(1817) -1 --> (1817) -1:NI3, pass, PEGB0
			10'd27 : rdata = 48'b110001010000001100000000000000000000000010000000;
			// PEs: 1 -> 
			// srcs: (532, 28)(2588) 8 --> (2588) 8:PEGB1, pass, 
			10'd28 : rdata = 48'b110001110000001000000000000000000000000000000000;
			// PEs: 3, 5 -> 0
			// srcs: (535, 29)(2588) 8, (2590) 6 --> (2591) 14:ALU, PEGB5, +, PEGB0
			10'd29 : rdata = 48'b000010011111111111100001010000000000000010000000;
			// PEs: 0, 3 -> 4
			// srcs: (1517, 30)(3140) 47, (6) 0 --> (3143) 0:PEGB0, ND0, *, PENB
			10'd30 : rdata = 48'b000111110000000001100000000000000000000100000000;
			// PEs: 3, 2 -> 2
			// srcs: (1519, 44)(3) 1, (3142) -47 --> (3926) -47:NM0, PENB, *, PEGB2
			10'd31 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 3, 4 -> 3
			// srcs: (1526, 59)(791) -2, (3927) 0 --> (4711) -2:NW0, PEGB4, -, NW0
			10'd32 : rdata = 48'b000100100000000011100001000000000100000000000000;
			// PEs: 0, 3 -> 
			// srcs: (1578, 31)(3140) 47, (68) 0 --> (3205) 0:PEGB0, ND10, *, 
			10'd33 : rdata = 48'b000111110000000001100001010000000000000000000000;
			// PEs: 3, 3 -> 
			// srcs: (1581, 45)(3) 1, (3205) 0 --> (3989) 0:NM0, ALU, *, 
			10'd34 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 3, 3 -> 3
			// srcs: (1584, 60)(853) 2, (3989) 0 --> (4773) 2:NW10, ALU, -, NW10
			10'd35 : rdata = 48'b000100100000101000111111111000000110100000000000;
			// PEs: 0, 3 -> 4
			// srcs: (1597, 32)(3140) 47, (87) 1 --> (3224) 47:PEGB0, ND1, *, PENB
			10'd36 : rdata = 48'b000111110000000001100000001000000000000100000000;
			// PEs: 3, 2 -> 2
			// srcs: (1598, 46)(3) 1, (3222) 94 --> (4006) 94:NM0, PENB, *, PEGB2
			10'd37 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 3, 4 -> 3
			// srcs: (1606, 61)(872) 0, (4008) 47 --> (4792) -47:NW1, PEGB4, -, NW1
			10'd38 : rdata = 48'b000100100000000111100001000000000100010000000000;
			// PEs: 0, 3 -> 4
			// srcs: (1677, 33)(3140) 47, (167) 1 --> (3304) 47:PEGB0, ND2, *, PENB
			10'd39 : rdata = 48'b000111110000000001100000010000000000000100000000;
			// PEs: 3, 2 -> 2
			// srcs: (1678, 47)(3) 1, (3302) -47 --> (4086) -47:NM0, PENB, *, PEGB2
			10'd40 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 3, 4 -> 3
			// srcs: (1686, 62)(952) -2, (4088) 47 --> (4872) -49:NW2, PEGB4, -, NW2
			10'd41 : rdata = 48'b000100100000001011100001000000000100100000000000;
			// PEs: 0, 3 -> 4
			// srcs: (1758, 34)(3140) 47, (248) 1 --> (3385) 47:PEGB0, ND11, *, PENB
			10'd42 : rdata = 48'b000111110000000001100001011000000000000100000000;
			// PEs: 0, 3 -> 3
			// srcs: (1759, 35)(3140) 47, (249) 1 --> (3386) 47:PEGB0, ND3, *, NI0
			10'd43 : rdata = 48'b000111110000000001100000011100000000000000000000;
			// PEs: 3, 2 -> 2
			// srcs: (1760, 48)(3) 1, (3384) 0 --> (4168) 0:NM0, PENB, *, PEGB2
			10'd44 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 3, 3 -> 
			// srcs: (1762, 49)(3) 1, (3386) 47 --> (4170) 47:NM0, NI0, *, 
			10'd45 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 3, 3 -> 3
			// srcs: (1765, 64)(1034) 2, (4170) 47 --> (4954) -45:NW3, ALU, -, NW3
			10'd46 : rdata = 48'b000100100000001100111111111000000100110000000000;
			// PEs: 3, 4 -> 3
			// srcs: (1767, 63)(1033) -1, (4169) 47 --> (4953) -48:NW11, PEGB4, -, NW11
			10'd47 : rdata = 48'b000100100000101111100001000000000110110000000000;
			// PEs: 0, 3 -> 4
			// srcs: (1839, 36)(3140) 47, (329) 2 --> (3466) 94:PEGB0, ND4, *, PENB
			10'd48 : rdata = 48'b000111110000000001100000100000000000000100000000;
			// PEs: 3, 2 -> 2
			// srcs: (1840, 50)(3) 1, (3464) 47 --> (4248) 47:NM0, PENB, *, PEGB2
			10'd49 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 3, 4 -> 3
			// srcs: (1848, 65)(1114) 2, (4250) 94 --> (5034) -92:NW4, PEGB4, -, NW4
			10'd50 : rdata = 48'b000100100000010011100001000000000101000000000000;
			// PEs: 0, 3 -> 4
			// srcs: (1919, 37)(3140) 47, (409) 0 --> (3546) 0:PEGB0, ND5, *, PENB
			10'd51 : rdata = 48'b000111110000000001100000101000000000000100000000;
			// PEs: 3, 2 -> 2
			// srcs: (1920, 51)(3) 1, (3544) 47 --> (4328) 47:NM0, PENB, *, PEGB2
			10'd52 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 3, 4 -> 3
			// srcs: (1928, 66)(1194) -2, (4330) 0 --> (5114) -2:NW5, PEGB4, -, NW5
			10'd53 : rdata = 48'b000100100000010111100001000000000101010000000000;
			// PEs: 0, 3 -> 
			// srcs: (1942, 38)(3140) 47, (432) -2 --> (3569) -94:PEGB0, ND12, *, 
			10'd54 : rdata = 48'b000111110000000001100001100000000000000000000000;
			// PEs: 3, 3 -> 
			// srcs: (1945, 52)(3) 1, (3569) -94 --> (4353) -94:NM0, ALU, *, 
			10'd55 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 3, 3 -> 3
			// srcs: (1948, 67)(1217) 0, (4353) -94 --> (5137) 94:NW12, ALU, -, NW12
			10'd56 : rdata = 48'b000100100000110000111111111000000111000000000000;
			// PEs: 0, 3 -> 3
			// srcs: (2001, 39)(3140) 47, (491) -3 --> (3628) -141:PEGB0, ND6, *, NI0
			10'd57 : rdata = 48'b000111110000000001100000110100000000000000000000;
			// PEs: 3, 2 -> 2
			// srcs: (2002, 53)(3) 1, (3626) 47 --> (4410) 47:NM0, PENB, *, PEGB2
			10'd58 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 3, 3 -> 
			// srcs: (2004, 54)(3) 1, (3628) -141 --> (4412) -141:NM0, NI0, *, 
			10'd59 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 3, 3 -> 3
			// srcs: (2007, 68)(1276) 2, (4412) -141 --> (5196) 143:NW6, ALU, -, NW6
			10'd60 : rdata = 48'b000100100000011000111111111000000101100000000000;
			// PEs: 0, 3 -> 4
			// srcs: (2081, 40)(3140) 47, (571) -2 --> (3708) -94:PEGB0, ND7, *, PENB
			10'd61 : rdata = 48'b000111110000000001100000111000000000000100000000;
			// PEs: 3, 2 -> 2
			// srcs: (2082, 55)(3) 1, (3706) 0 --> (4490) 0:NM0, PENB, *, PEGB2
			10'd62 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 3, 4 -> 3
			// srcs: (2090, 69)(1356) -1, (4492) -94 --> (5276) 93:NW7, PEGB4, -, NW7
			10'd63 : rdata = 48'b000100100000011111100001000000000101110000000000;
			// PEs: 0, 3 -> 
			// srcs: (2126, 41)(3140) 47, (616) -2 --> (3753) -94:PEGB0, ND13, *, 
			10'd64 : rdata = 48'b000111110000000001100001101000000000000000000000;
			// PEs: 3, 3 -> 
			// srcs: (2129, 56)(3) 1, (3753) -94 --> (4537) -94:NM0, ALU, *, 
			10'd65 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 3, 3 -> 3
			// srcs: (2132, 70)(1401) 1, (4537) -94 --> (5321) 95:NW13, ALU, -, NW13
			10'd66 : rdata = 48'b000100100000110100111111111000000111010000000000;
			// PEs: 0, 3 -> 4
			// srcs: (2161, 42)(3140) 47, (651) 1 --> (3788) 47:PEGB0, ND8, *, PENB
			10'd67 : rdata = 48'b000111110000000001100001000000000000000100000000;
			// PEs: 3, 2 -> 2
			// srcs: (2162, 57)(3) 1, (3786) -47 --> (4570) -47:NM0, PENB, *, PEGB2
			10'd68 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 3, 4 -> 3
			// srcs: (2170, 71)(1436) -3, (4572) 47 --> (5356) -50:NW8, PEGB4, -, NW8
			10'd69 : rdata = 48'b000100100000100011100001000000000110000000000000;
			// PEs: 0, 3 -> 4
			// srcs: (2243, 43)(3140) 47, (733) 0 --> (3870) 0:PEGB0, ND9, *, PENB
			10'd70 : rdata = 48'b000111110000000001100001001000000000000100000000;
			// PEs: 3, 2 -> 2
			// srcs: (2244, 58)(3) 1, (3868) 47 --> (4652) 47:NM0, PENB, *, PEGB2
			10'd71 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 3, 4 -> 3
			// srcs: (2252, 72)(1518) 0, (4654) 0 --> (5438) 0:NW9, PEGB4, -, NW9
			10'd72 : rdata = 48'b000100100000100111100001000000000110010000000000;
			default : rdata = 48'b000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 4) begin
	always @(*) begin
		case(address)
			// PEs: 4, 4 -> 4
			// srcs: (1, 0)(7) 0, (792) 1 --> (1576) 0:ND0, NW0, *, NI0
			10'd0 : rdata = 48'b000110110000000001000000000100000000000000000000;
			// PEs: 4, 4 -> 0
			// srcs: (2, 1)(88) -1, (873) -1 --> (1657) 1:ND1, NW1, *, PEGB0
			10'd1 : rdata = 48'b000110110000000101000000001000000000000010000000;
			// PEs: 4, 4 -> 0
			// srcs: (3, 2)(168) 0, (953) -2 --> (1737) 0:ND2, NW2, *, PEGB0
			10'd2 : rdata = 48'b000110110000001001000000010000000000000010000000;
			// PEs: 4, 4 -> 4
			// srcs: (4, 3)(250) -3, (1035) -3 --> (1819) 9:ND3, NW3, *, NI1
			10'd3 : rdata = 48'b000110110000001101000000011100001000000000000000;
			// PEs: 4, 4 -> 0
			// srcs: (5, 4)(330) 1, (1115) 0 --> (1899) 0:ND4, NW4, *, PEGB0
			10'd4 : rdata = 48'b000110110000010001000000100000000000000010000000;
			// PEs: 4, 4 -> 0
			// srcs: (6, 5)(410) 1, (1195) 0 --> (1979) 0:ND5, NW5, *, PEGB0
			10'd5 : rdata = 48'b000110110000010101000000101000000000000010000000;
			// PEs: 4, 4 -> 0
			// srcs: (7, 6)(492) -1, (1277) 2 --> (2061) -2:ND6, NW6, *, PEGB0
			10'd6 : rdata = 48'b000110110000011001000000110000000000000010000000;
			// PEs: 4, 4 -> 0
			// srcs: (8, 7)(572) 2, (1357) -1 --> (2141) -2:ND7, NW7, *, PEGB0
			10'd7 : rdata = 48'b000110110000011101000000111000000000000010000000;
			// PEs: 4, 4 -> 5
			// srcs: (9, 8)(652) -3, (1437) -1 --> (2221) 3:ND8, NW8, *, PENB
			10'd8 : rdata = 48'b000110110000100001000001000000000000000100000000;
			// PEs: 4, 4 -> 5
			// srcs: (10, 9)(734) 0, (1519) 1 --> (2303) 0:ND9, NW9, *, PENB
			10'd9 : rdata = 48'b000110110000100101000001001000000000000100000000;
			// PEs: 4, 4 -> 4
			// srcs: (11, 10)(71) -1, (856) 1 --> (1640) -1:ND10, NW10, *, NI2
			10'd10 : rdata = 48'b000110110000101001000001010100010000000000000000;
			// PEs: 4, 4 -> 4
			// srcs: (12, 11)(255) -3, (1040) -1 --> (1824) 3:ND11, NW11, *, NI3
			10'd11 : rdata = 48'b000110110000101101000001011100011000000000000000;
			// PEs: 4, 4 -> 4
			// srcs: (13, 12)(435) -2, (1220) 1 --> (2004) -2:ND12, NW12, *, NI4
			10'd12 : rdata = 48'b000110110000110001000001100100100000000000000000;
			// PEs: 4, 4 -> 4
			// srcs: (14, 13)(619) 2, (1404) 0 --> (2188) 0:ND13, NW13, *, NI5
			10'd13 : rdata = 48'b000110110000110101000001101100101000000000000000;
			// PEs: 2 -> 
			// srcs: (15, 18)(2218) 1 --> (2218) 1:PEGB2, pass, 
			10'd14 : rdata = 48'b110001110000010000000000000000000000000000000000;
			// PEs: 1, 4 -> 4
			// srcs: (17, 19)(2217) 0, (2218) 1 --> (2997) 1:PEGB1, ALU, +, NI6
			10'd15 : rdata = 48'b000011110000001000111111111100110000000000000000;
			// PEs: 0 -> 
			// srcs: (20, 14)(1587) 3 --> (1587) 3:PEGB0, pass, 
			10'd16 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 0, 4 -> 0
			// srcs: (29, 15)(1586) -4, (1587) 3 --> (2369) -1:PEGB0, ALU, +, PEGB0
			10'd17 : rdata = 48'b000011110000000000111111111000000000000010000000;
			// PEs: 0 -> 
			// srcs: (41, 16)(1731) -2 --> (1731) -2:PEGB0, pass, 
			10'd18 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 0, 4 -> 4
			// srcs: (50, 17)(1730) 0, (1731) -2 --> (2510) -2:PEGB0, ALU, +, NI7
			10'd19 : rdata = 48'b000011110000000000111111111100111000000000000000;
			// PEs: 4 -> 0
			// srcs: (113, 22)(1640) -1 --> (1640) -1:NI2, pass, PEGB0
			10'd20 : rdata = 48'b110001010000001000000000000000000000000010000000;
			// PEs: 4 -> 0
			// srcs: (119, 20)(1576) 0 --> (1576) 0:NI0, pass, PEGB0
			10'd21 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 4 -> 0
			// srcs: (120, 21)(1819) 9 --> (1819) 9:NI1, pass, PEGB0
			10'd22 : rdata = 48'b110001010000000100000000000000000000000010000000;
			// PEs: 4 -> 0
			// srcs: (131, 23)(2510) -2 --> (2510) -2:NI7, pass, PEGB0
			10'd23 : rdata = 48'b110001010000011100000000000000000000000010000000;
			// PEs: 4 -> 0
			// srcs: (146, 24)(1824) 3 --> (1824) 3:NI3, pass, PEGB0
			10'd24 : rdata = 48'b110001010000001100000000000000000000000010000000;
			// PEs: 4 -> 0
			// srcs: (192, 26)(2188) 0 --> (2188) 0:NI5, pass, PEGB0
			10'd25 : rdata = 48'b110001010000010100000000000000000000000010000000;
			// PEs: 4 -> 0
			// srcs: (220, 25)(2004) -2 --> (2004) -2:NI4, pass, PEGB0
			10'd26 : rdata = 48'b110001010000010000000000000000000000000010000000;
			// PEs: 4 -> 0
			// srcs: (253, 27)(2997) 1 --> (2997) 1:NI6, pass, PEGB0
			10'd27 : rdata = 48'b110001010000011000000000000000000000000010000000;
			// PEs: 0 -> 
			// srcs: (996, 28)(3095) -3 --> (3095) -3:PEGB0, pass, 
			10'd28 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 4, 1 -> 0
			// srcs: (998, 29)(3095) -3, (3097) 2 --> (3098) -1:ALU, PEGB1, +, PEGB0
			10'd29 : rdata = 48'b000010011111111111100000010000000000000010000000;
			// PEs: 0, 4 -> 5
			// srcs: (1518, 30)(3140) 47, (7) 0 --> (3144) 0:PEGB0, ND0, *, PENB
			10'd30 : rdata = 48'b000111110000000001100000000000000000000100000000;
			// PEs: 4, 3 -> 3
			// srcs: (1520, 44)(3) 1, (3143) 0 --> (3927) 0:NM0, PENB, *, PEGB3
			10'd31 : rdata = 48'b000111000000000011011111110000000000000010110000;
			// PEs: 4, 5 -> 4
			// srcs: (1527, 59)(792) 1, (3928) 0 --> (4712) 1:NW0, PEGB5, -, NW0
			10'd32 : rdata = 48'b000100100000000011100001010000000100000000000000;
			// PEs: 0, 4 -> 
			// srcs: (1581, 31)(3140) 47, (71) -1 --> (3208) -47:PEGB0, ND10, *, 
			10'd33 : rdata = 48'b000111110000000001100001010000000000000000000000;
			// PEs: 4, 4 -> 
			// srcs: (1584, 45)(3) 1, (3208) -47 --> (3992) -47:NM0, ALU, *, 
			10'd34 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 4, 4 -> 4
			// srcs: (1587, 60)(856) 1, (3992) -47 --> (4776) 48:NW10, ALU, -, NW10
			10'd35 : rdata = 48'b000100100000101000111111111000000110100000000000;
			// PEs: 0, 4 -> 5
			// srcs: (1598, 32)(3140) 47, (88) -1 --> (3225) -47:PEGB0, ND1, *, PENB
			10'd36 : rdata = 48'b000111110000000001100000001000000000000100000000;
			// PEs: 4, 3 -> 3
			// srcs: (1600, 46)(3) 1, (3224) 47 --> (4008) 47:NM0, PENB, *, PEGB3
			10'd37 : rdata = 48'b000111000000000011011111110000000000000010110000;
			// PEs: 4, 5 -> 4
			// srcs: (1607, 61)(873) -1, (4009) -47 --> (4793) 46:NW1, PEGB5, -, NW1
			10'd38 : rdata = 48'b000100100000000111100001010000000100010000000000;
			// PEs: 0, 4 -> 5
			// srcs: (1678, 33)(3140) 47, (168) 0 --> (3305) 0:PEGB0, ND2, *, PENB
			10'd39 : rdata = 48'b000111110000000001100000010000000000000100000000;
			// PEs: 4, 3 -> 3
			// srcs: (1680, 47)(3) 1, (3304) 47 --> (4088) 47:NM0, PENB, *, PEGB3
			10'd40 : rdata = 48'b000111000000000011011111110000000000000010110000;
			// PEs: 4, 5 -> 4
			// srcs: (1687, 62)(953) -2, (4089) 0 --> (4873) -2:NW2, PEGB5, -, NW2
			10'd41 : rdata = 48'b000100100000001011100001010000000100100000000000;
			// PEs: 0, 4 -> 5
			// srcs: (1760, 34)(3140) 47, (250) -3 --> (3387) -141:PEGB0, ND3, *, PENB
			10'd42 : rdata = 48'b000111110000000001100000011000000000000100000000;
			// PEs: 4, 3 -> 3
			// srcs: (1761, 48)(3) 1, (3385) 47 --> (4169) 47:NM0, PENB, *, PEGB3
			10'd43 : rdata = 48'b000111000000000011011111110000000000000010110000;
			// PEs: 0, 4 -> 
			// srcs: (1765, 35)(3140) 47, (255) -3 --> (3392) -141:PEGB0, ND11, *, 
			10'd44 : rdata = 48'b000111110000000001100001011000000000000000000000;
			// PEs: 4, 4 -> 4
			// srcs: (1768, 49)(3) 1, (3392) -141 --> (4176) -141:NM0, ALU, *, NI0
			10'd45 : rdata = 48'b000111000000000000111111111100000000000000000000;
			// PEs: 4, 5 -> 4
			// srcs: (1769, 63)(1035) -3, (4171) -141 --> (4955) 138:NW3, PEGB5, -, NW3
			10'd46 : rdata = 48'b000100100000001111100001010000000100110000000000;
			// PEs: 4, 4 -> 4
			// srcs: (1771, 64)(1040) -1, (4176) -141 --> (4960) 140:NW11, NI0, -, NW11
			10'd47 : rdata = 48'b000100100000101110100000000000000110110000000000;
			// PEs: 0, 4 -> 5
			// srcs: (1840, 36)(3140) 47, (330) 1 --> (3467) 47:PEGB0, ND4, *, PENB
			10'd48 : rdata = 48'b000111110000000001100000100000000000000100000000;
			// PEs: 4, 3 -> 3
			// srcs: (1842, 50)(3) 1, (3466) 94 --> (4250) 94:NM0, PENB, *, PEGB3
			10'd49 : rdata = 48'b000111000000000011011111110000000000000010110000;
			// PEs: 4, 5 -> 4
			// srcs: (1849, 65)(1115) 0, (4251) 47 --> (5035) -47:NW4, PEGB5, -, NW4
			10'd50 : rdata = 48'b000100100000010011100001010000000101000000000000;
			// PEs: 0, 4 -> 4
			// srcs: (1920, 37)(3140) 47, (410) 1 --> (3547) 47:PEGB0, ND5, *, NI0
			10'd51 : rdata = 48'b000111110000000001100000101100000000000000000000;
			// PEs: 4, 3 -> 3
			// srcs: (1922, 51)(3) 1, (3546) 0 --> (4330) 0:NM0, PENB, *, PEGB3
			10'd52 : rdata = 48'b000111000000000011011111110000000000000010110000;
			// PEs: 4, 4 -> 
			// srcs: (1923, 52)(3) 1, (3547) 47 --> (4331) 47:NM0, NI0, *, 
			10'd53 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 4, 4 -> 4
			// srcs: (1926, 66)(1195) 0, (4331) 47 --> (5115) -47:NW5, ALU, -, NW5
			10'd54 : rdata = 48'b000100100000010100111111111000000101010000000000;
			// PEs: 0, 4 -> 
			// srcs: (1945, 38)(3140) 47, (435) -2 --> (3572) -94:PEGB0, ND12, *, 
			10'd55 : rdata = 48'b000111110000000001100001100000000000000000000000;
			// PEs: 4, 4 -> 
			// srcs: (1948, 53)(3) 1, (3572) -94 --> (4356) -94:NM0, ALU, *, 
			10'd56 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 4, 4 -> 4
			// srcs: (1951, 67)(1220) 1, (4356) -94 --> (5140) 95:NW12, ALU, -, NW12
			10'd57 : rdata = 48'b000100100000110000111111111000000111000000000000;
			// PEs: 0, 4 -> 
			// srcs: (2002, 39)(3140) 47, (492) -1 --> (3629) -47:PEGB0, ND6, *, 
			10'd58 : rdata = 48'b000111110000000001100000110000000000000000000000;
			// PEs: 4, 4 -> 
			// srcs: (2005, 54)(3) 1, (3629) -47 --> (4413) -47:NM0, ALU, *, 
			10'd59 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 4, 4 -> 4
			// srcs: (2008, 68)(1277) 2, (4413) -47 --> (5197) 49:NW6, ALU, -, NW6
			10'd60 : rdata = 48'b000100100000011000111111111000000101100000000000;
			// PEs: 0, 4 -> 5
			// srcs: (2082, 40)(3140) 47, (572) 2 --> (3709) 94:PEGB0, ND7, *, PENB
			10'd61 : rdata = 48'b000111110000000001100000111000000000000100000000;
			// PEs: 4, 3 -> 3
			// srcs: (2084, 55)(3) 1, (3708) -94 --> (4492) -94:NM0, PENB, *, PEGB3
			10'd62 : rdata = 48'b000111000000000011011111110000000000000010110000;
			// PEs: 4, 5 -> 4
			// srcs: (2091, 69)(1357) -1, (4493) 94 --> (5277) -95:NW7, PEGB5, -, NW7
			10'd63 : rdata = 48'b000100100000011111100001010000000101110000000000;
			// PEs: 0, 4 -> 
			// srcs: (2129, 41)(3140) 47, (619) 2 --> (3756) 94:PEGB0, ND13, *, 
			10'd64 : rdata = 48'b000111110000000001100001101000000000000000000000;
			// PEs: 4, 4 -> 
			// srcs: (2132, 56)(3) 1, (3756) 94 --> (4540) 94:NM0, ALU, *, 
			10'd65 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 4, 4 -> 4
			// srcs: (2135, 70)(1404) 0, (4540) 94 --> (5324) -94:NW13, ALU, -, NW13
			10'd66 : rdata = 48'b000100100000110100111111111000000111010000000000;
			// PEs: 0, 4 -> 5
			// srcs: (2162, 42)(3140) 47, (652) -3 --> (3789) -141:PEGB0, ND8, *, PENB
			10'd67 : rdata = 48'b000111110000000001100001000000000000000100000000;
			// PEs: 4, 3 -> 3
			// srcs: (2164, 57)(3) 1, (3788) 47 --> (4572) 47:NM0, PENB, *, PEGB3
			10'd68 : rdata = 48'b000111000000000011011111110000000000000010110000;
			// PEs: 4, 5 -> 4
			// srcs: (2171, 71)(1437) -1, (4573) -141 --> (5357) 140:NW8, PEGB5, -, NW8
			10'd69 : rdata = 48'b000100100000100011100001010000000110000000000000;
			// PEs: 0, 4 -> 5
			// srcs: (2244, 43)(3140) 47, (734) 0 --> (3871) 0:PEGB0, ND9, *, PENB
			10'd70 : rdata = 48'b000111110000000001100001001000000000000100000000;
			// PEs: 4, 3 -> 3
			// srcs: (2246, 58)(3) 1, (3870) 0 --> (4654) 0:NM0, PENB, *, PEGB3
			10'd71 : rdata = 48'b000111000000000011011111110000000000000010110000;
			// PEs: 4, 5 -> 4
			// srcs: (2253, 72)(1519) 1, (4655) 0 --> (5439) 1:NW9, PEGB5, -, NW9
			10'd72 : rdata = 48'b000100100000100111100001010000000110010000000000;
			default : rdata = 48'b000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 5) begin
	always @(*) begin
		case(address)
			// PEs: 5, 5 -> 0
			// srcs: (1, 0)(8) 2, (793) -2 --> (1577) -4:ND0, NW0, *, PEGB0
			10'd0 : rdata = 48'b000110110000000001000000000000000000000010000000;
			// PEs: 5, 5 -> 0
			// srcs: (2, 1)(90) -2, (875) -1 --> (1659) 2:ND1, NW1, *, PEGB0
			10'd1 : rdata = 48'b000110110000000101000000001000000000000010000000;
			// PEs: 5, 5 -> 0
			// srcs: (3, 2)(170) -1, (955) 1 --> (1739) -1:ND2, NW2, *, PEGB0
			10'd2 : rdata = 48'b000110110000001001000000010000000000000010000000;
			// PEs: 5, 5 -> 5
			// srcs: (4, 3)(251) 1, (1036) 2 --> (1820) 2:ND3, NW3, *, NI0
			10'd3 : rdata = 48'b000110110000001101000000011100000000000000000000;
			// PEs: 5, 5 -> 0
			// srcs: (5, 4)(332) 2, (1117) -1 --> (1901) -2:ND4, NW4, *, PEGB0
			10'd4 : rdata = 48'b000110110000010001000000100000000000000010000000;
			// PEs: 5, 5 -> 0
			// srcs: (6, 5)(412) -3, (1197) 2 --> (1981) -6:ND5, NW5, *, PEGB0
			10'd5 : rdata = 48'b000110110000010101000000101000000000000010000000;
			// PEs: 5, 5 -> 5
			// srcs: (7, 6)(494) 0, (1279) 2 --> (2063) 0:ND6, NW6, *, NI1
			10'd6 : rdata = 48'b000110110000011001000000110100001000000000000000;
			// PEs: 5, 5 -> 0
			// srcs: (8, 7)(574) -2, (1359) 0 --> (2143) 0:ND7, NW7, *, PEGB0
			10'd7 : rdata = 48'b000110110000011101000000111000000000000010000000;
			// PEs: 5, 5 -> 7
			// srcs: (9, 8)(654) 1, (1439) 0 --> (2223) 0:ND8, NW8, *, PEGB7
			10'd8 : rdata = 48'b000110110000100001000001000000000000000011110000;
			// PEs: 5, 5 -> 7
			// srcs: (10, 9)(736) 2, (1521) 0 --> (2305) 0:ND9, NW9, *, PEGB7
			10'd9 : rdata = 48'b000110110000100101000001001000000000000011110000;
			// PEs: 5, 5 -> 1
			// srcs: (11, 10)(74) -2, (859) -1 --> (1643) 2:ND10, NW10, *, PEGB1
			10'd10 : rdata = 48'b000110110000101001000001010000000000000010010000;
			// PEs: 5, 5 -> 5
			// srcs: (12, 11)(258) -3, (1043) -1 --> (1827) 3:ND11, NW11, *, NI2
			10'd11 : rdata = 48'b000110110000101101000001011100010000000000000000;
			// PEs: 5, 5 -> 5
			// srcs: (13, 12)(438) 0, (1223) 2 --> (2007) 0:ND12, NW12, *, NI3
			10'd12 : rdata = 48'b000110110000110001000001100100011000000000000000;
			// PEs: 5, 5 -> 5
			// srcs: (14, 13)(622) -2, (1407) -3 --> (2191) 6:ND13, NW13, *, NI4
			10'd13 : rdata = 48'b000110110000110101000001101100100000000000000000;
			// PEs: 3, 4 -> 5
			// srcs: (15, 18)(2220) -3, (2221) 3 --> (2999) 0:PEGB3, PENB, +, NI5
			10'd14 : rdata = 48'b000011110000011011011111110100101000000000000000;
			// PEs: 3, 4 -> 5
			// srcs: (16, 19)(2302) 0, (2303) 0 --> (3080) 0:PEGB3, PENB, +, NI6
			10'd15 : rdata = 48'b000011110000011011011111110100110000000000000000;
			// PEs: 0 -> 
			// srcs: (22, 14)(1590) 3 --> (1590) 3:PEGB0, pass, 
			10'd16 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 0, 5 -> 0
			// srcs: (31, 15)(1589) 6, (1590) 3 --> (2371) 9:PEGB0, ALU, +, PEGB0
			10'd17 : rdata = 48'b000011110000000000111111111000000000000010000000;
			// PEs: 0 -> 
			// srcs: (54, 16)(1804) -4 --> (1804) -4:PEGB0, pass, 
			10'd18 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 0, 5 -> 1
			// srcs: (64, 17)(1803) 0, (1804) -4 --> (2583) -4:PEGB0, ALU, +, PEGB1
			10'd19 : rdata = 48'b000011110000000000111111111000000000000010010000;
			// PEs: 7 -> 
			// srcs: (73, 22)(2589) 6 --> (2589) 6:PEGB7, pass, 
			10'd20 : rdata = 48'b110001110000111000000000000000000000000000000000;
			// PEs: 5, 1 -> 3
			// srcs: (76, 23)(2589) 6, (1811) 0 --> (2590) 6:ALU, PEGB1, +, PEGB3
			10'd21 : rdata = 48'b000010011111111111100000010000000000000010110000;
			// PEs: 5 -> 0
			// srcs: (129, 20)(1820) 2 --> (1820) 2:NI0, pass, PEGB0
			10'd22 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 5 -> 0
			// srcs: (145, 21)(2063) 0 --> (2063) 0:NI1, pass, PEGB0
			10'd23 : rdata = 48'b110001010000000100000000000000000000000010000000;
			// PEs: 5 -> 0
			// srcs: (146, 24)(1827) 3 --> (1827) 3:NI2, pass, PEGB0
			10'd24 : rdata = 48'b110001010000001000000000000000000000000010000000;
			// PEs: 5 -> 0
			// srcs: (158, 25)(2007) 0 --> (2007) 0:NI3, pass, PEGB0
			10'd25 : rdata = 48'b110001010000001100000000000000000000000010000000;
			// PEs: 5 -> 0
			// srcs: (171, 28)(3080) 0 --> (3080) 0:NI6, pass, PEGB0
			10'd26 : rdata = 48'b110001010000011000000000000000000000000010000000;
			// PEs: 5 -> 0
			// srcs: (192, 26)(2191) 6 --> (2191) 6:NI4, pass, PEGB0
			10'd27 : rdata = 48'b110001010000010000000000000000000000000010000000;
			// PEs: 5 -> 0
			// srcs: (261, 27)(2999) 0 --> (2999) 0:NI5, pass, PEGB0
			10'd28 : rdata = 48'b110001010000010100000000000000000000000010000000;
			// PEs: 0, 5 -> 6
			// srcs: (1519, 29)(3140) 47, (8) 2 --> (3145) 94:PEGB0, ND0, *, PENB
			10'd29 : rdata = 48'b000111110000000001100000000000000000000100000000;
			// PEs: 5, 4 -> 4
			// srcs: (1521, 43)(3) 1, (3144) 0 --> (3928) 0:NM0, PENB, *, PEGB4
			10'd30 : rdata = 48'b000111000000000011011111110000000000000011000000;
			// PEs: 5, 6 -> 5
			// srcs: (1528, 60)(793) -2, (3929) 94 --> (4713) -96:NW0, PEGB6, -, NW0
			10'd31 : rdata = 48'b000100100000000011100001100000000100000000000000;
			// PEs: 0, 5 -> 
			// srcs: (1584, 30)(3140) 47, (74) -2 --> (3211) -94:PEGB0, ND10, *, 
			10'd32 : rdata = 48'b000111110000000001100001010000000000000000000000;
			// PEs: 5, 5 -> 
			// srcs: (1587, 44)(3) 1, (3211) -94 --> (3995) -94:NM0, ALU, *, 
			10'd33 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 5, 5 -> 5
			// srcs: (1590, 61)(859) -1, (3995) -94 --> (4779) 93:NW10, ALU, -, NW10
			10'd34 : rdata = 48'b000100100000101000111111111000000110100000000000;
			// PEs: 0, 5 -> 5
			// srcs: (1600, 31)(3140) 47, (90) -2 --> (3227) -94:PEGB0, ND1, *, NI0
			10'd35 : rdata = 48'b000111110000000001100000001100000000000000000000;
			// PEs: 5, 4 -> 4
			// srcs: (1601, 45)(3) 1, (3225) -47 --> (4009) -47:NM0, PENB, *, PEGB4
			10'd36 : rdata = 48'b000111000000000011011111110000000000000011000000;
			// PEs: 5, 5 -> 
			// srcs: (1603, 46)(3) 1, (3227) -94 --> (4011) -94:NM0, NI0, *, 
			10'd37 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 5, 5 -> 5
			// srcs: (1606, 62)(875) -1, (4011) -94 --> (4795) 93:NW1, ALU, -, NW1
			10'd38 : rdata = 48'b000100100000000100111111111000000100010000000000;
			// PEs: 0, 5 -> 6
			// srcs: (1680, 32)(3140) 47, (170) -1 --> (3307) -47:PEGB0, ND2, *, PENB
			10'd39 : rdata = 48'b000111110000000001100000010000000000000100000000;
			// PEs: 5, 4 -> 4
			// srcs: (1681, 47)(3) 1, (3305) 0 --> (4089) 0:NM0, PENB, *, PEGB4
			10'd40 : rdata = 48'b000111000000000011011111110000000000000011000000;
			// PEs: 5, 6 -> 5
			// srcs: (1689, 63)(955) 1, (4091) -47 --> (4875) 48:NW2, PEGB6, -, NW2
			10'd41 : rdata = 48'b000100100000001011100001100000000100100000000000;
			// PEs: 0, 5 -> 6
			// srcs: (1761, 33)(3140) 47, (251) 1 --> (3388) 47:PEGB0, ND3, *, PENB
			10'd42 : rdata = 48'b000111110000000001100000011000000000000100000000;
			// PEs: 5, 4 -> 4
			// srcs: (1763, 48)(3) 1, (3387) -141 --> (4171) -141:NM0, PENB, *, PEGB4
			10'd43 : rdata = 48'b000111000000000011011111110000000000000011000000;
			// PEs: 0, 5 -> 5
			// srcs: (1768, 34)(3140) 47, (258) -3 --> (3395) -141:PEGB0, ND11, *, NI0
			10'd44 : rdata = 48'b000111110000000001100001011100000000000000000000;
			// PEs: 5, 6 -> 5
			// srcs: (1770, 64)(1036) 2, (4172) 47 --> (4956) -45:NW3, PEGB6, -, NW3
			10'd45 : rdata = 48'b000100100000001111100001100000000100110000000000;
			// PEs: 5, 5 -> 
			// srcs: (1771, 49)(3) 1, (3395) -141 --> (4179) -141:NM0, NI0, *, 
			10'd46 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 5, 5 -> 5
			// srcs: (1774, 65)(1043) -1, (4179) -141 --> (4963) 140:NW11, ALU, -, NW11
			10'd47 : rdata = 48'b000100100000101100111111111000000110110000000000;
			// PEs: 0, 5 -> 5
			// srcs: (1842, 35)(3140) 47, (332) 2 --> (3469) 94:PEGB0, ND4, *, NI0
			10'd48 : rdata = 48'b000111110000000001100000100100000000000000000000;
			// PEs: 5, 4 -> 4
			// srcs: (1843, 50)(3) 1, (3467) 47 --> (4251) 47:NM0, PENB, *, PEGB4
			10'd49 : rdata = 48'b000111000000000011011111110000000000000011000000;
			// PEs: 5, 5 -> 
			// srcs: (1845, 51)(3) 1, (3469) 94 --> (4253) 94:NM0, NI0, *, 
			10'd50 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 5, 5 -> 5
			// srcs: (1848, 66)(1117) -1, (4253) 94 --> (5037) -95:NW4, ALU, -, NW4
			10'd51 : rdata = 48'b000100100000010000111111111000000101000000000000;
			// PEs: 0, 5 -> 
			// srcs: (1922, 36)(3140) 47, (412) -3 --> (3549) -141:PEGB0, ND5, *, 
			10'd52 : rdata = 48'b000111110000000001100000101000000000000000000000;
			// PEs: 5, 5 -> 
			// srcs: (1925, 52)(3) 1, (3549) -141 --> (4333) -141:NM0, ALU, *, 
			10'd53 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 5, 5 -> 5
			// srcs: (1928, 67)(1197) 2, (4333) -141 --> (5117) 143:NW5, ALU, -, NW5
			10'd54 : rdata = 48'b000100100000010100111111111000000101010000000000;
			// PEs: 0, 5 -> 
			// srcs: (1948, 37)(3140) 47, (438) 0 --> (3575) 0:PEGB0, ND12, *, 
			10'd55 : rdata = 48'b000111110000000001100001100000000000000000000000;
			// PEs: 5, 5 -> 
			// srcs: (1951, 53)(3) 1, (3575) 0 --> (4359) 0:NM0, ALU, *, 
			10'd56 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 5, 5 -> 5
			// srcs: (1954, 68)(1223) 2, (4359) 0 --> (5143) 2:NW12, ALU, -, NW12
			10'd57 : rdata = 48'b000100100000110000111111111000000111000000000000;
			// PEs: 0, 5 -> 
			// srcs: (2004, 38)(3140) 47, (494) 0 --> (3631) 0:PEGB0, ND6, *, 
			10'd58 : rdata = 48'b000111110000000001100000110000000000000000000000;
			// PEs: 5, 5 -> 
			// srcs: (2007, 54)(3) 1, (3631) 0 --> (4415) 0:NM0, ALU, *, 
			10'd59 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 5, 5 -> 5
			// srcs: (2010, 69)(1279) 2, (4415) 0 --> (5199) 2:NW6, ALU, -, NW6
			10'd60 : rdata = 48'b000100100000011000111111111000000101100000000000;
			// PEs: 0, 5 -> 6
			// srcs: (2084, 39)(3140) 47, (574) -2 --> (3711) -94:PEGB0, ND7, *, PENB
			10'd61 : rdata = 48'b000111110000000001100000111000000000000100000000;
			// PEs: 5, 4 -> 4
			// srcs: (2085, 55)(3) 1, (3709) 94 --> (4493) 94:NM0, PENB, *, PEGB4
			10'd62 : rdata = 48'b000111000000000011011111110000000000000011000000;
			// PEs: 5, 6 -> 5
			// srcs: (2093, 70)(1359) 0, (4495) -94 --> (5279) 94:NW7, PEGB6, -, NW7
			10'd63 : rdata = 48'b000100100000011111100001100000000101110000000000;
			// PEs: 0, 5 -> 
			// srcs: (2132, 40)(3140) 47, (622) -2 --> (3759) -94:PEGB0, ND13, *, 
			10'd64 : rdata = 48'b000111110000000001100001101000000000000000000000;
			// PEs: 5, 5 -> 
			// srcs: (2135, 56)(3) 1, (3759) -94 --> (4543) -94:NM0, ALU, *, 
			10'd65 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 5, 5 -> 5
			// srcs: (2138, 71)(1407) -3, (4543) -94 --> (5327) 91:NW13, ALU, -, NW13
			10'd66 : rdata = 48'b000100100000110100111111111000000111010000000000;
			// PEs: 0, 5 -> 6
			// srcs: (2164, 41)(3140) 47, (654) 1 --> (3791) 47:PEGB0, ND8, *, PENB
			10'd67 : rdata = 48'b000111110000000001100001000000000000000100000000;
			// PEs: 5, 4 -> 4
			// srcs: (2165, 57)(3) 1, (3789) -141 --> (4573) -141:NM0, PENB, *, PEGB4
			10'd68 : rdata = 48'b000111000000000011011111110000000000000011000000;
			// PEs: 5, 6 -> 5
			// srcs: (2173, 72)(1439) 0, (4575) 47 --> (5359) -47:NW8, PEGB6, -, NW8
			10'd69 : rdata = 48'b000100100000100011100001100000000110000000000000;
			// PEs: 0, 5 -> 5
			// srcs: (2246, 42)(3140) 47, (736) 2 --> (3873) 94:PEGB0, ND9, *, NI0
			10'd70 : rdata = 48'b000111110000000001100001001100000000000000000000;
			// PEs: 5, 4 -> 4
			// srcs: (2247, 58)(3) 1, (3871) 0 --> (4655) 0:NM0, PENB, *, PEGB4
			10'd71 : rdata = 48'b000111000000000011011111110000000000000011000000;
			// PEs: 5, 5 -> 
			// srcs: (2249, 59)(3) 1, (3873) 94 --> (4657) 94:NM0, NI0, *, 
			10'd72 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 5, 5 -> 5
			// srcs: (2252, 73)(1521) 0, (4657) 94 --> (5441) -94:NW9, ALU, -, NW9
			10'd73 : rdata = 48'b000100100000100100111111111000000110010000000000;
			default : rdata = 48'b000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 6) begin
	always @(*) begin
		case(address)
			// PEs: 6, 6 -> 0
			// srcs: (1, 0)(9) 2, (794) -3 --> (1578) -6:ND0, NW0, *, PEGB0
			10'd0 : rdata = 48'b000110110000000001000000000000000000000010000000;
			// PEs: 6, 6 -> 0
			// srcs: (2, 1)(91) 0, (876) -1 --> (1660) 0:ND1, NW1, *, PEGB0
			10'd1 : rdata = 48'b000110110000000101000000001000000000000010000000;
			// PEs: 6, 6 -> 0
			// srcs: (3, 2)(171) 0, (956) 1 --> (1740) 0:ND2, NW2, *, PEGB0
			10'd2 : rdata = 48'b000110110000001001000000010000000000000010000000;
			// PEs: 6, 6 -> 6
			// srcs: (4, 3)(252) 0, (1037) 2 --> (1821) 0:ND3, NW3, *, NI0
			10'd3 : rdata = 48'b000110110000001101000000011100000000000000000000;
			// PEs: 6, 6 -> 0
			// srcs: (5, 4)(333) 2, (1118) -3 --> (1902) -6:ND4, NW4, *, PEGB0
			10'd4 : rdata = 48'b000110110000010001000000100000000000000010000000;
			// PEs: 6, 6 -> 0
			// srcs: (6, 5)(413) -1, (1198) 0 --> (1982) 0:ND5, NW5, *, PEGB0
			10'd5 : rdata = 48'b000110110000010101000000101000000000000010000000;
			// PEs: 6, 6 -> 6
			// srcs: (7, 6)(495) -3, (1280) 1 --> (2064) -3:ND6, NW6, *, NI1
			10'd6 : rdata = 48'b000110110000011001000000110100001000000000000000;
			// PEs: 6, 6 -> 0
			// srcs: (8, 7)(575) 2, (1360) 0 --> (2144) 0:ND7, NW7, *, PEGB0
			10'd7 : rdata = 48'b000110110000011101000000111000000000000010000000;
			// PEs: 6, 6 -> 7
			// srcs: (9, 8)(655) 1, (1440) 0 --> (2224) 0:ND8, NW8, *, PENB
			10'd8 : rdata = 48'b000110110000100001000001000000000000000100000000;
			// PEs: 6, 6 -> 7
			// srcs: (10, 9)(737) -2, (1522) 2 --> (2306) -4:ND9, NW9, *, PENB
			10'd9 : rdata = 48'b000110110000100101000001001000000000000100000000;
			// PEs: 6, 6 -> 0
			// srcs: (11, 10)(77) 0, (862) -3 --> (1646) 0:ND10, NW10, *, PEGB0
			10'd10 : rdata = 48'b000110110000101001000001010000000000000010000000;
			// PEs: 6, 6 -> 6
			// srcs: (12, 11)(261) -1, (1046) 0 --> (1830) 0:ND11, NW11, *, NI2
			10'd11 : rdata = 48'b000110110000101101000001011100010000000000000000;
			// PEs: 6, 6 -> 6
			// srcs: (13, 12)(441) 2, (1226) -1 --> (2010) -2:ND12, NW12, *, NI3
			10'd12 : rdata = 48'b000110110000110001000001100100011000000000000000;
			// PEs: 6, 6 -> 6
			// srcs: (14, 13)(625) -1, (1410) 1 --> (2194) -1:ND13, NW13, *, NI4
			10'd13 : rdata = 48'b000110110000110101000001101100100000000000000000;
			// PEs: 2 -> 
			// srcs: (15, 18)(2300) -3 --> (2300) -3:PEGB2, pass, 
			10'd14 : rdata = 48'b110001110000010000000000000000000000000000000000;
			// PEs: 1, 6 -> 6
			// srcs: (18, 19)(2299) 1, (2300) -3 --> (3077) -2:PEGB1, ALU, +, NI5
			10'd15 : rdata = 48'b000011110000001000111111111100101000000000000000;
			// PEs: 0 -> 
			// srcs: (24, 14)(1593) -3 --> (1593) -3:PEGB0, pass, 
			10'd16 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 0, 6 -> 0
			// srcs: (33, 15)(1592) 9, (1593) -3 --> (2374) 6:PEGB0, ALU, +, PEGB0
			10'd17 : rdata = 48'b000011110000000000111111111000000000000010000000;
			// PEs: 0 -> 
			// srcs: (56, 16)(1807) 4 --> (1807) 4:PEGB0, pass, 
			10'd18 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 0, 6 -> 1
			// srcs: (65, 17)(1806) 4, (1807) 4 --> (2587) 8:PEGB0, ALU, +, PEGB1
			10'd19 : rdata = 48'b000011110000000000111111111000000000000010010000;
			// PEs: 6 -> 0
			// srcs: (137, 20)(1821) 0 --> (1821) 0:NI0, pass, PEGB0
			10'd20 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 6 -> 0
			// srcs: (138, 22)(1830) 0 --> (1830) 0:NI2, pass, PEGB0
			10'd21 : rdata = 48'b110001010000001000000000000000000000000010000000;
			// PEs: 6 -> 0
			// srcs: (139, 25)(2010) -2 --> (2010) -2:NI3, pass, PEGB0
			10'd22 : rdata = 48'b110001010000001100000000000000000000000010000000;
			// PEs: 6 -> 0
			// srcs: (153, 21)(2064) -3 --> (2064) -3:NI1, pass, PEGB0
			10'd23 : rdata = 48'b110001010000000100000000000000000000000010000000;
			// PEs: 6 -> 0
			// srcs: (159, 26)(2194) -1 --> (2194) -1:NI4, pass, PEGB0
			10'd24 : rdata = 48'b110001010000010000000000000000000000000010000000;
			// PEs: 0 -> 
			// srcs: (556, 23)(1974) 6 --> (1974) 6:PEGB0, pass, 
			10'd25 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 1, 6 -> 6
			// srcs: (558, 24)(2754) -8, (1974) 6 --> (2755) -2:PEGB1, ALU, +, NI0
			10'd26 : rdata = 48'b000011110000001000111111111100000000000000000000;
			// PEs: 6 -> 1
			// srcs: (596, 27)(3077) -2 --> (3077) -2:NI5, pass, PEGB1
			10'd27 : rdata = 48'b110001010000010100000000000000000000000010010000;
			// PEs: 6 -> 1
			// srcs: (971, 28)(2755) -2 --> (2755) -2:NI0, pass, PEGB1
			10'd28 : rdata = 48'b110001010000000000000000000000000000000010010000;
			// PEs: 0, 6 -> 6
			// srcs: (1520, 29)(3140) 47, (9) 2 --> (3146) 94:PEGB0, ND0, *, NI0
			10'd29 : rdata = 48'b000111110000000001100000000100000000000000000000;
			// PEs: 6, 5 -> 5
			// srcs: (1522, 43)(3) 1, (3145) 94 --> (3929) 94:NM0, PENB, *, PEGB5
			10'd30 : rdata = 48'b000111000000000011011111110000000000000011010000;
			// PEs: 6, 6 -> 
			// srcs: (1523, 44)(3) 1, (3146) 94 --> (3930) 94:NM0, NI0, *, 
			10'd31 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 6, 6 -> 6
			// srcs: (1526, 60)(794) -3, (3930) 94 --> (4714) -97:NW0, ALU, -, NW0
			10'd32 : rdata = 48'b000100100000000000111111111000000100000000000000;
			// PEs: 0, 6 -> 
			// srcs: (1587, 30)(3140) 47, (77) 0 --> (3214) 0:PEGB0, ND10, *, 
			10'd33 : rdata = 48'b000111110000000001100001010000000000000000000000;
			// PEs: 6, 6 -> 
			// srcs: (1590, 45)(3) 1, (3214) 0 --> (3998) 0:NM0, ALU, *, 
			10'd34 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 6, 6 -> 6
			// srcs: (1593, 61)(862) -3, (3998) 0 --> (4782) -3:NW10, ALU, -, NW10
			10'd35 : rdata = 48'b000100100000101000111111111000000110100000000000;
			// PEs: 0, 6 -> 
			// srcs: (1601, 31)(3140) 47, (91) 0 --> (3228) 0:PEGB0, ND1, *, 
			10'd36 : rdata = 48'b000111110000000001100000001000000000000000000000;
			// PEs: 6, 6 -> 
			// srcs: (1604, 46)(3) 1, (3228) 0 --> (4012) 0:NM0, ALU, *, 
			10'd37 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 6, 6 -> 6
			// srcs: (1607, 62)(876) -1, (4012) 0 --> (4796) -1:NW1, ALU, -, NW1
			10'd38 : rdata = 48'b000100100000000100111111111000000100010000000000;
			// PEs: 0, 6 -> 7
			// srcs: (1681, 32)(3140) 47, (171) 0 --> (3308) 0:PEGB0, ND2, *, PENB
			10'd39 : rdata = 48'b000111110000000001100000010000000000000100000000;
			// PEs: 6, 5 -> 5
			// srcs: (1683, 47)(3) 1, (3307) -47 --> (4091) -47:NM0, PENB, *, PEGB5
			10'd40 : rdata = 48'b000111000000000011011111110000000000000011010000;
			// PEs: 6, 7 -> 6
			// srcs: (1690, 63)(956) 1, (4092) 0 --> (4876) 1:NW2, PEGB7, -, NW2
			10'd41 : rdata = 48'b000100100000001011100001110000000100100000000000;
			// PEs: 0, 6 -> 6
			// srcs: (1762, 33)(3140) 47, (252) 0 --> (3389) 0:PEGB0, ND3, *, NI0
			10'd42 : rdata = 48'b000111110000000001100000011100000000000000000000;
			// PEs: 6, 5 -> 5
			// srcs: (1764, 48)(3) 1, (3388) 47 --> (4172) 47:NM0, PENB, *, PEGB5
			10'd43 : rdata = 48'b000111000000000011011111110000000000000011010000;
			// PEs: 6, 6 -> 
			// srcs: (1765, 49)(3) 1, (3389) 0 --> (4173) 0:NM0, NI0, *, 
			10'd44 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 6, 6 -> 6
			// srcs: (1768, 64)(1037) 2, (4173) 0 --> (4957) 2:NW3, ALU, -, NW3
			10'd45 : rdata = 48'b000100100000001100111111111000000100110000000000;
			// PEs: 0, 6 -> 
			// srcs: (1771, 34)(3140) 47, (261) -1 --> (3398) -47:PEGB0, ND11, *, 
			10'd46 : rdata = 48'b000111110000000001100001011000000000000000000000;
			// PEs: 6, 6 -> 
			// srcs: (1774, 50)(3) 1, (3398) -47 --> (4182) -47:NM0, ALU, *, 
			10'd47 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 6, 6 -> 6
			// srcs: (1777, 65)(1046) 0, (4182) -47 --> (4966) 47:NW11, ALU, -, NW11
			10'd48 : rdata = 48'b000100100000101100111111111000000110110000000000;
			// PEs: 0, 6 -> 
			// srcs: (1843, 35)(3140) 47, (333) 2 --> (3470) 94:PEGB0, ND4, *, 
			10'd49 : rdata = 48'b000111110000000001100000100000000000000000000000;
			// PEs: 6, 6 -> 
			// srcs: (1846, 51)(3) 1, (3470) 94 --> (4254) 94:NM0, ALU, *, 
			10'd50 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 6, 6 -> 6
			// srcs: (1849, 66)(1118) -3, (4254) 94 --> (5038) -97:NW4, ALU, -, NW4
			10'd51 : rdata = 48'b000100100000010000111111111000000101000000000000;
			// PEs: 0, 6 -> 
			// srcs: (1923, 36)(3140) 47, (413) -1 --> (3550) -47:PEGB0, ND5, *, 
			10'd52 : rdata = 48'b000111110000000001100000101000000000000000000000;
			// PEs: 6, 6 -> 
			// srcs: (1926, 52)(3) 1, (3550) -47 --> (4334) -47:NM0, ALU, *, 
			10'd53 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 6, 6 -> 6
			// srcs: (1929, 67)(1198) 0, (4334) -47 --> (5118) 47:NW5, ALU, -, NW5
			10'd54 : rdata = 48'b000100100000010100111111111000000101010000000000;
			// PEs: 0, 6 -> 
			// srcs: (1951, 37)(3140) 47, (441) 2 --> (3578) 94:PEGB0, ND12, *, 
			10'd55 : rdata = 48'b000111110000000001100001100000000000000000000000;
			// PEs: 6, 6 -> 
			// srcs: (1954, 53)(3) 1, (3578) 94 --> (4362) 94:NM0, ALU, *, 
			10'd56 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 6, 6 -> 6
			// srcs: (1957, 68)(1226) -1, (4362) 94 --> (5146) -95:NW12, ALU, -, NW12
			10'd57 : rdata = 48'b000100100000110000111111111000000111000000000000;
			// PEs: 0, 6 -> 
			// srcs: (2005, 38)(3140) 47, (495) -3 --> (3632) -141:PEGB0, ND6, *, 
			10'd58 : rdata = 48'b000111110000000001100000110000000000000000000000;
			// PEs: 6, 6 -> 
			// srcs: (2008, 54)(3) 1, (3632) -141 --> (4416) -141:NM0, ALU, *, 
			10'd59 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 6, 6 -> 6
			// srcs: (2011, 69)(1280) 1, (4416) -141 --> (5200) 142:NW6, ALU, -, NW6
			10'd60 : rdata = 48'b000100100000011000111111111000000101100000000000;
			// PEs: 0, 6 -> 7
			// srcs: (2085, 39)(3140) 47, (575) 2 --> (3712) 94:PEGB0, ND7, *, PENB
			10'd61 : rdata = 48'b000111110000000001100000111000000000000100000000;
			// PEs: 6, 5 -> 5
			// srcs: (2087, 55)(3) 1, (3711) -94 --> (4495) -94:NM0, PENB, *, PEGB5
			10'd62 : rdata = 48'b000111000000000011011111110000000000000011010000;
			// PEs: 6, 7 -> 6
			// srcs: (2094, 70)(1360) 0, (4496) 94 --> (5280) -94:NW7, PEGB7, -, NW7
			10'd63 : rdata = 48'b000100100000011111100001110000000101110000000000;
			// PEs: 0, 6 -> 
			// srcs: (2135, 40)(3140) 47, (625) -1 --> (3762) -47:PEGB0, ND13, *, 
			10'd64 : rdata = 48'b000111110000000001100001101000000000000000000000;
			// PEs: 6, 6 -> 
			// srcs: (2138, 56)(3) 1, (3762) -47 --> (4546) -47:NM0, ALU, *, 
			10'd65 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 6, 6 -> 6
			// srcs: (2141, 71)(1410) 1, (4546) -47 --> (5330) 48:NW13, ALU, -, NW13
			10'd66 : rdata = 48'b000100100000110100111111111000000111010000000000;
			// PEs: 0, 6 -> 6
			// srcs: (2165, 41)(3140) 47, (655) 1 --> (3792) 47:PEGB0, ND8, *, NI0
			10'd67 : rdata = 48'b000111110000000001100001000100000000000000000000;
			// PEs: 6, 5 -> 5
			// srcs: (2167, 57)(3) 1, (3791) 47 --> (4575) 47:NM0, PENB, *, PEGB5
			10'd68 : rdata = 48'b000111000000000011011111110000000000000011010000;
			// PEs: 6, 6 -> 
			// srcs: (2168, 58)(3) 1, (3792) 47 --> (4576) 47:NM0, NI0, *, 
			10'd69 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 6, 6 -> 6
			// srcs: (2171, 72)(1440) 0, (4576) 47 --> (5360) -47:NW8, ALU, -, NW8
			10'd70 : rdata = 48'b000100100000100000111111111000000110000000000000;
			// PEs: 0, 6 -> 
			// srcs: (2247, 42)(3140) 47, (737) -2 --> (3874) -94:PEGB0, ND9, *, 
			10'd71 : rdata = 48'b000111110000000001100001001000000000000000000000;
			// PEs: 6, 6 -> 
			// srcs: (2250, 59)(3) 1, (3874) -94 --> (4658) -94:NM0, ALU, *, 
			10'd72 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 6, 6 -> 6
			// srcs: (2253, 73)(1522) 2, (4658) -94 --> (5442) 96:NW9, ALU, -, NW9
			10'd73 : rdata = 48'b000100100000100100111111111000000110010000000000;
			default : rdata = 48'b000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 7) begin
	always @(*) begin
		case(address)
			// PEs: 7, 7 -> 2
			// srcs: (1, 0)(11) 2, (796) -3 --> (1580) -6:ND0, NW0, *, PEGB2
			10'd0 : rdata = 48'b000110110000000001000000000000000000000010100000;
			// PEs: 7, 7 -> 1
			// srcs: (2, 1)(93) 1, (878) -3 --> (1662) -3:ND1, NW1, *, PEGB1
			10'd1 : rdata = 48'b000110110000000101000000001000000000000010010000;
			// PEs: 7, 7 -> 1
			// srcs: (3, 2)(173) -3, (958) -1 --> (1742) 3:ND2, NW2, *, PEGB1
			10'd2 : rdata = 48'b000110110000001001000000010000000000000010010000;
			// PEs: 7, 7 -> 0
			// srcs: (4, 3)(253) 0, (1038) 2 --> (1822) 0:ND3, NW3, *, PENB
			10'd3 : rdata = 48'b000110110000001101000000011000000000000100000000;
			// PEs: 7, 7 -> 0
			// srcs: (5, 4)(335) 2, (1120) -1 --> (1904) -2:ND4, NW4, *, PENB
			10'd4 : rdata = 48'b000110110000010001000000100000000000000100000000;
			// PEs: 7, 7 -> 0
			// srcs: (6, 5)(415) 1, (1200) -3 --> (1984) -3:ND5, NW5, *, PENB
			10'd5 : rdata = 48'b000110110000010101000000101000000000000100000000;
			// PEs: 7, 7 -> 7
			// srcs: (7, 6)(496) -1, (1281) 0 --> (2065) 0:ND6, NW6, *, NI0
			10'd6 : rdata = 48'b000110110000011001000000110100000000000000000000;
			// PEs: 7, 7 -> 0
			// srcs: (8, 7)(577) -2, (1362) 2 --> (2146) -4:ND7, NW7, *, PENB
			10'd7 : rdata = 48'b000110110000011101000000111000000000000100000000;
			// PEs: 7, 7 -> 0
			// srcs: (9, 8)(657) 0, (1442) 1 --> (2226) 0:ND8, NW8, *, PENB
			10'd8 : rdata = 48'b000110110000100001000001000000000000000100000000;
			// PEs: 7, 7 -> 7
			// srcs: (10, 9)(739) -2, (1524) -3 --> (2308) 6:ND9, NW9, *, NI1
			10'd9 : rdata = 48'b000110110000100101000001001100001000000000000000;
			// PEs: 7, 7 -> 7
			// srcs: (11, 10)(80) 2, (865) 0 --> (1649) 0:ND10, NW10, *, NI2
			10'd10 : rdata = 48'b000110110000101001000001010100010000000000000000;
			// PEs: 7, 7 -> 7
			// srcs: (12, 11)(264) 1, (1049) 0 --> (1833) 0:ND11, NW11, *, NI3
			10'd11 : rdata = 48'b000110110000101101000001011100011000000000000000;
			// PEs: 7, 7 -> 7
			// srcs: (13, 12)(444) -2, (1229) -1 --> (2013) 2:ND12, NW12, *, NI4
			10'd12 : rdata = 48'b000110110000110001000001100100100000000000000000;
			// PEs: 7, 7 -> 7
			// srcs: (14, 13)(628) 1, (1413) 0 --> (2197) 0:ND13, NW13, *, NI5
			10'd13 : rdata = 48'b000110110000110101000001101100101000000000000000;
			// PEs: 5, 6 -> 7
			// srcs: (15, 18)(2223) 0, (2224) 0 --> (3003) 0:PEGB5, PENB, +, NI6
			10'd14 : rdata = 48'b000011110000101011011111110100110000000000000000;
			// PEs: 5, 6 -> 7
			// srcs: (16, 19)(2305) 0, (2306) -4 --> (3082) -4:PEGB5, PENB, +, NI7
			10'd15 : rdata = 48'b000011110000101011011111110100111000000000000000;
			// PEs: 0 -> 
			// srcs: (26, 14)(1596) -6 --> (1596) -6:PEGB0, pass, 
			10'd16 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 0, 7 -> 0
			// srcs: (35, 15)(1595) 0, (1596) -6 --> (2376) -6:PEGB0, ALU, +, PENB
			10'd17 : rdata = 48'b000011110000000000111111111000000000000100000000;
			// PEs: 0 -> 
			// srcs: (59, 16)(1810) 3 --> (1810) 3:PEGB0, pass, 
			10'd18 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 0, 7 -> 5
			// srcs: (68, 17)(1809) 3, (1810) 3 --> (2589) 6:PEGB0, ALU, +, PEGB5
			10'd19 : rdata = 48'b000011110000000000111111111000000000000011010000;
			// PEs: 7 -> 0
			// srcs: (131, 22)(1649) 0 --> (1649) 0:NI2, pass, PENB
			10'd20 : rdata = 48'b110001010000001000000000000000000000000100000000;
			// PEs: 7 -> 0
			// srcs: (149, 24)(2013) 2 --> (2013) 2:NI4, pass, PENB
			10'd21 : rdata = 48'b110001010000010000000000000000000000000100000000;
			// PEs: 7 -> 0
			// srcs: (156, 23)(1833) 0 --> (1833) 0:NI3, pass, PENB
			10'd22 : rdata = 48'b110001010000001100000000000000000000000100000000;
			// PEs: 7 -> 0
			// srcs: (161, 20)(2065) 0 --> (2065) 0:NI0, pass, PENB
			10'd23 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 7 -> 0
			// srcs: (166, 21)(2308) 6 --> (2308) 6:NI1, pass, PENB
			10'd24 : rdata = 48'b110001010000000100000000000000000000000100000000;
			// PEs: 7 -> 0
			// srcs: (171, 26)(3003) 0 --> (3003) 0:NI6, pass, PENB
			10'd25 : rdata = 48'b110001010000011000000000000000000000000100000000;
			// PEs: 7 -> 0
			// srcs: (201, 25)(2197) 0 --> (2197) 0:NI5, pass, PENB
			10'd26 : rdata = 48'b110001010000010100000000000000000000000100000000;
			// PEs: 7 -> 0
			// srcs: (206, 27)(3082) -4 --> (3082) -4:NI7, pass, PENB
			10'd27 : rdata = 48'b110001010000011100000000000000000000000100000000;
			// PEs: 0 -> 
			// srcs: (1167, 28)(2580) -21 --> (2580) -21:PEGB0, pass, 
			10'd28 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 7, 1 -> 0
			// srcs: (1169, 29)(2580) -21, (2585) -3 --> (2586) -24:ALU, PEGB1, +, PENB
			10'd29 : rdata = 48'b000010011111111111100000010000000000000100000000;
			// PEs: 0, 7 -> 
			// srcs: (1522, 30)(3140) 47, (11) 2 --> (3148) 94:PEGB0, ND0, *, 
			10'd30 : rdata = 48'b000111110000000001100000000000000000000000000000;
			// PEs: 7, 7 -> 
			// srcs: (1525, 44)(3) 1, (3148) 94 --> (3932) 94:NM0, ALU, *, 
			10'd31 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 7, 7 -> 7
			// srcs: (1528, 60)(796) -3, (3932) 94 --> (4716) -97:NW0, ALU, -, NW0
			10'd32 : rdata = 48'b000100100000000000111111111000000100000000000000;
			// PEs: 0, 7 -> 
			// srcs: (1590, 31)(3140) 47, (80) 2 --> (3217) 94:PEGB0, ND10, *, 
			10'd33 : rdata = 48'b000111110000000001100001010000000000000000000000;
			// PEs: 7, 7 -> 
			// srcs: (1593, 45)(3) 1, (3217) 94 --> (4001) 94:NM0, ALU, *, 
			10'd34 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 7, 7 -> 7
			// srcs: (1596, 61)(865) 0, (4001) 94 --> (4785) -94:NW10, ALU, -, NW10
			10'd35 : rdata = 48'b000100100000101000111111111000000110100000000000;
			// PEs: 0, 7 -> 
			// srcs: (1603, 32)(3140) 47, (93) 1 --> (3230) 47:PEGB0, ND1, *, 
			10'd36 : rdata = 48'b000111110000000001100000001000000000000000000000;
			// PEs: 7, 7 -> 
			// srcs: (1606, 46)(3) 1, (3230) 47 --> (4014) 47:NM0, ALU, *, 
			10'd37 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 7, 7 -> 7
			// srcs: (1609, 62)(878) -3, (4014) 47 --> (4798) -50:NW1, ALU, -, NW1
			10'd38 : rdata = 48'b000100100000000100111111111000000100010000000000;
			// PEs: 0, 7 -> 7
			// srcs: (1683, 33)(3140) 47, (173) -3 --> (3310) -141:PEGB0, ND2, *, NI0
			10'd39 : rdata = 48'b000111110000000001100000010100000000000000000000;
			// PEs: 7, 6 -> 6
			// srcs: (1684, 47)(3) 1, (3308) 0 --> (4092) 0:NM0, PENB, *, PEGB6
			10'd40 : rdata = 48'b000111000000000011011111110000000000000011100000;
			// PEs: 7, 7 -> 
			// srcs: (1686, 48)(3) 1, (3310) -141 --> (4094) -141:NM0, NI0, *, 
			10'd41 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 7, 7 -> 7
			// srcs: (1689, 63)(958) -1, (4094) -141 --> (4878) 140:NW2, ALU, -, NW2
			10'd42 : rdata = 48'b000100100000001000111111111000000100100000000000;
			// PEs: 0, 7 -> 
			// srcs: (1763, 34)(3140) 47, (253) 0 --> (3390) 0:PEGB0, ND3, *, 
			10'd43 : rdata = 48'b000111110000000001100000011000000000000000000000;
			// PEs: 7, 7 -> 
			// srcs: (1766, 49)(3) 1, (3390) 0 --> (4174) 0:NM0, ALU, *, 
			10'd44 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 7, 7 -> 7
			// srcs: (1769, 64)(1038) 2, (4174) 0 --> (4958) 2:NW3, ALU, -, NW3
			10'd45 : rdata = 48'b000100100000001100111111111000000100110000000000;
			// PEs: 0, 7 -> 
			// srcs: (1774, 35)(3140) 47, (264) 1 --> (3401) 47:PEGB0, ND11, *, 
			10'd46 : rdata = 48'b000111110000000001100001011000000000000000000000;
			// PEs: 7, 7 -> 
			// srcs: (1777, 50)(3) 1, (3401) 47 --> (4185) 47:NM0, ALU, *, 
			10'd47 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 7, 7 -> 7
			// srcs: (1780, 65)(1049) 0, (4185) 47 --> (4969) -47:NW11, ALU, -, NW11
			10'd48 : rdata = 48'b000100100000101100111111111000000110110000000000;
			// PEs: 0, 7 -> 
			// srcs: (1845, 36)(3140) 47, (335) 2 --> (3472) 94:PEGB0, ND4, *, 
			10'd49 : rdata = 48'b000111110000000001100000100000000000000000000000;
			// PEs: 7, 7 -> 
			// srcs: (1848, 51)(3) 1, (3472) 94 --> (4256) 94:NM0, ALU, *, 
			10'd50 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 7, 7 -> 7
			// srcs: (1851, 66)(1120) -1, (4256) 94 --> (5040) -95:NW4, ALU, -, NW4
			10'd51 : rdata = 48'b000100100000010000111111111000000101000000000000;
			// PEs: 0, 7 -> 
			// srcs: (1925, 37)(3140) 47, (415) 1 --> (3552) 47:PEGB0, ND5, *, 
			10'd52 : rdata = 48'b000111110000000001100000101000000000000000000000;
			// PEs: 7, 7 -> 
			// srcs: (1928, 52)(3) 1, (3552) 47 --> (4336) 47:NM0, ALU, *, 
			10'd53 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 7, 7 -> 7
			// srcs: (1931, 67)(1200) -3, (4336) 47 --> (5120) -50:NW5, ALU, -, NW5
			10'd54 : rdata = 48'b000100100000010100111111111000000101010000000000;
			// PEs: 0, 7 -> 
			// srcs: (1954, 38)(3140) 47, (444) -2 --> (3581) -94:PEGB0, ND12, *, 
			10'd55 : rdata = 48'b000111110000000001100001100000000000000000000000;
			// PEs: 7, 7 -> 
			// srcs: (1957, 53)(3) 1, (3581) -94 --> (4365) -94:NM0, ALU, *, 
			10'd56 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 7, 7 -> 7
			// srcs: (1960, 68)(1229) -1, (4365) -94 --> (5149) 93:NW12, ALU, -, NW12
			10'd57 : rdata = 48'b000100100000110000111111111000000111000000000000;
			// PEs: 0, 7 -> 
			// srcs: (2006, 39)(3140) 47, (496) -1 --> (3633) -47:PEGB0, ND6, *, 
			10'd58 : rdata = 48'b000111110000000001100000110000000000000000000000;
			// PEs: 7, 7 -> 
			// srcs: (2009, 54)(3) 1, (3633) -47 --> (4417) -47:NM0, ALU, *, 
			10'd59 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 7, 7 -> 7
			// srcs: (2012, 69)(1281) 0, (4417) -47 --> (5201) 47:NW6, ALU, -, NW6
			10'd60 : rdata = 48'b000100100000011000111111111000000101100000000000;
			// PEs: 0, 7 -> 7
			// srcs: (2087, 40)(3140) 47, (577) -2 --> (3714) -94:PEGB0, ND7, *, NI0
			10'd61 : rdata = 48'b000111110000000001100000111100000000000000000000;
			// PEs: 7, 6 -> 6
			// srcs: (2088, 55)(3) 1, (3712) 94 --> (4496) 94:NM0, PENB, *, PEGB6
			10'd62 : rdata = 48'b000111000000000011011111110000000000000011100000;
			// PEs: 7, 7 -> 
			// srcs: (2090, 56)(3) 1, (3714) -94 --> (4498) -94:NM0, NI0, *, 
			10'd63 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 7, 7 -> 7
			// srcs: (2093, 70)(1362) 2, (4498) -94 --> (5282) 96:NW7, ALU, -, NW7
			10'd64 : rdata = 48'b000100100000011100111111111000000101110000000000;
			// PEs: 0, 7 -> 
			// srcs: (2138, 41)(3140) 47, (628) 1 --> (3765) 47:PEGB0, ND13, *, 
			10'd65 : rdata = 48'b000111110000000001100001101000000000000000000000;
			// PEs: 7, 7 -> 
			// srcs: (2141, 57)(3) 1, (3765) 47 --> (4549) 47:NM0, ALU, *, 
			10'd66 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 7, 7 -> 7
			// srcs: (2144, 71)(1413) 0, (4549) 47 --> (5333) -47:NW13, ALU, -, NW13
			10'd67 : rdata = 48'b000100100000110100111111111000000111010000000000;
			// PEs: 0, 7 -> 
			// srcs: (2167, 42)(3140) 47, (657) 0 --> (3794) 0:PEGB0, ND8, *, 
			10'd68 : rdata = 48'b000111110000000001100001000000000000000000000000;
			// PEs: 7, 7 -> 
			// srcs: (2170, 58)(3) 1, (3794) 0 --> (4578) 0:NM0, ALU, *, 
			10'd69 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 7, 7 -> 7
			// srcs: (2173, 72)(1442) 1, (4578) 0 --> (5362) 1:NW8, ALU, -, NW8
			10'd70 : rdata = 48'b000100100000100000111111111000000110000000000000;
			// PEs: 0, 7 -> 
			// srcs: (2249, 43)(3140) 47, (739) -2 --> (3876) -94:PEGB0, ND9, *, 
			10'd71 : rdata = 48'b000111110000000001100001001000000000000000000000;
			// PEs: 7, 7 -> 
			// srcs: (2252, 59)(3) 1, (3876) -94 --> (4660) -94:NM0, ALU, *, 
			10'd72 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 7, 7 -> 7
			// srcs: (2255, 73)(1524) -3, (4660) -94 --> (5444) 91:NW9, ALU, -, NW9
			10'd73 : rdata = 48'b000100100000100100111111111000000110010000000000;
			default : rdata = 48'b000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 8) begin
	always @(*) begin
		case(address)
			// PEs: 9 -> 0
			// srcs: (6, 0)(1581) 1 --> (1581) 1:PEGB1, pass, PUGB0
			10'd0 : rdata = 48'b110001110000001000000000000000000000000000001000;
			// PEs: 10 -> 0
			// srcs: (7, 1)(1583) -4 --> (1583) -4:PEGB2, pass, PUGB0
			10'd1 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 11 -> 0
			// srcs: (8, 2)(1584) -4 --> (1584) -4:PEGB3, pass, PUGB0
			10'd2 : rdata = 48'b110001110000011000000000000000000000000000001000;
			// PEs: 12 -> 0
			// srcs: (9, 3)(1586) -4 --> (1586) -4:PEGB4, pass, PUGB0
			10'd3 : rdata = 48'b110001110000100000000000000000000000000000001000;
			// PEs: 13 -> 0
			// srcs: (10, 4)(1587) 3 --> (1587) 3:PEGB5, pass, PUGB0
			10'd4 : rdata = 48'b110001110000101000000000000000000000000000001000;
			// PEs: 14 -> 0
			// srcs: (11, 5)(1589) 6 --> (1589) 6:PEGB6, pass, PUGB0
			10'd5 : rdata = 48'b110001110000110000000000000000000000000000001000;
			// PEs: 15 -> 0
			// srcs: (12, 6)(1590) 3 --> (1590) 3:PENB, pass, PUGB0
			10'd6 : rdata = 48'b110001101111111000000000000000000000000000001000;
			// PEs: 24 -> 8
			// srcs: (13, 11)(1602) -4 --> (1602) -4:PUGB3, pass, NI0
			10'd7 : rdata = 48'b110001110000011100000000000100000000000000000000;
			// PEs: 24 -> 8
			// srcs: (14, 13)(1604) -1 --> (1604) -1:PUGB3, pass, NI1
			10'd8 : rdata = 48'b110001110000011100000000000100001000000000000000;
			// PEs: 16 -> 8
			// srcs: (15, 7)(1598) 4 --> (1598) 4:PUGB2, pass, NI2
			10'd9 : rdata = 48'b110001110000010100000000000100010000000000000000;
			// PEs: 24 -> 12
			// srcs: (16, 14)(1605) -2 --> (1605) -2:PUGB3, pass, PEGB4
			10'd10 : rdata = 48'b110001110000011100000000000000000000000011000000;
			// PEs: 24 -> 8
			// srcs: (17, 16)(1607) -2 --> (1607) -2:PUGB3, pass, NI3
			10'd11 : rdata = 48'b110001110000011100000000000100011000000000000000;
			// PEs: 16 -> 10
			// srcs: (18, 8)(1599) -2 --> (1599) -2:PUGB2, pass, PEGB2
			10'd12 : rdata = 48'b110001110000010100000000000000000000000010100000;
			// PEs: 16 -> 11
			// srcs: (19, 10)(1601) 4 --> (1601) 4:PUGB2, pass, PEGB3
			10'd13 : rdata = 48'b110001110000010100000000000000000000000010110000;
			// PEs: 24 -> 13
			// srcs: (20, 17)(1608) 0 --> (1608) 0:PUGB3, pass, PEGB5
			10'd14 : rdata = 48'b110001110000011100000000000000000000000011010000;
			// PEs: 24 -> 8
			// srcs: (21, 19)(1610) -6 --> (1610) -6:PUGB3, pass, NI4
			10'd15 : rdata = 48'b110001110000011100000000000100100000000000000000;
			// PEs: 24 -> 14
			// srcs: (22, 20)(1611) -2 --> (1611) -2:PUGB3, pass, PEGB6
			10'd16 : rdata = 48'b110001110000011100000000000000000000000011100000;
			// PEs: 32 -> 8
			// srcs: (23, 22)(1613) 0 --> (1613) 0:PUGB4, pass, NI5
			10'd17 : rdata = 48'b110001110000100100000000000100101000000000000000;
			// PEs: 32 -> 15
			// srcs: (24, 23)(1614) 6 --> (1614) 6:PUGB4, pass, PEGB7
			10'd18 : rdata = 48'b110001110000100100000000000000000000000011110000;
			// PEs: 8 -> 12
			// srcs: (25, 15)(1604) -1 --> (1604) -1:NI1, pass, PEGB4
			10'd19 : rdata = 48'b110001010000000100000000000000000000000011000000;
			// PEs: 9 -> 0
			// srcs: (26, 25)(1663) -3 --> (1663) -3:PEGB1, pass, PUGB0
			10'd20 : rdata = 48'b110001110000001000000000000000000000000000001000;
			// PEs: 8 -> 10
			// srcs: (27, 9)(1598) 4 --> (1598) 4:NI2, pass, PEGB2
			10'd21 : rdata = 48'b110001010000001000000000000000000000000010100000;
			// PEs: 8 -> 11
			// srcs: (28, 12)(1602) -4 --> (1602) -4:NI0, pass, PEGB3
			10'd22 : rdata = 48'b110001010000000000000000000000000000000010110000;
			// PEs: 8 -> 13
			// srcs: (29, 18)(1607) -2 --> (1607) -2:NI3, pass, PEGB5
			10'd23 : rdata = 48'b110001010000001100000000000000000000000011010000;
			// PEs: 10 -> 40
			// srcs: (30, 26)(1665) -1 --> (1665) -1:PEGB2, pass, PUGB5
			10'd24 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 8 -> 14
			// srcs: (31, 21)(1610) -6 --> (1610) -6:NI4, pass, PEGB6
			10'd25 : rdata = 48'b110001010000010000000000000000000000000011100000;
			// PEs: 11 -> 40
			// srcs: (32, 27)(1666) 0 --> (1666) 0:PEGB3, pass, PUGB5
			10'd26 : rdata = 48'b110001110000011000000000000000000000000000001101;
			// PEs: 8 -> 15
			// srcs: (33, 24)(1613) 0 --> (1613) 0:NI5, pass, PEGB7
			10'd27 : rdata = 48'b110001010000010100000000000000000000000011110000;
			// PEs: 12 -> 48
			// srcs: (34, 28)(1668) 9 --> (1668) 9:PEGB4, pass, PUGB6
			10'd28 : rdata = 48'b110001110000100000000000000000000000000000001110;
			// PEs: 13 -> 48
			// srcs: (35, 29)(1669) 0 --> (1669) 0:PEGB5, pass, PUGB6
			10'd29 : rdata = 48'b110001110000101000000000000000000000000000001110;
			// PEs: 16 -> 8
			// srcs: (36, 30)(1675) 4 --> (1675) 4:PUGB2, pass, NI0
			10'd30 : rdata = 48'b110001110000010100000000000100000000000000000000;
			// PEs: 9 -> 0
			// srcs: (37, 42)(1743) 1 --> (1743) 1:PEGB1, pass, PUGB0
			10'd31 : rdata = 48'b110001110000001000000000000000000000000000001000;
			// PEs: 16 -> 9
			// srcs: (38, 31)(1676) -6 --> (1676) -6:PUGB2, pass, PENB
			10'd32 : rdata = 48'b110001110000010100000000000000000000000100000000;
			// PEs: 0 -> 8
			// srcs: (39, 33)(1733) 4 --> (1733) 4:PUNB, pass, NI1
			10'd33 : rdata = 48'b110001101111111100000000000100001000000000000000;
			// PEs: 0 -> 10
			// srcs: (40, 34)(1734) -1 --> (1734) -1:PUNB, pass, PEGB2
			10'd34 : rdata = 48'b110001101111111100000000000000000000000010100000;
			// PEs: 0 -> 8
			// srcs: (41, 36)(1736) -2 --> (1736) -2:PUNB, pass, NI2
			10'd35 : rdata = 48'b110001101111111100000000000100010000000000000000;
			// PEs: 0 -> 11
			// srcs: (42, 37)(1737) 0 --> (1737) 0:PUNB, pass, PEGB3
			10'd36 : rdata = 48'b110001101111111100000000000000000000000010110000;
			// PEs: 10 -> 0
			// srcs: (43, 43)(1745) 2 --> (1745) 2:PEGB2, pass, PUGB0
			10'd37 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 8 -> 9
			// srcs: (44, 32)(1675) 4 --> (1675) 4:NI0, pass, PENB
			10'd38 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 0 -> 8
			// srcs: (45, 39)(1739) -1 --> (1739) -1:PUNB, pass, NI0
			10'd39 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 0 -> 12
			// srcs: (46, 40)(1740) 0 --> (1740) 0:PUNB, pass, PEGB4
			10'd40 : rdata = 48'b110001101111111100000000000000000000000011000000;
			// PEs: 11 -> 0
			// srcs: (47, 44)(1746) -2 --> (1746) -2:PEGB3, pass, PUGB0
			10'd41 : rdata = 48'b110001110000011000000000000000000000000000001000;
			// PEs: 12 -> 16
			// srcs: (48, 45)(1748) -3 --> (1748) -3:PEGB4, pass, PUNB
			10'd42 : rdata = 48'b110001110000100000000000000000000000001000000000;
			// PEs: 8 -> 10
			// srcs: (49, 35)(1733) 4 --> (1733) 4:NI1, pass, PEGB2
			10'd43 : rdata = 48'b110001010000000100000000000000000000000010100000;
			// PEs: 13 -> 16
			// srcs: (50, 46)(1749) 2 --> (1749) 2:PEGB5, pass, PUNB
			10'd44 : rdata = 48'b110001110000101000000000000000000000001000000000;
			// PEs: 8 -> 11
			// srcs: (51, 38)(1736) -2 --> (1736) -2:NI2, pass, PEGB3
			10'd45 : rdata = 48'b110001010000001000000000000000000000000010110000;
			// PEs: 14 -> 16
			// srcs: (52, 47)(1751) 0 --> (1751) 0:PEGB6, pass, PUNB
			10'd46 : rdata = 48'b110001110000110000000000000000000000001000000000;
			// PEs: 15 -> 16
			// srcs: (53, 48)(1752) 2 --> (1752) 2:PENB, pass, PUNB
			10'd47 : rdata = 48'b110001101111111000000000000000000000001000000000;
			// PEs: 16 -> 8
			// srcs: (54, 49)(1754) 0 --> (1754) 0:PUGB2, pass, NI1
			10'd48 : rdata = 48'b110001110000010100000000000100001000000000000000;
			// PEs: 8 -> 12
			// srcs: (55, 41)(1739) -1 --> (1739) -1:NI0, pass, PEGB4
			10'd49 : rdata = 48'b110001010000000000000000000000000000000011000000;
			// PEs: 16 -> 9
			// srcs: (56, 50)(1755) -4 --> (1755) -4:PUGB2, pass, PENB
			10'd50 : rdata = 48'b110001110000010100000000000000000000000100000000;
			// PEs: 0 -> 8
			// srcs: (57, 52)(1815) -3 --> (1815) -3:PUNB, pass, NI0
			10'd51 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 0 -> 13
			// srcs: (58, 53)(1816) 0 --> (1816) 0:PUNB, pass, PEGB5
			10'd52 : rdata = 48'b110001101111111100000000000000000000000011010000;
			// PEs: 9 -> 16
			// srcs: (59, 55)(1823) 0 --> (1823) 0:PEGB1, pass, PUNB
			10'd53 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 10 -> 16
			// srcs: (60, 56)(1825) 1 --> (1825) 1:PEGB2, pass, PUNB
			10'd54 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 11 -> 16
			// srcs: (61, 57)(1826) -2 --> (1826) -2:PEGB3, pass, PUNB
			10'd55 : rdata = 48'b110001110000011000000000000000000000001000000000;
			// PEs: 8 -> 9
			// srcs: (62, 51)(1754) 0 --> (1754) 0:NI1, pass, PENB
			10'd56 : rdata = 48'b110001010000000100000000000000000000000100000000;
			// PEs: 12 -> 16
			// srcs: (63, 58)(1828) 0 --> (1828) 0:PEGB4, pass, PUNB
			10'd57 : rdata = 48'b110001110000100000000000000000000000001000000000;
			// PEs: 13 -> 16
			// srcs: (64, 59)(1829) 0 --> (1829) 0:PEGB5, pass, PUNB
			10'd58 : rdata = 48'b110001110000101000000000000000000000001000000000;
			// PEs: 14 -> 16
			// srcs: (65, 60)(1831) -3 --> (1831) -3:PEGB6, pass, PUNB
			10'd59 : rdata = 48'b110001110000110000000000000000000000001000000000;
			// PEs: 15 -> 16
			// srcs: (66, 61)(1832) 9 --> (1832) 9:PENB, pass, PUNB
			10'd60 : rdata = 48'b110001101111111000000000000000000000001000000000;
			// PEs: 8 -> 13
			// srcs: (67, 54)(1815) -3 --> (1815) -3:NI0, pass, PEGB5
			10'd61 : rdata = 48'b110001010000000000000000000000000000000011010000;
			// PEs: 0 -> 8
			// srcs: (68, 62)(1895) -4 --> (1895) -4:PUNB, pass, NI0
			10'd62 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 0 -> 9
			// srcs: (69, 63)(1896) -3 --> (1896) -3:PUNB, pass, PENB
			10'd63 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 10 -> 16
			// srcs: (70, 72)(1907) 0 --> (1907) 0:PEGB2, pass, PUNB
			10'd64 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 11 -> 16
			// srcs: (71, 73)(1908) -3 --> (1908) -3:PEGB3, pass, PUNB
			10'd65 : rdata = 48'b110001110000011000000000000000000000001000000000;
			// PEs: 12 -> 16
			// srcs: (72, 74)(1910) -2 --> (1910) -2:PEGB4, pass, PUNB
			10'd66 : rdata = 48'b110001110000100000000000000000000000001000000000;
			// PEs: 13 -> 16
			// srcs: (73, 75)(1911) 0 --> (1911) 0:PEGB5, pass, PUNB
			10'd67 : rdata = 48'b110001110000101000000000000000000000001000000000;
			// PEs: 14 -> 16
			// srcs: (74, 76)(1913) 2 --> (1913) 2:PEGB6, pass, PUNB
			10'd68 : rdata = 48'b110001110000110000000000000000000000001000000000;
			// PEs: 8 -> 9
			// srcs: (75, 64)(1895) -4 --> (1895) -4:NI0, pass, PENB
			10'd69 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 0 -> 8
			// srcs: (76, 65)(1898) 4 --> (1898) 4:PUNB, pass, NI0
			10'd70 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 0 -> 9
			// srcs: (77, 66)(1899) 0 --> (1899) 0:PUNB, pass, PENB
			10'd71 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 15 -> 16
			// srcs: (78, 77)(1914) -4 --> (1914) -4:PENB, pass, PUNB
			10'd72 : rdata = 48'b110001101111111000000000000000000000001000000000;
			// PEs: 10 -> 16
			// srcs: (79, 88)(1987) 4 --> (1987) 4:PEGB2, pass, PUNB
			10'd73 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 11 -> 16
			// srcs: (80, 89)(1988) -2 --> (1988) -2:PEGB3, pass, PUNB
			10'd74 : rdata = 48'b110001110000011000000000000000000000001000000000;
			// PEs: 12 -> 16
			// srcs: (81, 90)(1990) -2 --> (1990) -2:PEGB4, pass, PUNB
			10'd75 : rdata = 48'b110001110000100000000000000000000000001000000000;
			// PEs: 13 -> 16
			// srcs: (82, 91)(1991) 1 --> (1991) 1:PEGB5, pass, PUNB
			10'd76 : rdata = 48'b110001110000101000000000000000000000001000000000;
			// PEs: 8 -> 9
			// srcs: (83, 67)(1898) 4 --> (1898) 4:NI0, pass, PENB
			10'd77 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 0 -> 8
			// srcs: (84, 68)(1901) -2 --> (1901) -2:PUNB, pass, NI0
			10'd78 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 0 -> 9
			// srcs: (85, 69)(1902) -6 --> (1902) -6:PUNB, pass, PENB
			10'd79 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 0 -> 14
			// srcs: (86, 71)(1904) -2 --> (1904) -2:PUNB, pass, PEGB6
			10'd80 : rdata = 48'b110001101111111100000000000000000000000011100000;
			// PEs: 14 -> 16
			// srcs: (87, 92)(1993) 0 --> (1993) 0:PEGB6, pass, PUNB
			10'd81 : rdata = 48'b110001110000110000000000000000000000001000000000;
			// PEs: 15 -> 16
			// srcs: (88, 93)(1994) 0 --> (1994) 0:PENB, pass, PUNB
			10'd82 : rdata = 48'b110001101111111000000000000000000000001000000000;
			// PEs: 10 -> 16
			// srcs: (89, 100)(2067) -1 --> (2067) -1:PEGB2, pass, PUNB
			10'd83 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 11 -> 16
			// srcs: (90, 101)(2068) 0 --> (2068) 0:PEGB3, pass, PUNB
			10'd84 : rdata = 48'b110001110000011000000000000000000000001000000000;
			// PEs: 8 -> 9
			// srcs: (91, 70)(1901) -2 --> (1901) -2:NI0, pass, PENB
			10'd85 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 0 -> 8
			// srcs: (92, 78)(1975) -2 --> (1975) -2:PUNB, pass, NI0
			10'd86 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 0 -> 9
			// srcs: (93, 79)(1976) -3 --> (1976) -3:PUNB, pass, PENB
			10'd87 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 12 -> 16
			// srcs: (94, 102)(2070) 4 --> (2070) 4:PEGB4, pass, PUNB
			10'd88 : rdata = 48'b110001110000100000000000000000000000001000000000;
			// PEs: 13 -> 16
			// srcs: (95, 103)(2071) 2 --> (2071) 2:PEGB5, pass, PUNB
			10'd89 : rdata = 48'b110001110000101000000000000000000000001000000000;
			// PEs: 14 -> 16
			// srcs: (96, 104)(2073) 2 --> (2073) 2:PEGB6, pass, PUNB
			10'd90 : rdata = 48'b110001110000110000000000000000000000001000000000;
			// PEs: 15 -> 16
			// srcs: (97, 105)(2074) 4 --> (2074) 4:PENB, pass, PUNB
			10'd91 : rdata = 48'b110001101111111000000000000000000000001000000000;
			// PEs: 10 -> 16
			// srcs: (98, 116)(2149) 4 --> (2149) 4:PEGB2, pass, PUNB
			10'd92 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 8 -> 9
			// srcs: (99, 80)(1975) -2 --> (1975) -2:NI0, pass, PENB
			10'd93 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 0 -> 8
			// srcs: (100, 81)(1978) 0 --> (1978) 0:PUNB, pass, NI0
			10'd94 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 0 -> 9
			// srcs: (101, 82)(1979) 0 --> (1979) 0:PUNB, pass, PENB
			10'd95 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 11 -> 16
			// srcs: (102, 117)(2150) 1 --> (2150) 1:PEGB3, pass, PUNB
			10'd96 : rdata = 48'b110001110000011000000000000000000000001000000000;
			// PEs: 12 -> 16
			// srcs: (103, 118)(2152) 0 --> (2152) 0:PEGB4, pass, PUNB
			10'd97 : rdata = 48'b110001110000100000000000000000000000001000000000;
			// PEs: 13 -> 16
			// srcs: (104, 119)(2153) 4 --> (2153) 4:PEGB5, pass, PUNB
			10'd98 : rdata = 48'b110001110000101000000000000000000000001000000000;
			// PEs: 14 -> 16
			// srcs: (105, 120)(2155) 2 --> (2155) 2:PEGB6, pass, PUNB
			10'd99 : rdata = 48'b110001110000110000000000000000000000001000000000;
			// PEs: 15 -> 16
			// srcs: (106, 121)(2156) 2 --> (2156) 2:PENB, pass, PUNB
			10'd100 : rdata = 48'b110001101111111000000000000000000000001000000000;
			// PEs: 8 -> 9
			// srcs: (107, 83)(1978) 0 --> (1978) 0:NI0, pass, PENB
			10'd101 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 0 -> 8
			// srcs: (108, 84)(1981) -6 --> (1981) -6:PUNB, pass, NI0
			10'd102 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 0 -> 9
			// srcs: (109, 85)(1982) 0 --> (1982) 0:PUNB, pass, PENB
			10'd103 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 0 -> 15
			// srcs: (110, 87)(1984) -3 --> (1984) -3:PUNB, pass, PEGB7
			10'd104 : rdata = 48'b110001101111111100000000000000000000000011110000;
			// PEs: 12 -> 24
			// srcs: (111, 141)(2386) -3 --> (2386) -3:PEGB4, pass, PUGB3
			10'd105 : rdata = 48'b110001110000100000000000000000000000000000001011;
			// PEs: 13 -> 32
			// srcs: (112, 142)(2388) -2 --> (2388) -2:PEGB5, pass, PUGB4
			10'd106 : rdata = 48'b110001110000101000000000000000000000000000001100;
			// PEs: 14 -> 0
			// srcs: (113, 143)(2392) -8 --> (2392) -8:PEGB6, pass, PUGB0
			10'd107 : rdata = 48'b110001110000110000000000000000000000000000001000;
			// PEs: 15 -> 56
			// srcs: (114, 144)(2394) 6 --> (2394) 6:PENB, pass, PUGB7
			10'd108 : rdata = 48'b110001101111111000000000000000000000000000001111;
			// PEs: 8 -> 9
			// srcs: (115, 86)(1981) -6 --> (1981) -6:NI0, pass, PENB
			10'd109 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 0 -> 8
			// srcs: (116, 94)(2057) 0 --> (2057) 0:PUNB, pass, NI0
			10'd110 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 0 -> 9
			// srcs: (117, 95)(2058) 0 --> (2058) 0:PUNB, pass, PENB
			10'd111 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 14 -> 16
			// srcs: (118, 126)(1671) 2 --> (1671) 2:PEGB6, pass, PUNB
			10'd112 : rdata = 48'b110001110000110000000000000000000000001000000000;
			// PEs: 11 -> 40
			// srcs: (119, 151)(1658) 4 --> (1658) 4:PEGB3, pass, PUGB5
			10'd113 : rdata = 48'b110001110000011000000000000000000000000000001101;
			// PEs: 11 -> 40
			// srcs: (120, 164)(2516) -2 --> (2516) -2:PEGB3, pass, PUGB5
			10'd114 : rdata = 48'b110001110000011000000000000000000000000000001101;
			// PEs: 9 -> 40
			// srcs: (121, 174)(1836) 6 --> (1836) 6:PEGB1, pass, PUGB5
			10'd115 : rdata = 48'b110001110000001000000000000000000000000000001101;
			// PEs: 8 -> 9
			// srcs: (123, 96)(2057) 0 --> (2057) 0:NI0, pass, PENB
			10'd116 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 0 -> 8
			// srcs: (124, 97)(2060) -6 --> (2060) -6:PUNB, pass, NI0
			10'd117 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 0 -> 9
			// srcs: (125, 98)(2061) -2 --> (2061) -2:PUNB, pass, PENB
			10'd118 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 15 -> 16
			// srcs: (126, 127)(1672) 1 --> (1672) 1:PENB, pass, PUNB
			10'd119 : rdata = 48'b110001101111111000000000000000000000001000000000;
			// PEs: 10 -> 16
			// srcs: (127, 150)(1655) 6 --> (1655) 6:PEGB2, pass, PUNB
			10'd120 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 12 -> 48
			// srcs: (128, 152)(1661) 0 --> (1661) 0:PEGB4, pass, PUGB6
			10'd121 : rdata = 48'b110001110000100000000000000000000000000000001110;
			// PEs: 9 -> 16
			// srcs: (129, 156)(2457) -2 --> (2457) -2:PEGB1, pass, PUNB
			10'd122 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 10 -> 32
			// srcs: (130, 163)(2514) 3 --> (2514) 3:PEGB2, pass, PUGB4
			10'd123 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 8 -> 9
			// srcs: (131, 99)(2060) -6 --> (2060) -6:NI0, pass, PENB
			10'd124 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 0 -> 8
			// srcs: (132, 106)(2137) 0 --> (2137) 0:PUNB, pass, NI0
			10'd125 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 0 -> 9
			// srcs: (133, 107)(2138) 0 --> (2138) 0:PUNB, pass, PENB
			10'd126 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 15 -> 48
			// srcs: (134, 155)(1670) -6 --> (1670) -6:PENB, pass, PUGB6
			10'd127 : rdata = 48'b110001101111111000000000000000000000000000001110;
			// PEs: 9 -> 48
			// srcs: (135, 169)(2533) -4 --> (2533) -4:PEGB1, pass, PUGB6
			10'd128 : rdata = 48'b110001110000001000000000000000000000000000001110;
			// PEs: 12 -> 24
			// srcs: (136, 177)(1845) 0 --> (1845) 0:PEGB4, pass, PUGB3
			10'd129 : rdata = 48'b110001110000100000000000000000000000000000001011;
			// PEs: 14 -> 0
			// srcs: (137, 179)(1851) 0 --> (1851) 0:PEGB6, pass, PUGB0
			10'd130 : rdata = 48'b110001110000110000000000000000000000000000001000;
			// PEs: 8 -> 9
			// srcs: (139, 108)(2137) 0 --> (2137) 0:NI0, pass, PENB
			10'd131 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 0 -> 8
			// srcs: (140, 109)(2140) 2 --> (2140) 2:PUNB, pass, NI0
			10'd132 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 0 -> 9
			// srcs: (141, 110)(2141) -2 --> (2141) -2:PUNB, pass, PENB
			10'd133 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 15 -> 32
			// srcs: (142, 180)(1854) 0 --> (1854) 0:PENB, pass, PUGB4
			10'd134 : rdata = 48'b110001101111111000000000000000000000000000001100;
			// PEs: 10 -> 16
			// srcs: (143, 175)(1839) -6 --> (1839) -6:PEGB2, pass, PUNB
			10'd135 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 9 -> 16
			// srcs: (144, 185)(2678) 4 --> (2678) 4:PEGB1, pass, PUNB
			10'd136 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 9 -> 0
			// srcs: (145, 186)(2680) -8 --> (2680) -8:PEGB1, pass, PUGB0
			10'd137 : rdata = 48'b110001110000001000000000000000000000000000001000;
			// PEs: 11 -> 48
			// srcs: (146, 203)(2026) -1 --> (2026) -1:PEGB3, pass, PUGB6
			10'd138 : rdata = 48'b110001110000011000000000000000000000000000001110;
			// PEs: 8 -> 9
			// srcs: (147, 111)(2140) 2 --> (2140) 2:NI0, pass, PENB
			10'd139 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 0 -> 8
			// srcs: (148, 112)(2143) 0 --> (2143) 0:PUNB, pass, NI0
			10'd140 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 0 -> 9
			// srcs: (149, 113)(2144) 0 --> (2144) 0:PUNB, pass, PENB
			10'd141 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 15 -> 0
			// srcs: (150, 194)(2765) -4 --> (2765) -4:PENB, pass, PUGB0
			10'd142 : rdata = 48'b110001101111111000000000000000000000000000001000;
			// PEs: 10 -> 16
			// srcs: (153, 202)(2023) 1 --> (2023) 1:PEGB2, pass, PUNB
			10'd143 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 8 -> 9
			// srcs: (155, 114)(2143) 0 --> (2143) 0:NI0, pass, PENB
			10'd144 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 0 -> 9
			// srcs: (156, 115)(2146) -4 --> (2146) -4:PUNB, pass, PENB
			10'd145 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 0 -> 9
			// srcs: (157, 122)(2226) 0 --> (2226) 0:PUNB, pass, PENB
			10'd146 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 14 -> 32
			// srcs: (158, 206)(2035) -1 --> (2035) -1:PEGB6, pass, PUGB4
			10'd147 : rdata = 48'b110001110000110000000000000000000000000000001100;
			// PEs: 13 -> 16
			// srcs: (161, 205)(2032) 0 --> (2032) 0:PEGB5, pass, PUNB
			10'd148 : rdata = 48'b110001110000101000000000000000000000001000000000;
			// PEs: 40 -> 8
			// srcs: (196, 123)(1624) 0 --> (1624) 0:PUGB5, pass, NI0
			10'd149 : rdata = 48'b110001110000101100000000000100000000000000000000;
			// PEs: 40 -> 15
			// srcs: (213, 124)(1625) 4 --> (1625) 4:PUGB5, pass, PEGB7
			10'd150 : rdata = 48'b110001110000101100000000000000000000000011110000;
			// PEs: 0 -> 8
			// srcs: (220, 128)(1818) 2 --> (1818) 2:PUNB, pass, NI1
			10'd151 : rdata = 48'b110001101111111100000000000100001000000000000000;
			// PEs: 8 -> 15
			// srcs: (222, 125)(1624) 0 --> (1624) 0:NI0, pass, PEGB7
			10'd152 : rdata = 48'b110001010000000000000000000000000000000011110000;
			// PEs: 15 -> 56
			// srcs: (229, 145)(2406) 4 --> (2406) 4:PENB, pass, PUGB7
			10'd153 : rdata = 48'b110001101111111000000000000000000000000000001111;
			// PEs: 14 -> 56
			// srcs: (237, 154)(1667) 4 --> (1667) 4:PEGB6, pass, PUGB7
			10'd154 : rdata = 48'b110001110000110000000000000000000000000000001111;
			// PEs: 0 -> 10
			// srcs: (242, 129)(1819) 9 --> (1819) 9:PUNB, pass, PEGB2
			10'd155 : rdata = 48'b110001101111111100000000000000000000000010100000;
			// PEs: 11 -> 56
			// srcs: (245, 176)(1842) 3 --> (1842) 3:PEGB3, pass, PUGB7
			10'd156 : rdata = 48'b110001110000011000000000000000000000000000001111;
			// PEs: 9 -> 56
			// srcs: (246, 191)(2756) -5 --> (2756) -5:PEGB1, pass, PUGB7
			10'd157 : rdata = 48'b110001110000001000000000000000000000000000001111;
			// PEs: 9 -> 24
			// srcs: (247, 192)(2760) 0 --> (2760) 0:PEGB1, pass, PUGB3
			10'd158 : rdata = 48'b110001110000001000000000000000000000000000001011;
			// PEs: 9 -> 56
			// srcs: (248, 193)(2762) -6 --> (2762) -6:PEGB1, pass, PUGB7
			10'd159 : rdata = 48'b110001110000001000000000000000000000000000001111;
			// PEs: 9 -> 0
			// srcs: (249, 201)(2020) 1 --> (2020) 1:PEGB1, pass, PUGB0
			10'd160 : rdata = 48'b110001110000001000000000000000000000000000001000;
			// PEs: 9 -> 32
			// srcs: (250, 221)(2922) 0 --> (2922) 0:PEGB1, pass, PUGB4
			10'd161 : rdata = 48'b110001110000001000000000000000000000000000001100;
			// PEs: 8 -> 10
			// srcs: (251, 130)(1818) 2 --> (1818) 2:NI1, pass, PEGB2
			10'd162 : rdata = 48'b110001010000000100000000000000000000000010100000;
			// PEs: 12 -> 0
			// srcs: (257, 204)(2029) 0 --> (2029) 0:PEGB4, pass, PUGB0
			10'd163 : rdata = 48'b110001110000100000000000000000000000000000001000;
			// PEs: 9 -> 16
			// srcs: (258, 211)(2836) 0 --> (2836) 0:PEGB1, pass, PUNB
			10'd164 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 0 -> 8
			// srcs: (259, 131)(1820) 2 --> (1820) 2:PUNB, pass, NI0
			10'd165 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 9 -> 24
			// srcs: (260, 212)(2838) -8 --> (2838) -8:PEGB1, pass, PUGB3
			10'd166 : rdata = 48'b110001110000001000000000000000000000000000001011;
			// PEs: 9 -> 48
			// srcs: (261, 219)(2917) 0 --> (2917) 0:PEGB1, pass, PUGB6
			10'd167 : rdata = 48'b110001110000001000000000000000000000000000001110;
			// PEs: 15 -> 0
			// srcs: (262, 207)(2038) -2 --> (2038) -2:PENB, pass, PUGB0
			10'd168 : rdata = 48'b110001101111111000000000000000000000000000001000;
			// PEs: 9 -> 40
			// srcs: (263, 220)(2919) 0 --> (2919) 0:PEGB1, pass, PUGB5
			10'd169 : rdata = 48'b110001110000001000000000000000000000000000001101;
			// PEs: 13 -> 56
			// srcs: (264, 238)(3094) -3 --> (3094) -3:PEGB5, pass, PUGB7
			10'd170 : rdata = 48'b110001110000101000000000000000000000000000001111;
			// PEs: 9 -> 48
			// srcs: (271, 222)(2924) -3 --> (2924) -3:PEGB1, pass, PUGB6
			10'd171 : rdata = 48'b110001110000001000000000000000000000000000001110;
			// PEs: 10 -> 40
			// srcs: (272, 224)(2203) 1 --> (2203) 1:PEGB2, pass, PUGB5
			10'd172 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 11 -> 24
			// srcs: (273, 225)(2206) -2 --> (2206) -2:PEGB3, pass, PUGB3
			10'd173 : rdata = 48'b110001110000011000000000000000000000000000001011;
			// PEs: 12 -> 0
			// srcs: (274, 226)(2209) 0 --> (2209) 0:PEGB4, pass, PUGB0
			10'd174 : rdata = 48'b110001110000100000000000000000000000000000001000;
			// PEs: 0 -> 13
			// srcs: (275, 132)(1821) 0 --> (1821) 0:PUNB, pass, PEGB5
			10'd175 : rdata = 48'b110001101111111100000000000000000000000011010000;
			// PEs: 9 -> 16
			// srcs: (276, 230)(3005) 1 --> (3005) 1:PEGB1, pass, PUNB
			10'd176 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 8 -> 13
			// srcs: (284, 133)(1820) 2 --> (1820) 2:NI0, pass, PEGB5
			10'd177 : rdata = 48'b110001010000000000000000000000000000000011010000;
			// PEs: 10 -> 16
			// srcs: (285, 231)(3008) -12 --> (3008) -12:PEGB2, pass, PUNB
			10'd178 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 0 -> 8
			// srcs: (288, 134)(2063) 0 --> (2063) 0:PUNB, pass, NI0
			10'd179 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 11 -> 16
			// srcs: (293, 232)(3010) -4 --> (3010) -4:PEGB3, pass, PUNB
			10'd180 : rdata = 48'b110001110000011000000000000000000000001000000000;
			// PEs: 12 -> 16
			// srcs: (301, 233)(3015) -3 --> (3015) -3:PEGB4, pass, PUNB
			10'd181 : rdata = 48'b110001110000100000000000000000000000001000000000;
			// PEs: 0 -> 9
			// srcs: (304, 135)(2064) -3 --> (2064) -3:PUNB, pass, PENB
			10'd182 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 8 -> 9
			// srcs: (310, 136)(2063) 0 --> (2063) 0:NI0, pass, PENB
			10'd183 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 0 -> 14
			// srcs: (317, 137)(2065) 0 --> (2065) 0:PUNB, pass, PEGB6
			10'd184 : rdata = 48'b110001101111111100000000000000000000000011100000;
			// PEs: 0 -> 9
			// srcs: (324, 138)(2308) 6 --> (2308) 6:PUNB, pass, PENB
			10'd185 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 48 -> 9
			// srcs: (325, 139)(1600) -2 --> (1600) -2:PUGB6, pass, PENB
			10'd186 : rdata = 48'b110001110000110100000000000000000000000100000000;
			// PEs: 48 -> 9
			// srcs: (326, 140)(1603) -3 --> (1603) -3:PUGB6, pass, PENB
			10'd187 : rdata = 48'b110001110000110100000000000000000000000100000000;
			// PEs: 16 -> 8
			// srcs: (327, 146)(2413) -6 --> (2413) -6:PUGB2, pass, NI0
			10'd188 : rdata = 48'b110001110000010100000000000100000000000000000000;
			// PEs: 0 -> 9
			// srcs: (336, 147)(1634) 3 --> (1634) 3:PUNB, pass, PENB
			10'd189 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 8 -> 9
			// srcs: (342, 148)(2413) -6 --> (2413) -6:NI0, pass, PENB
			10'd190 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 24 -> 9
			// srcs: (343, 149)(2431) 7 --> (2431) 7:PUGB3, pass, PENB
			10'd191 : rdata = 48'b110001110000011100000000000000000000000100000000;
			// PEs: 0 -> 9
			// srcs: (344, 153)(2442) -6 --> (2442) -6:PUNB, pass, PENB
			10'd192 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 32 -> 8
			// srcs: (345, 157)(2471) 15 --> (2471) 15:PUGB4, pass, NI0
			10'd193 : rdata = 48'b110001110000100100000000000100000000000000000000;
			// PEs: 9 -> 48
			// srcs: (349, 245)(2414) -3 --> (2414) -3:PEGB1, pass, PUGB6
			10'd194 : rdata = 48'b110001110000001000000000000000000000000000001110;
			// PEs: 9 -> 24
			// srcs: (350, 249)(2432) 7 --> (2432) 7:PEGB1, pass, PUGB3
			10'd195 : rdata = 48'b110001110000001000000000000000000000000000001011;
			// PEs: 9 -> 40
			// srcs: (351, 250)(2443) 0 --> (2443) 0:PEGB1, pass, PUGB5
			10'd196 : rdata = 48'b110001110000001000000000000000000000000000001101;
			// PEs: 11 -> 24
			// srcs: (352, 258)(2602) 13 --> (2602) 13:PEGB3, pass, PUGB3
			10'd197 : rdata = 48'b110001110000011000000000000000000000000000001011;
			// PEs: 10 -> 48
			// srcs: (353, 287)(2385) -3 --> (2385) -3:PEGB2, pass, PUGB6
			10'd198 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 16 -> 9
			// srcs: (367, 158)(1692) 0 --> (1692) 0:PUGB2, pass, PENB
			10'd199 : rdata = 48'b110001110000010100000000000000000000000100000000;
			// PEs: 8 -> 9
			// srcs: (373, 159)(2471) 15 --> (2471) 15:NI0, pass, PENB
			10'd200 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 56 -> 8
			// srcs: (374, 160)(2496) 2 --> (2496) 2:PUGB7, pass, NI0
			10'd201 : rdata = 48'b110001110000111100000000000100000000000000000000;
			// PEs: 32 -> 9
			// srcs: (375, 161)(1719) 6 --> (1719) 6:PUGB4, pass, PENB
			10'd202 : rdata = 48'b110001110000100100000000000000000000000100000000;
			// PEs: 9 -> 0
			// srcs: (380, 251)(2472) 15 --> (2472) 15:PEGB1, pass, PUGB0
			10'd203 : rdata = 48'b110001110000001000000000000000000000000000001000;
			// PEs: 8 -> 9
			// srcs: (381, 162)(2496) 2 --> (2496) 2:NI0, pass, PENB
			10'd204 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 32 -> 9
			// srcs: (382, 165)(1741) 0 --> (1741) 0:PUGB4, pass, PENB
			10'd205 : rdata = 48'b110001110000100100000000000000000000000100000000;
			// PEs: 16 -> 8
			// srcs: (383, 166)(2531) 2 --> (2531) 2:PUGB2, pass, NI0
			10'd206 : rdata = 48'b110001110000010100000000000100000000000000000000;
			// PEs: 40 -> 9
			// srcs: (384, 167)(1753) -4 --> (1753) -4:PUGB5, pass, PENB
			10'd207 : rdata = 48'b110001110000101100000000000000000000000100000000;
			// PEs: 9 -> 0
			// srcs: (389, 256)(2520) -1 --> (2520) -1:PEGB1, pass, PUGB0
			10'd208 : rdata = 48'b110001110000001000000000000000000000000000001000;
			// PEs: 8 -> 9
			// srcs: (390, 168)(2531) 2 --> (2531) 2:NI0, pass, PENB
			10'd209 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 32 -> 8
			// srcs: (391, 170)(2592) 5 --> (2592) 5:PUGB4, pass, NI0
			10'd210 : rdata = 48'b110001110000100100000000000100000000000000000000;
			// PEs: 0 -> 9
			// srcs: (392, 171)(1814) -6 --> (1814) -6:PUNB, pass, PENB
			10'd211 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 9 -> 16
			// srcs: (397, 257)(2532) -2 --> (2532) -2:PEGB1, pass, PUNB
			10'd212 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 8 -> 9
			// srcs: (398, 172)(2592) 5 --> (2592) 5:NI0, pass, PENB
			10'd213 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 0 -> 9
			// srcs: (399, 173)(1817) -1 --> (1817) -1:PUNB, pass, PENB
			10'd214 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 32 -> 9
			// srcs: (400, 178)(2626) 0 --> (2626) 0:PUGB4, pass, PENB
			10'd215 : rdata = 48'b110001110000100100000000000000000000000100000000;
			// PEs: 48 -> 8
			// srcs: (401, 181)(2652) 3 --> (2652) 3:PUGB6, pass, NI0
			10'd216 : rdata = 48'b110001110000110100000000000100000000000000000000;
			// PEs: 16 -> 9
			// srcs: (402, 182)(1873) 2 --> (1873) 2:PUGB2, pass, PENB
			10'd217 : rdata = 48'b110001110000010100000000000000000000000100000000;
			// PEs: 8 -> 9
			// srcs: (413, 183)(2652) 3 --> (2652) 3:NI0, pass, PENB
			10'd218 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 24 -> 9
			// srcs: (414, 184)(1897) -2 --> (1897) -2:PUGB3, pass, PENB
			10'd219 : rdata = 48'b110001110000011100000000000000000000000100000000;
			// PEs: 32 -> 9
			// srcs: (415, 187)(1906) 6 --> (1906) 6:PUGB4, pass, PENB
			10'd220 : rdata = 48'b110001110000100100000000000000000000000100000000;
			// PEs: 0 -> 8
			// srcs: (416, 188)(2751) -4 --> (2751) -4:PUNB, pass, NI0
			10'd221 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 48 -> 9
			// srcs: (417, 189)(1971) -6 --> (1971) -6:PUGB6, pass, PENB
			10'd222 : rdata = 48'b110001110000110100000000000000000000000100000000;
			// PEs: 9 -> 0
			// srcs: (418, 259)(2627) 6 --> (2627) 6:PEGB1, pass, PUGB0
			10'd223 : rdata = 48'b110001110000001000000000000000000000000000001000;
			// PEs: 9 -> 16
			// srcs: (420, 263)(2653) 5 --> (2653) 5:PEGB1, pass, PUNB
			10'd224 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 9 -> 56
			// srcs: (421, 264)(2676) -9 --> (2676) -9:PEGB1, pass, PUGB7
			10'd225 : rdata = 48'b110001110000001000000000000000000000000000001111;
			// PEs: 9 -> 0
			// srcs: (422, 265)(2685) 4 --> (2685) 4:PEGB1, pass, PUGB0
			10'd226 : rdata = 48'b110001110000001000000000000000000000000000001000;
			// PEs: 8 -> 9
			// srcs: (423, 190)(2751) -4 --> (2751) -4:NI0, pass, PENB
			10'd227 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 24 -> 8
			// srcs: (424, 195)(2777) -3 --> (2777) -3:PUGB3, pass, NI0
			10'd228 : rdata = 48'b110001110000011100000000000100000000000000000000;
			// PEs: 0 -> 9
			// srcs: (425, 196)(1998) 0 --> (1998) 0:PUNB, pass, PENB
			10'd229 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 8 -> 9
			// srcs: (431, 197)(2777) -3 --> (2777) -3:NI0, pass, PENB
			10'd230 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 24 -> 8
			// srcs: (432, 198)(2783) -2 --> (2783) -2:PUGB3, pass, NI0
			10'd231 : rdata = 48'b110001110000011100000000000100000000000000000000;
			// PEs: 0 -> 9
			// srcs: (433, 199)(2004) -2 --> (2004) -2:PUNB, pass, PENB
			10'd232 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 9 -> 24
			// srcs: (438, 270)(2778) -3 --> (2778) -3:PEGB1, pass, PUGB3
			10'd233 : rdata = 48'b110001110000001000000000000000000000000000001011;
			// PEs: 8 -> 9
			// srcs: (439, 200)(2783) -2 --> (2783) -2:NI0, pass, PENB
			10'd234 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 0 -> 8
			// srcs: (440, 208)(2827) 1 --> (2827) 1:PUNB, pass, NI0
			10'd235 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 16 -> 9
			// srcs: (441, 209)(2050) 0 --> (2050) 0:PUGB2, pass, PENB
			10'd236 : rdata = 48'b110001110000010100000000000000000000000100000000;
			// PEs: 9 -> 56
			// srcs: (446, 271)(2784) -4 --> (2784) -4:PEGB1, pass, PUGB7
			10'd237 : rdata = 48'b110001110000001000000000000000000000000000001111;
			// PEs: 8 -> 9
			// srcs: (447, 210)(2827) 1 --> (2827) 1:NI0, pass, PENB
			10'd238 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 56 -> 8
			// srcs: (448, 213)(2901) 6 --> (2901) 6:PUGB7, pass, NI0
			10'd239 : rdata = 48'b110001110000111100000000000100000000000000000000;
			// PEs: 40 -> 9
			// srcs: (449, 214)(2124) -3 --> (2124) -3:PUGB5, pass, PENB
			10'd240 : rdata = 48'b110001110000101100000000000000000000000100000000;
			// PEs: 9 -> 56
			// srcs: (454, 272)(2828) 1 --> (2828) 1:PEGB1, pass, PUGB7
			10'd241 : rdata = 48'b110001110000001000000000000000000000000000001111;
			// PEs: 8 -> 9
			// srcs: (455, 215)(2901) 6 --> (2901) 6:NI0, pass, PENB
			10'd242 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 0 -> 8
			// srcs: (456, 216)(2907) 2 --> (2907) 2:PUNB, pass, NI0
			10'd243 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 40 -> 9
			// srcs: (457, 217)(2130) -4 --> (2130) -4:PUGB5, pass, PENB
			10'd244 : rdata = 48'b110001110000101100000000000000000000000100000000;
			// PEs: 0 -> 11
			// srcs: (458, 227)(2994) -1 --> (2994) -1:PUNB, pass, PEGB3
			10'd245 : rdata = 48'b110001101111111100000000000000000000000010110000;
			// PEs: 8 -> 9
			// srcs: (463, 218)(2907) 2 --> (2907) 2:NI0, pass, PENB
			10'd246 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 56 -> 9
			// srcs: (464, 223)(2978) -4 --> (2978) -4:PUGB7, pass, PENB
			10'd247 : rdata = 48'b110001110000111100000000000000000000000100000000;
			// PEs: 9 -> 16
			// srcs: (470, 275)(2908) -2 --> (2908) -2:PEGB1, pass, PUNB
			10'd248 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 9 -> 40
			// srcs: (471, 279)(2979) -7 --> (2979) -7:PEGB1, pass, PUGB5
			10'd249 : rdata = 48'b110001110000001000000000000000000000000000001101;
			// PEs: 0 -> 9
			// srcs: (494, 228)(2997) 1 --> (2997) 1:PUNB, pass, PENB
			10'd250 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 0 -> 9
			// srcs: (513, 229)(2999) 0 --> (2999) 0:PUNB, pass, PENB
			10'd251 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 56 -> 8
			// srcs: (514, 234)(3071) -1 --> (3071) -1:PUGB7, pass, NI0
			10'd252 : rdata = 48'b110001110000111100000000000100000000000000000000;
			// PEs: 40 -> 9
			// srcs: (515, 235)(2295) 1 --> (2295) 1:PUGB5, pass, PENB
			10'd253 : rdata = 48'b110001110000101100000000000000000000000100000000;
			// PEs: 8 -> 9
			// srcs: (521, 236)(3071) -1 --> (3071) -1:NI0, pass, PENB
			10'd254 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 40 -> 9
			// srcs: (522, 237)(2314) 4 --> (2314) 4:PUGB5, pass, PENB
			10'd255 : rdata = 48'b110001110000101100000000000000000000000100000000;
			// PEs: 24 -> 8
			// srcs: (523, 239)(3114) 4 --> (3114) 4:PUGB3, pass, NI0
			10'd256 : rdata = 48'b110001110000011100000000000100000000000000000000;
			// PEs: 9 -> 32
			// srcs: (528, 281)(3072) 0 --> (3072) 0:PEGB1, pass, PUGB4
			10'd257 : rdata = 48'b110001110000001000000000000000000000000000001100;
			// PEs: 56 -> 9
			// srcs: (532, 240)(2338) 0 --> (2338) 0:PUGB7, pass, PENB
			10'd258 : rdata = 48'b110001110000111100000000000000000000000100000000;
			// PEs: 8 -> 9
			// srcs: (538, 241)(3114) 4 --> (3114) 4:NI0, pass, PENB
			10'd259 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 40 -> 8
			// srcs: (539, 242)(3128) 8 --> (3128) 8:PUGB5, pass, NI0
			10'd260 : rdata = 48'b110001110000101100000000000100000000000000000000;
			// PEs: 9 -> 0
			// srcs: (545, 282)(3115) 4 --> (3115) 4:PEGB1, pass, PUGB0
			10'd261 : rdata = 48'b110001110000001000000000000000000000000000001000;
			// PEs: 56 -> 9
			// srcs: (548, 243)(2353) 1 --> (2353) 1:PUGB7, pass, PENB
			10'd262 : rdata = 48'b110001110000111100000000000000000000000100000000;
			// PEs: 8 -> 9
			// srcs: (554, 244)(3128) 8 --> (3128) 8:NI0, pass, PENB
			10'd263 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 0 -> 8
			// srcs: (555, 246)(2423) -3 --> (2423) -3:PUNB, pass, NI0
			10'd264 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 16 -> 9
			// srcs: (556, 247)(2425) -5 --> (2425) -5:PUGB2, pass, PENB
			10'd265 : rdata = 48'b110001110000010100000000000000000000000100000000;
			// PEs: 9 -> 24
			// srcs: (561, 286)(3129) 9 --> (3129) 9:PEGB1, pass, PUGB3
			10'd266 : rdata = 48'b110001110000001000000000000000000000000000001011;
			// PEs: 8 -> 9
			// srcs: (562, 248)(2423) -3 --> (2423) -3:NI0, pass, PENB
			10'd267 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 0 -> 8
			// srcs: (563, 252)(2484) -3 --> (2484) -3:PUNB, pass, NI0
			10'd268 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 16 -> 9
			// srcs: (564, 253)(2486) 17 --> (2486) 17:PUGB2, pass, PENB
			10'd269 : rdata = 48'b110001110000010100000000000000000000000100000000;
			// PEs: 9 -> 56
			// srcs: (569, 288)(2426) -8 --> (2426) -8:PEGB1, pass, PUGB7
			10'd270 : rdata = 48'b110001110000001000000000000000000000000000001111;
			// PEs: 8 -> 9
			// srcs: (570, 254)(2484) -3 --> (2484) -3:NI0, pass, PENB
			10'd271 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 0 -> 9
			// srcs: (571, 255)(2495) 5 --> (2495) 5:PUNB, pass, PENB
			10'd272 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 0 -> 8
			// srcs: (572, 260)(2630) 3 --> (2630) 3:PUNB, pass, NI0
			10'd273 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 32 -> 9
			// srcs: (573, 261)(2632) 0 --> (2632) 0:PUGB4, pass, PENB
			10'd274 : rdata = 48'b110001110000100100000000000000000000000100000000;
			// PEs: 9 -> 40
			// srcs: (577, 292)(2487) 14 --> (2487) 14:PEGB1, pass, PUGB5
			10'd275 : rdata = 48'b110001110000001000000000000000000000000000001101;
			// PEs: 9 -> 0
			// srcs: (578, 293)(2498) 13 --> (2498) 13:PEGB1, pass, PUGB0
			10'd276 : rdata = 48'b110001110000001000000000000000000000000000001000;
			// PEs: 8 -> 9
			// srcs: (579, 262)(2630) 3 --> (2630) 3:NI0, pass, PENB
			10'd277 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 0 -> 9
			// srcs: (580, 266)(2750) -1 --> (2750) -1:PUNB, pass, PENB
			10'd278 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 24 -> 8
			// srcs: (594, 267)(2761) 0 --> (2761) 0:PUGB3, pass, NI0
			10'd279 : rdata = 48'b110001110000011100000000000100000000000000000000;
			// PEs: 56 -> 9
			// srcs: (595, 268)(2763) -4 --> (2763) -4:PUGB7, pass, PENB
			10'd280 : rdata = 48'b110001110000111100000000000000000000000100000000;
			// PEs: 8 -> 9
			// srcs: (601, 269)(2761) 0 --> (2761) 0:NI0, pass, PENB
			10'd281 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 9 -> 16
			// srcs: (608, 297)(2764) -4 --> (2764) -4:PEGB1, pass, PUNB
			10'd282 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 24 -> 9
			// srcs: (627, 273)(2849) -1 --> (2849) -1:PUGB3, pass, PENB
			10'd283 : rdata = 48'b110001110000011100000000000000000000000100000000;
			// PEs: 56 -> 9
			// srcs: (628, 274)(2900) 13 --> (2900) 13:PUGB7, pass, PENB
			10'd284 : rdata = 48'b110001110000111100000000000000000000000100000000;
			// PEs: 32 -> 8
			// srcs: (629, 276)(2956) 11 --> (2956) 11:PUGB4, pass, NI0
			10'd285 : rdata = 48'b110001110000100100000000000100000000000000000000;
			// PEs: 48 -> 9
			// srcs: (630, 277)(2958) 0 --> (2958) 0:PUGB6, pass, PENB
			10'd286 : rdata = 48'b110001110000110100000000000000000000000100000000;
			// PEs: 9 -> 0
			// srcs: (635, 298)(2850) -4 --> (2850) -4:PEGB1, pass, PUGB0
			10'd287 : rdata = 48'b110001110000001000000000000000000000000000001000;
			// PEs: 8 -> 9
			// srcs: (636, 278)(2956) 11 --> (2956) 11:NI0, pass, PENB
			10'd288 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 0 -> 9
			// srcs: (637, 280)(2993) -2 --> (2993) -2:PUNB, pass, PENB
			10'd289 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 9 -> 16
			// srcs: (643, 303)(2959) 11 --> (2959) 11:PEGB1, pass, PUNB
			10'd290 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 40 -> 8
			// srcs: (717, 283)(3118) -5 --> (3118) -5:PUGB5, pass, NI0
			10'd291 : rdata = 48'b110001110000101100000000000100000000000000000000;
			// PEs: 0 -> 9
			// srcs: (718, 284)(3120) -4 --> (3120) -4:PUNB, pass, PENB
			10'd292 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 8 -> 9
			// srcs: (724, 285)(3118) -5 --> (3118) -5:NI0, pass, PENB
			10'd293 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 40 -> 8
			// srcs: (734, 289)(2444) 2 --> (2444) 2:PUGB5, pass, NI0
			10'd294 : rdata = 48'b110001110000101100000000000100000000000000000000;
			// PEs: 56 -> 9
			// srcs: (735, 290)(2449) 6 --> (2449) 6:PUGB7, pass, PENB
			10'd295 : rdata = 48'b110001110000111100000000000000000000000100000000;
			// PEs: 8 -> 9
			// srcs: (741, 291)(2444) 2 --> (2444) 2:NI0, pass, PENB
			10'd296 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 0 -> 9
			// srcs: (742, 294)(2591) 14 --> (2591) 14:PUNB, pass, PENB
			10'd297 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 9 -> 48
			// srcs: (748, 306)(2450) 8 --> (2450) 8:PEGB1, pass, PUGB6
			10'd298 : rdata = 48'b110001110000001000000000000000000000000000001110;
			// PEs: 0 -> 9
			// srcs: (967, 295)(2628) 16 --> (2628) 16:PUNB, pass, PENB
			10'd299 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 9 -> 32
			// srcs: (975, 308)(2634) 19 --> (2634) 19:PEGB1, pass, PUGB4
			10'd300 : rdata = 48'b110001110000001000000000000000000000000000001100;
			// PEs: 0 -> 9
			// srcs: (985, 296)(2758) -7 --> (2758) -7:PUNB, pass, PENB
			10'd301 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 56 -> 9
			// srcs: (986, 299)(2898) 11 --> (2898) 11:PUGB7, pass, PENB
			10'd302 : rdata = 48'b110001110000111100000000000000000000000100000000;
			// PEs: 9 -> 16
			// srcs: (992, 309)(2759) -18 --> (2759) -18:PEGB1, pass, PUNB
			10'd303 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 9 -> 16
			// srcs: (993, 313)(2904) 27 --> (2904) 27:PEGB1, pass, PUNB
			10'd304 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 32 -> 8
			// srcs: (1118, 300)(2948) 10 --> (2948) 10:PUGB4, pass, NI0
			10'd305 : rdata = 48'b110001110000100100000000000100000000000000000000;
			// PEs: 0 -> 9
			// srcs: (1119, 301)(2953) -4 --> (2953) -4:PUNB, pass, PENB
			10'd306 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 8 -> 9
			// srcs: (1125, 302)(2948) 10 --> (2948) 10:NI0, pass, PENB
			10'd307 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 0 -> 9
			// srcs: (1126, 304)(3098) -1 --> (3098) -1:PUNB, pass, PENB
			10'd308 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 0 -> 9
			// srcs: (1127, 305)(3116) -2 --> (3116) -2:PUNB, pass, PENB
			10'd309 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 9 -> 16
			// srcs: (1132, 314)(2954) 6 --> (2954) 6:PEGB1, pass, PUNB
			10'd310 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 10 -> 16
			// srcs: (1133, 315)(3002) -9 --> (3002) -9:PEGB2, pass, PUNB
			10'd311 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 9 -> 0
			// srcs: (1134, 316)(3099) 15 --> (3099) 15:PEGB1, pass, PUGB0
			10'd312 : rdata = 48'b110001110000001000000000000000000000000000001000;
			// PEs: 0 -> 9
			// srcs: (1173, 307)(2586) -24 --> (2586) -24:PUNB, pass, PENB
			10'd313 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 24 -> 8
			// srcs: (1174, 310)(2807) 6 --> (2807) 6:PUGB3, pass, NI0
			10'd314 : rdata = 48'b110001110000011100000000000100000000000000000000;
			// PEs: 48 -> 9
			// srcs: (1397, 311)(2818) -3 --> (2818) -3:PUGB6, pass, PENB
			10'd315 : rdata = 48'b110001110000110100000000000000000000000100000000;
			// PEs: 8 -> 9
			// srcs: (1404, 312)(2807) 6 --> (2807) 6:NI0, pass, PENB
			10'd316 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 32 -> 9
			// srcs: (1405, 317)(3133) 11 --> (3133) 11:PUGB4, pass, PENB
			10'd317 : rdata = 48'b110001110000100100000000000000000000000100000000;
			// PEs: 56 -> 9
			// srcs: (1406, 318)(2575) 19 --> (2575) 19:PUGB7, pass, PENB
			10'd318 : rdata = 48'b110001110000111100000000000000000000000100000000;
			// PEs: 16 -> 8
			// srcs: (1407, 319)(2771) -20 --> (2771) -20:PUGB2, pass, NI0
			10'd319 : rdata = 48'b110001110000010100000000000100000000000000000000;
			// PEs: 32 -> 9
			// srcs: (1408, 320)(2794) -1 --> (2794) -1:PUGB4, pass, PENB
			10'd320 : rdata = 48'b110001110000100100000000000000000000000100000000;
			// PEs: 9 -> 24
			// srcs: (1411, 322)(2819) 3 --> (2819) 3:PEGB1, pass, PUGB3
			10'd321 : rdata = 48'b110001110000001000000000000000000000000000001011;
			// PEs: 9 -> 48
			// srcs: (1413, 324)(2599) 4 --> (2599) 4:PEGB1, pass, PUGB6
			10'd322 : rdata = 48'b110001110000001000000000000000000000000000001110;
			// PEs: 8 -> 9
			// srcs: (1414, 321)(2771) -20 --> (2771) -20:NI0, pass, PENB
			10'd323 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 0 -> 9
			// srcs: (1415, 323)(3111) 3 --> (3111) 3:PUNB, pass, PENB
			10'd324 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 9 -> 16
			// srcs: (1421, 325)(2795) -21 --> (2795) -21:PEGB1, pass, PUNB
			10'd325 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 0 -> 9
			// srcs: (1434, 326)(3087) -28 --> (3087) -28:PUNB, pass, PENB
			10'd326 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 9 -> 40
			// srcs: (1442, 327)(3136) -25 --> (3136) -25:PEGB1, pass, PUGB5
			10'd327 : rdata = 48'b110001110000001000000000000000000000000000001101;
			// PEs: 0 -> 8
			// srcs: (1456, 328)(2747) 88 --> (2747) 88:PUNB, pass, NI0
			10'd328 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 48 -> 9
			// srcs: (1485, 329)(3138) -39 --> (3138) -39:PUGB6, pass, PENB
			10'd329 : rdata = 48'b110001110000110100000000000000000000000100000000;
			// PEs: 8 -> 9
			// srcs: (1492, 330)(2747) 88 --> (2747) 88:NI0, pass, PENB
			10'd330 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 10 -> 0
			// srcs: (1502, 331)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd331 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 0
			// srcs: (1506, 332)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd332 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 0
			// srcs: (1507, 333)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd333 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 0
			// srcs: (1508, 334)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd334 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 0
			// srcs: (1509, 335)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd335 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 0
			// srcs: (1510, 336)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd336 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 40
			// srcs: (1511, 337)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd337 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 0
			// srcs: (1512, 338)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd338 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 40
			// srcs: (1514, 339)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd339 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 48
			// srcs: (1516, 340)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd340 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 48
			// srcs: (1519, 341)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd341 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 48
			// srcs: (1522, 342)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd342 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 16
			// srcs: (1523, 343)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd343 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 16
			// srcs: (1524, 344)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd344 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 48
			// srcs: (1525, 345)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd345 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 16
			// srcs: (1526, 346)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd346 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 16
			// srcs: (1527, 347)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd347 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 48
			// srcs: (1528, 348)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd348 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 16
			// srcs: (1529, 349)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd349 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 16
			// srcs: (1530, 350)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd350 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 48
			// srcs: (1531, 351)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd351 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 16
			// srcs: (1532, 352)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd352 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 24
			// srcs: (1533, 353)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd353 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 48
			// srcs: (1534, 354)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd354 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 24
			// srcs: (1535, 355)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd355 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 24
			// srcs: (1536, 356)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd356 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 56
			// srcs: (1537, 357)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd357 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 24
			// srcs: (1538, 358)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd358 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 24
			// srcs: (1539, 359)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd359 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 56
			// srcs: (1540, 360)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd360 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 24
			// srcs: (1541, 361)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd361 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 24
			// srcs: (1542, 362)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd362 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 56
			// srcs: (1543, 363)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd363 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 32
			// srcs: (1544, 364)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd364 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 32
			// srcs: (1545, 365)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd365 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 56
			// srcs: (1546, 366)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd366 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 32
			// srcs: (1547, 367)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd367 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 32
			// srcs: (1548, 368)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd368 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 56
			// srcs: (1549, 369)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd369 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 32
			// srcs: (1550, 370)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd370 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 32
			// srcs: (1551, 371)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd371 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 56
			// srcs: (1552, 372)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd372 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 32
			// srcs: (1553, 373)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd373 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 40
			// srcs: (1554, 374)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd374 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 40
			// srcs: (1555, 375)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd375 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 40
			// srcs: (1556, 376)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd376 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 40
			// srcs: (1557, 377)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd377 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 40
			// srcs: (1558, 378)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd378 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 56
			// srcs: (1559, 379)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd379 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 40
			// srcs: (1560, 380)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd380 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 40
			// srcs: (1561, 381)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd381 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 0
			// srcs: (1562, 382)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd382 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 48
			// srcs: (1563, 383)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd383 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 48
			// srcs: (1564, 384)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd384 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 0
			// srcs: (1565, 385)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd385 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 48
			// srcs: (1566, 386)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd386 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 48
			// srcs: (1567, 387)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd387 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 0
			// srcs: (1568, 388)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd388 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 48
			// srcs: (1569, 389)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd389 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 48
			// srcs: (1570, 390)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd390 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 0
			// srcs: (1571, 391)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd391 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 48
			// srcs: (1572, 392)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd392 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 56
			// srcs: (1573, 393)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd393 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 0
			// srcs: (1574, 394)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd394 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 56
			// srcs: (1575, 395)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd395 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 56
			// srcs: (1576, 396)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd396 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 0
			// srcs: (1577, 397)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd397 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 56
			// srcs: (1578, 398)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd398 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 56
			// srcs: (1579, 399)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd399 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 0
			// srcs: (1580, 400)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd400 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 56
			// srcs: (1581, 401)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd401 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 56
			// srcs: (1582, 402)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd402 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 0
			// srcs: (1584, 403)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd403 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 0
			// srcs: (1585, 404)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd404 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 0
			// srcs: (1587, 405)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd405 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 0
			// srcs: (1588, 406)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd406 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 0
			// srcs: (1590, 407)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd407 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 0
			// srcs: (1591, 408)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd408 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 0
			// srcs: (1593, 409)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd409 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 16
			// srcs: (1604, 410)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd410 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 16
			// srcs: (1605, 411)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd411 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 16
			// srcs: (1606, 412)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd412 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 16
			// srcs: (1607, 413)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd413 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 16
			// srcs: (1608, 414)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd414 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 16
			// srcs: (1609, 415)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd415 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 16
			// srcs: (1610, 416)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd416 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 16
			// srcs: (1611, 417)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd417 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 16
			// srcs: (1612, 418)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd418 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 24
			// srcs: (1613, 419)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd419 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 16
			// srcs: (1614, 420)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd420 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 24
			// srcs: (1615, 421)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd421 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 24
			// srcs: (1616, 422)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd422 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 16
			// srcs: (1617, 423)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd423 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 24
			// srcs: (1618, 424)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd424 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 24
			// srcs: (1619, 425)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd425 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 16
			// srcs: (1620, 426)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd426 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 24
			// srcs: (1621, 427)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd427 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 24
			// srcs: (1622, 428)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd428 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 16
			// srcs: (1623, 429)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd429 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 32
			// srcs: (1624, 430)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd430 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 32
			// srcs: (1625, 431)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd431 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 16
			// srcs: (1626, 432)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd432 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 32
			// srcs: (1627, 433)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd433 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 32
			// srcs: (1628, 434)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd434 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 24
			// srcs: (1629, 435)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd435 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 32
			// srcs: (1630, 436)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd436 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 32
			// srcs: (1631, 437)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd437 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 24
			// srcs: (1632, 438)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd438 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 32
			// srcs: (1633, 439)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd439 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 40
			// srcs: (1634, 440)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd440 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 24
			// srcs: (1635, 441)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd441 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 40
			// srcs: (1636, 442)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd442 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 40
			// srcs: (1637, 443)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd443 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 24
			// srcs: (1638, 444)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd444 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 40
			// srcs: (1639, 445)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd445 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 40
			// srcs: (1640, 446)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd446 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 24
			// srcs: (1641, 447)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd447 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 40
			// srcs: (1642, 448)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd448 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 40
			// srcs: (1643, 449)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd449 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 24
			// srcs: (1644, 450)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd450 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 48
			// srcs: (1645, 451)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd451 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 48
			// srcs: (1646, 452)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd452 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 24
			// srcs: (1647, 453)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd453 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 48
			// srcs: (1648, 454)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd454 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 48
			// srcs: (1649, 455)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd455 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 32
			// srcs: (1650, 456)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd456 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 48
			// srcs: (1651, 457)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd457 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 48
			// srcs: (1652, 458)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd458 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 48
			// srcs: (1653, 459)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd459 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 56
			// srcs: (1654, 460)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd460 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 56
			// srcs: (1655, 461)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd461 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 56
			// srcs: (1656, 462)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd462 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 32
			// srcs: (1657, 463)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd463 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 56
			// srcs: (1658, 464)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd464 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 56
			// srcs: (1659, 465)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd465 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 32
			// srcs: (1660, 466)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd466 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 56
			// srcs: (1661, 467)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd467 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 56
			// srcs: (1662, 468)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd468 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 32
			// srcs: (1663, 469)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd469 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 0
			// srcs: (1664, 470)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd470 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 0
			// srcs: (1665, 471)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd471 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 32
			// srcs: (1666, 472)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd472 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 0
			// srcs: (1667, 473)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd473 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 0
			// srcs: (1668, 474)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd474 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 32
			// srcs: (1669, 475)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd475 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 0
			// srcs: (1670, 476)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd476 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 0
			// srcs: (1671, 477)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd477 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 32
			// srcs: (1672, 478)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd478 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 0
			// srcs: (1673, 479)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd479 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 40
			// srcs: (1675, 480)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd480 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 40
			// srcs: (1678, 481)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd481 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 40
			// srcs: (1681, 482)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd482 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 40
			// srcs: (1684, 483)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd483 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 16
			// srcs: (1685, 484)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd484 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 16
			// srcs: (1686, 485)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd485 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 40
			// srcs: (1687, 486)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd486 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 16
			// srcs: (1688, 487)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd487 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 16
			// srcs: (1689, 488)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd488 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 40
			// srcs: (1690, 489)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd489 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 16
			// srcs: (1691, 490)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd490 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 16
			// srcs: (1692, 491)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd491 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 40
			// srcs: (1693, 492)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd492 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 16
			// srcs: (1694, 493)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd493 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 24
			// srcs: (1695, 494)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd494 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 48
			// srcs: (1696, 495)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd495 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 24
			// srcs: (1697, 496)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd496 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 24
			// srcs: (1698, 497)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd497 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 48
			// srcs: (1699, 498)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd498 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 24
			// srcs: (1700, 499)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd499 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 24
			// srcs: (1701, 500)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd500 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 24
			// srcs: (1702, 501)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd501 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 24
			// srcs: (1703, 502)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd502 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 32
			// srcs: (1704, 503)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd503 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 32
			// srcs: (1705, 504)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd504 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 48
			// srcs: (1706, 505)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd505 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 32
			// srcs: (1707, 506)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd506 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 32
			// srcs: (1708, 507)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd507 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 48
			// srcs: (1709, 508)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd508 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 32
			// srcs: (1710, 509)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd509 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 32
			// srcs: (1711, 510)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd510 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 48
			// srcs: (1712, 511)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd511 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 32
			// srcs: (1713, 512)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd512 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 40
			// srcs: (1714, 513)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd513 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 48
			// srcs: (1715, 514)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd514 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 40
			// srcs: (1716, 515)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd515 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 40
			// srcs: (1717, 516)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd516 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 48
			// srcs: (1718, 517)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd517 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 40
			// srcs: (1719, 518)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd518 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 40
			// srcs: (1720, 519)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd519 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 56
			// srcs: (1721, 520)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd520 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 40
			// srcs: (1722, 521)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd521 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 40
			// srcs: (1723, 522)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd522 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 56
			// srcs: (1724, 523)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd523 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 48
			// srcs: (1725, 524)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd524 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 48
			// srcs: (1726, 525)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd525 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 56
			// srcs: (1727, 526)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd526 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 48
			// srcs: (1728, 527)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd527 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 48
			// srcs: (1729, 528)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd528 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 56
			// srcs: (1730, 529)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd529 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 48
			// srcs: (1731, 530)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd530 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 48
			// srcs: (1732, 531)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd531 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 56
			// srcs: (1733, 532)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd532 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 48
			// srcs: (1734, 533)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd533 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 56
			// srcs: (1735, 534)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd534 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 56
			// srcs: (1736, 535)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd535 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 56
			// srcs: (1737, 536)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd536 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 56
			// srcs: (1738, 537)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd537 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 56
			// srcs: (1739, 538)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd538 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 56
			// srcs: (1740, 539)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd539 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 56
			// srcs: (1741, 540)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd540 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 0
			// srcs: (1742, 541)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd541 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 56
			// srcs: (1743, 542)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd542 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 56
			// srcs: (1744, 543)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd543 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 0
			// srcs: (1745, 544)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd544 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 0
			// srcs: (1746, 545)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd545 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 0
			// srcs: (1747, 546)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd546 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 0
			// srcs: (1748, 547)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd547 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 0
			// srcs: (1749, 548)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd548 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 0
			// srcs: (1750, 549)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd549 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 0
			// srcs: (1751, 550)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd550 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 0
			// srcs: (1752, 551)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd551 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 0
			// srcs: (1753, 552)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd552 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 0
			// srcs: (1755, 553)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd553 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 0
			// srcs: (1758, 554)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd554 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 0
			// srcs: (1761, 555)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd555 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 0
			// srcs: (1764, 556)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd556 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 16
			// srcs: (1765, 557)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd557 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 16
			// srcs: (1766, 558)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd558 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 16
			// srcs: (1768, 559)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd559 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 16
			// srcs: (1769, 560)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd560 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 16
			// srcs: (1771, 561)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd561 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 16
			// srcs: (1772, 562)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd562 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 16
			// srcs: (1774, 563)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd563 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 24
			// srcs: (1775, 564)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd564 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 24
			// srcs: (1777, 565)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd565 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 24
			// srcs: (1778, 566)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd566 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 24
			// srcs: (1780, 567)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd567 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 24
			// srcs: (1781, 568)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd568 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 24
			// srcs: (1783, 569)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd569 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 24
			// srcs: (1784, 570)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd570 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 32
			// srcs: (1786, 571)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd571 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 32
			// srcs: (1787, 572)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd572 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 16
			// srcs: (1788, 573)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd573 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 32
			// srcs: (1789, 574)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd574 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 32
			// srcs: (1790, 575)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd575 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 16
			// srcs: (1791, 576)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd576 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 32
			// srcs: (1792, 577)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd577 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 32
			// srcs: (1793, 578)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd578 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 16
			// srcs: (1794, 579)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd579 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 32
			// srcs: (1795, 580)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd580 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 40
			// srcs: (1796, 581)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd581 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 16
			// srcs: (1797, 582)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd582 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 40
			// srcs: (1798, 583)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd583 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 40
			// srcs: (1799, 584)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd584 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 40
			// srcs: (1800, 585)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd585 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 40
			// srcs: (1801, 586)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd586 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 40
			// srcs: (1802, 587)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd587 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 40
			// srcs: (1803, 588)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd588 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 16
			// srcs: (1804, 589)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd589 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 48
			// srcs: (1805, 590)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd590 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 48
			// srcs: (1806, 591)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd591 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 16
			// srcs: (1807, 592)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd592 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 48
			// srcs: (1808, 593)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd593 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 48
			// srcs: (1809, 594)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd594 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 16
			// srcs: (1810, 595)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd595 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 48
			// srcs: (1811, 596)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd596 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 48
			// srcs: (1812, 597)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd597 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 24
			// srcs: (1813, 598)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd598 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 48
			// srcs: (1814, 599)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd599 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 56
			// srcs: (1815, 600)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd600 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 24
			// srcs: (1816, 601)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd601 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 56
			// srcs: (1817, 602)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd602 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 56
			// srcs: (1818, 603)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd603 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 24
			// srcs: (1819, 604)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd604 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 56
			// srcs: (1820, 605)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd605 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 56
			// srcs: (1821, 606)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd606 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 24
			// srcs: (1822, 607)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd607 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 56
			// srcs: (1823, 608)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd608 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 56
			// srcs: (1824, 609)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd609 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 24
			// srcs: (1825, 610)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd610 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 0
			// srcs: (1826, 611)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd611 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 0
			// srcs: (1827, 612)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd612 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 24
			// srcs: (1828, 613)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd613 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 0
			// srcs: (1829, 614)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd614 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 0
			// srcs: (1830, 615)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd615 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 24
			// srcs: (1831, 616)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd616 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 0
			// srcs: (1832, 617)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd617 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 0
			// srcs: (1833, 618)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd618 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 32
			// srcs: (1834, 619)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd619 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 0
			// srcs: (1835, 620)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd620 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 32
			// srcs: (1837, 621)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd621 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 32
			// srcs: (1840, 622)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd622 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 32
			// srcs: (1843, 623)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd623 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 32
			// srcs: (1846, 624)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd624 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 16
			// srcs: (1847, 625)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd625 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 16
			// srcs: (1848, 626)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd626 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 16
			// srcs: (1849, 627)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd627 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 16
			// srcs: (1850, 628)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd628 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 16
			// srcs: (1851, 629)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd629 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 16
			// srcs: (1852, 630)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd630 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 32
			// srcs: (1853, 631)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd631 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 16
			// srcs: (1854, 632)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd632 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 24
			// srcs: (1855, 633)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd633 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 32
			// srcs: (1856, 634)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd634 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 24
			// srcs: (1857, 635)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd635 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 24
			// srcs: (1858, 636)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd636 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 40
			// srcs: (1859, 637)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd637 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 24
			// srcs: (1860, 638)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd638 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 24
			// srcs: (1861, 639)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd639 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 40
			// srcs: (1862, 640)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd640 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 24
			// srcs: (1863, 641)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd641 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 24
			// srcs: (1864, 642)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd642 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 40
			// srcs: (1865, 643)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd643 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 32
			// srcs: (1866, 644)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd644 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 32
			// srcs: (1867, 645)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd645 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 40
			// srcs: (1868, 646)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd646 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 32
			// srcs: (1869, 647)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd647 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 32
			// srcs: (1870, 648)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd648 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 40
			// srcs: (1871, 649)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd649 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 32
			// srcs: (1872, 650)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd650 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 32
			// srcs: (1873, 651)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd651 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 40
			// srcs: (1874, 652)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd652 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 32
			// srcs: (1875, 653)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd653 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 40
			// srcs: (1876, 654)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd654 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 40
			// srcs: (1877, 655)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd655 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 40
			// srcs: (1878, 656)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd656 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 40
			// srcs: (1879, 657)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd657 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 48
			// srcs: (1880, 658)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd658 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 40
			// srcs: (1881, 659)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd659 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 40
			// srcs: (1882, 660)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd660 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 48
			// srcs: (1883, 661)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd661 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 40
			// srcs: (1884, 662)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd662 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 40
			// srcs: (1885, 663)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd663 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 48
			// srcs: (1886, 664)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd664 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 48
			// srcs: (1887, 665)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd665 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 48
			// srcs: (1888, 666)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd666 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 48
			// srcs: (1889, 667)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd667 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 48
			// srcs: (1890, 668)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd668 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 48
			// srcs: (1891, 669)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd669 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 48
			// srcs: (1892, 670)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd670 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 48
			// srcs: (1893, 671)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd671 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 48
			// srcs: (1894, 672)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd672 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 48
			// srcs: (1895, 673)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd673 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 48
			// srcs: (1896, 674)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd674 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 56
			// srcs: (1897, 675)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd675 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 56
			// srcs: (1898, 676)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd676 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 56
			// srcs: (1899, 677)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd677 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 56
			// srcs: (1900, 678)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd678 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 56
			// srcs: (1901, 679)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd679 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 48
			// srcs: (1902, 680)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd680 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 56
			// srcs: (1903, 681)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd681 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 56
			// srcs: (1904, 682)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd682 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 56
			// srcs: (1905, 683)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd683 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 0
			// srcs: (1906, 684)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd684 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 0
			// srcs: (1907, 685)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd685 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 56
			// srcs: (1908, 686)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd686 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 0
			// srcs: (1909, 687)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd687 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 0
			// srcs: (1910, 688)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd688 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 56
			// srcs: (1911, 689)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd689 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 0
			// srcs: (1912, 690)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd690 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 0
			// srcs: (1913, 691)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd691 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 56
			// srcs: (1914, 692)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd692 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 0
			// srcs: (1915, 693)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd693 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 56
			// srcs: (1917, 694)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd694 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 56
			// srcs: (1920, 695)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd695 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 56
			// srcs: (1923, 696)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd696 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 0
			// srcs: (1926, 697)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd697 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 16
			// srcs: (1927, 698)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd698 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 16
			// srcs: (1928, 699)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd699 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 0
			// srcs: (1929, 700)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd700 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 16
			// srcs: (1930, 701)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd701 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 16
			// srcs: (1931, 702)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd702 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 0
			// srcs: (1932, 703)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd703 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 16
			// srcs: (1933, 704)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd704 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 16
			// srcs: (1934, 705)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd705 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 0
			// srcs: (1935, 706)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd706 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 16
			// srcs: (1936, 707)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd707 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 24
			// srcs: (1937, 708)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd708 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 0
			// srcs: (1938, 709)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd709 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 24
			// srcs: (1939, 710)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd710 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 24
			// srcs: (1940, 711)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd711 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 0
			// srcs: (1941, 712)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd712 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 24
			// srcs: (1942, 713)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd713 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 24
			// srcs: (1943, 714)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd714 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 0
			// srcs: (1944, 715)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd715 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 24
			// srcs: (1945, 716)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd716 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 24
			// srcs: (1946, 717)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd717 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 32
			// srcs: (1947, 718)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd718 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 32
			// srcs: (1948, 719)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd719 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 32
			// srcs: (1949, 720)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd720 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 32
			// srcs: (1950, 721)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd721 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 32
			// srcs: (1952, 722)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd722 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 32
			// srcs: (1953, 723)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd723 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 32
			// srcs: (1955, 724)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd724 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 40
			// srcs: (1956, 725)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd725 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 40
			// srcs: (1958, 726)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd726 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 40
			// srcs: (1959, 727)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd727 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 40
			// srcs: (1961, 728)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd728 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 40
			// srcs: (1962, 729)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd729 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 40
			// srcs: (1964, 730)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd730 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 40
			// srcs: (1965, 731)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd731 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 48
			// srcs: (1967, 732)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd732 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 48
			// srcs: (1968, 733)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd733 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 48
			// srcs: (1970, 734)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd734 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 48
			// srcs: (1971, 735)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd735 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 16
			// srcs: (1972, 736)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd736 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 48
			// srcs: (1973, 737)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd737 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 48
			// srcs: (1974, 738)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd738 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 16
			// srcs: (1975, 739)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd739 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 48
			// srcs: (1976, 740)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd740 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 56
			// srcs: (1977, 741)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd741 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 16
			// srcs: (1978, 742)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd742 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 56
			// srcs: (1979, 743)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd743 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 56
			// srcs: (1980, 744)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd744 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 16
			// srcs: (1981, 745)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd745 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 56
			// srcs: (1982, 746)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd746 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 56
			// srcs: (1983, 747)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd747 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 16
			// srcs: (1984, 748)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd748 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 56
			// srcs: (1985, 749)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd749 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 56
			// srcs: (1986, 750)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd750 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 16
			// srcs: (1987, 751)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd751 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 0
			// srcs: (1988, 752)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd752 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 0
			// srcs: (1989, 753)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd753 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 16
			// srcs: (1990, 754)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd754 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 0
			// srcs: (1991, 755)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd755 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 0
			// srcs: (1992, 756)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd756 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 24
			// srcs: (1993, 757)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd757 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 0
			// srcs: (1994, 758)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd758 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 0
			// srcs: (1995, 759)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd759 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 0
			// srcs: (1996, 760)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd760 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 24
			// srcs: (2000, 761)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd761 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 24
			// srcs: (2003, 762)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd762 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 24
			// srcs: (2006, 763)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd763 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 16
			// srcs: (2007, 764)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd764 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 16
			// srcs: (2008, 765)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd765 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 24
			// srcs: (2009, 766)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd766 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 16
			// srcs: (2010, 767)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd767 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 16
			// srcs: (2011, 768)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd768 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 24
			// srcs: (2012, 769)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd769 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 16
			// srcs: (2013, 770)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd770 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 16
			// srcs: (2014, 771)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd771 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 24
			// srcs: (2015, 772)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd772 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 16
			// srcs: (2016, 773)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd773 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 24
			// srcs: (2017, 774)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd774 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 32
			// srcs: (2018, 775)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd775 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 24
			// srcs: (2019, 776)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd776 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 24
			// srcs: (2020, 777)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd777 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 32
			// srcs: (2021, 778)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd778 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 24
			// srcs: (2022, 779)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd779 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 24
			// srcs: (2023, 780)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd780 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 32
			// srcs: (2024, 781)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd781 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 24
			// srcs: (2025, 782)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd782 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 24
			// srcs: (2026, 783)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd783 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 32
			// srcs: (2027, 784)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd784 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 32
			// srcs: (2028, 785)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd785 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 32
			// srcs: (2029, 786)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd786 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 32
			// srcs: (2030, 787)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd787 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 32
			// srcs: (2031, 788)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd788 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 32
			// srcs: (2032, 789)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd789 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 32
			// srcs: (2033, 790)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd790 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 32
			// srcs: (2034, 791)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd791 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 32
			// srcs: (2035, 792)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd792 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 32
			// srcs: (2036, 793)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd793 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 32
			// srcs: (2037, 794)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd794 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 40
			// srcs: (2038, 795)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd795 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 40
			// srcs: (2039, 796)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd796 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 40
			// srcs: (2040, 797)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd797 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 40
			// srcs: (2041, 798)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd798 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 40
			// srcs: (2042, 799)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd799 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 40
			// srcs: (2043, 800)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd800 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 40
			// srcs: (2044, 801)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd801 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 40
			// srcs: (2045, 802)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd802 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 40
			// srcs: (2046, 803)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd803 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 48
			// srcs: (2047, 804)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd804 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 48
			// srcs: (2048, 805)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd805 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 40
			// srcs: (2049, 806)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd806 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 48
			// srcs: (2050, 807)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd807 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 48
			// srcs: (2051, 808)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd808 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 40
			// srcs: (2052, 809)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd809 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 48
			// srcs: (2053, 810)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd810 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 48
			// srcs: (2054, 811)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd811 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 40
			// srcs: (2055, 812)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd812 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 48
			// srcs: (2056, 813)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd813 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 56
			// srcs: (2057, 814)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd814 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 40
			// srcs: (2058, 815)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd815 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 56
			// srcs: (2059, 816)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd816 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 56
			// srcs: (2060, 817)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd817 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 40
			// srcs: (2061, 818)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd818 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 56
			// srcs: (2062, 819)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd819 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 56
			// srcs: (2063, 820)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd820 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 48
			// srcs: (2064, 821)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd821 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 56
			// srcs: (2065, 822)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd822 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 56
			// srcs: (2066, 823)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd823 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 48
			// srcs: (2067, 824)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd824 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 0
			// srcs: (2068, 825)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd825 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 0
			// srcs: (2069, 826)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd826 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 48
			// srcs: (2070, 827)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd827 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 0
			// srcs: (2071, 828)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd828 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 0
			// srcs: (2072, 829)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd829 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 48
			// srcs: (2073, 830)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd830 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 0
			// srcs: (2074, 831)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd831 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 0
			// srcs: (2075, 832)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd832 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 48
			// srcs: (2076, 833)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd833 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 0
			// srcs: (2077, 834)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd834 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 48
			// srcs: (2079, 835)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd835 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 48
			// srcs: (2082, 836)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd836 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 56
			// srcs: (2085, 837)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd837 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 56
			// srcs: (2088, 838)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd838 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 16
			// srcs: (2089, 839)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd839 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 16
			// srcs: (2090, 840)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd840 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 56
			// srcs: (2091, 841)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd841 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 16
			// srcs: (2092, 842)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd842 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 16
			// srcs: (2093, 843)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd843 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 16
			// srcs: (2094, 844)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd844 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 16
			// srcs: (2095, 845)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd845 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 16
			// srcs: (2096, 846)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd846 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 24
			// srcs: (2097, 847)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd847 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 56
			// srcs: (2098, 848)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd848 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 24
			// srcs: (2099, 849)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd849 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 24
			// srcs: (2100, 850)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd850 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 56
			// srcs: (2101, 851)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd851 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 24
			// srcs: (2102, 852)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd852 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 24
			// srcs: (2103, 853)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd853 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 56
			// srcs: (2104, 854)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd854 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 24
			// srcs: (2105, 855)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd855 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 24
			// srcs: (2106, 856)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd856 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 56
			// srcs: (2107, 857)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd857 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 32
			// srcs: (2108, 858)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd858 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 32
			// srcs: (2109, 859)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd859 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 0
			// srcs: (2110, 860)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd860 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 32
			// srcs: (2111, 861)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd861 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 32
			// srcs: (2112, 862)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd862 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 0
			// srcs: (2113, 863)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd863 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 32
			// srcs: (2114, 864)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd864 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 32
			// srcs: (2115, 865)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd865 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 0
			// srcs: (2116, 866)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd866 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 32
			// srcs: (2117, 867)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd867 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 40
			// srcs: (2118, 868)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd868 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 0
			// srcs: (2119, 869)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd869 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 40
			// srcs: (2120, 870)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd870 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 40
			// srcs: (2121, 871)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd871 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 0
			// srcs: (2122, 872)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd872 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 40
			// srcs: (2123, 873)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd873 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 40
			// srcs: (2124, 874)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd874 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 0
			// srcs: (2125, 875)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd875 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 40
			// srcs: (2126, 876)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd876 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 40
			// srcs: (2127, 877)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd877 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 0
			// srcs: (2128, 878)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd878 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 48
			// srcs: (2129, 879)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd879 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 48
			// srcs: (2130, 880)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd880 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 48
			// srcs: (2132, 881)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd881 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 48
			// srcs: (2133, 882)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd882 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 48
			// srcs: (2135, 883)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd883 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 48
			// srcs: (2136, 884)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd884 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 48
			// srcs: (2138, 885)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd885 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 56
			// srcs: (2139, 886)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd886 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 56
			// srcs: (2141, 887)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd887 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 56
			// srcs: (2142, 888)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd888 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 56
			// srcs: (2143, 889)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd889 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 56
			// srcs: (2144, 890)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd890 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 56
			// srcs: (2145, 891)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd891 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 56
			// srcs: (2146, 892)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd892 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 0
			// srcs: (2148, 893)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd893 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 0
			// srcs: (2149, 894)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd894 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 0
			// srcs: (2151, 895)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd895 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 0
			// srcs: (2152, 896)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd896 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 0
			// srcs: (2154, 897)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd897 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 0
			// srcs: (2155, 898)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd898 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 16
			// srcs: (2156, 899)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd899 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 0
			// srcs: (2157, 900)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd900 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 16
			// srcs: (2159, 901)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd901 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 16
			// srcs: (2162, 902)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd902 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 16
			// srcs: (2165, 903)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd903 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 16
			// srcs: (2168, 904)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd904 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 16
			// srcs: (2169, 905)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd905 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 16
			// srcs: (2170, 906)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd906 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 16
			// srcs: (2171, 907)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd907 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 16
			// srcs: (2172, 908)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd908 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 16
			// srcs: (2173, 909)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd909 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 16
			// srcs: (2174, 910)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd910 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 16
			// srcs: (2175, 911)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd911 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 16
			// srcs: (2176, 912)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd912 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 24
			// srcs: (2177, 913)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd913 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 16
			// srcs: (2178, 914)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd914 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 24
			// srcs: (2179, 915)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd915 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 24
			// srcs: (2180, 916)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd916 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 24
			// srcs: (2181, 917)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd917 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 24
			// srcs: (2182, 918)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd918 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 24
			// srcs: (2183, 919)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd919 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 24
			// srcs: (2184, 920)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd920 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 24
			// srcs: (2185, 921)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd921 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 24
			// srcs: (2186, 922)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd922 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 24
			// srcs: (2187, 923)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd923 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 24
			// srcs: (2188, 924)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd924 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 24
			// srcs: (2189, 925)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd925 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 32
			// srcs: (2190, 926)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd926 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 32
			// srcs: (2191, 927)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd927 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 32
			// srcs: (2192, 928)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd928 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 32
			// srcs: (2193, 929)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd929 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 32
			// srcs: (2194, 930)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd930 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 32
			// srcs: (2195, 931)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd931 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 24
			// srcs: (2196, 932)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd932 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 32
			// srcs: (2197, 933)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd933 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 40
			// srcs: (2198, 934)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd934 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 24
			// srcs: (2199, 935)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd935 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 40
			// srcs: (2200, 936)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd936 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 40
			// srcs: (2201, 937)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd937 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 32
			// srcs: (2202, 938)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd938 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 40
			// srcs: (2203, 939)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd939 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 40
			// srcs: (2204, 940)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd940 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 32
			// srcs: (2205, 941)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd941 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 40
			// srcs: (2206, 942)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd942 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 40
			// srcs: (2207, 943)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd943 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 32
			// srcs: (2208, 944)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd944 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 48
			// srcs: (2209, 945)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd945 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 48
			// srcs: (2210, 946)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd946 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 32
			// srcs: (2211, 947)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd947 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 48
			// srcs: (2212, 948)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd948 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 48
			// srcs: (2213, 949)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd949 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 32
			// srcs: (2214, 950)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd950 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 48
			// srcs: (2215, 951)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd951 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 48
			// srcs: (2216, 952)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd952 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 32
			// srcs: (2217, 953)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd953 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 48
			// srcs: (2218, 954)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd954 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 56
			// srcs: (2219, 955)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd955 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 32
			// srcs: (2220, 956)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd956 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 56
			// srcs: (2221, 957)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd957 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 56
			// srcs: (2222, 958)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd958 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 40
			// srcs: (2223, 959)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd959 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 56
			// srcs: (2224, 960)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd960 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 56
			// srcs: (2225, 961)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd961 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 40
			// srcs: (2226, 962)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd962 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 56
			// srcs: (2227, 963)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd963 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 56
			// srcs: (2228, 964)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd964 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 40
			// srcs: (2229, 965)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd965 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 0
			// srcs: (2230, 966)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd966 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 0
			// srcs: (2231, 967)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd967 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 40
			// srcs: (2232, 968)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd968 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 0
			// srcs: (2233, 969)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd969 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 0
			// srcs: (2234, 970)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd970 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 40
			// srcs: (2235, 971)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd971 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 0
			// srcs: (2236, 972)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd972 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 0
			// srcs: (2237, 973)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd973 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 40
			// srcs: (2238, 974)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd974 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 0
			// srcs: (2239, 975)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB0
			10'd975 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 10 -> 40
			// srcs: (2245, 976)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd976 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 48
			// srcs: (2248, 977)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd977 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 16
			// srcs: (2249, 978)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd978 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 16
			// srcs: (2250, 979)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd979 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 48
			// srcs: (2251, 980)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd980 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 16
			// srcs: (2252, 981)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd981 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 16
			// srcs: (2253, 982)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd982 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 48
			// srcs: (2254, 983)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd983 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 16
			// srcs: (2255, 984)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd984 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 16
			// srcs: (2256, 985)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd985 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 48
			// srcs: (2257, 986)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd986 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 16
			// srcs: (2258, 987)(3140) 47 --> (3140) 47:PEGB2, pass, PUNB
			10'd987 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 10 -> 24
			// srcs: (2259, 988)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd988 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 48
			// srcs: (2260, 989)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd989 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 24
			// srcs: (2261, 990)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd990 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 24
			// srcs: (2262, 991)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd991 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 48
			// srcs: (2263, 992)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd992 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 24
			// srcs: (2264, 993)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd993 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 24
			// srcs: (2265, 994)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd994 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 48
			// srcs: (2266, 995)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB6
			10'd995 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 10 -> 24
			// srcs: (2267, 996)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd996 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 24
			// srcs: (2268, 997)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB3
			10'd997 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 10 -> 56
			// srcs: (2269, 998)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd998 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 32
			// srcs: (2270, 999)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd999 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 32
			// srcs: (2271, 1000)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd1000 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 56
			// srcs: (2272, 1001)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd1001 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 32
			// srcs: (2273, 1002)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd1002 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 32
			// srcs: (2274, 1003)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd1003 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 56
			// srcs: (2275, 1004)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd1004 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 32
			// srcs: (2276, 1005)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd1005 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 32
			// srcs: (2277, 1006)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd1006 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 56
			// srcs: (2278, 1007)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd1007 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 32
			// srcs: (2279, 1008)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB4
			10'd1008 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 10 -> 40
			// srcs: (2280, 1009)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd1009 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 56
			// srcs: (2281, 1010)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd1010 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 40
			// srcs: (2282, 1011)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd1011 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 40
			// srcs: (2283, 1012)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd1012 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 56
			// srcs: (2284, 1013)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd1013 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 10 -> 40
			// srcs: (2285, 1014)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd1014 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 40
			// srcs: (2286, 1015)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB5
			10'd1015 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 10 -> 56
			// srcs: (2287, 1016)(3140) 47 --> (3140) 47:PEGB2, pass, PUGB7
			10'd1016 : rdata = 48'b110001110000010000000000000000000000000000001111;
			default : rdata = 48'b000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 9) begin
	always @(*) begin
		case(address)
			// PEs: 9, 9 -> 8
			// srcs: (1, 0)(12) -1, (797) -1 --> (1581) 1:ND0, NW0, *, PEGB0
			10'd0 : rdata = 48'b000110110000000001000000000000000000000010000000;
			// PEs: 9, 9 -> 8
			// srcs: (2, 1)(94) -3, (879) 1 --> (1663) -3:ND1, NW1, *, PEGB0
			10'd1 : rdata = 48'b000110110000000101000000001000000000000010000000;
			// PEs: 9, 9 -> 8
			// srcs: (3, 2)(174) -1, (959) -1 --> (1743) 1:ND2, NW2, *, PEGB0
			10'd2 : rdata = 48'b000110110000001001000000010000000000000010000000;
			// PEs: 9, 9 -> 8
			// srcs: (4, 3)(254) -1, (1039) 0 --> (1823) 0:ND3, NW3, *, PEGB0
			10'd3 : rdata = 48'b000110110000001101000000011000000000000010000000;
			// PEs: 9, 9 -> 14
			// srcs: (5, 4)(336) 1, (1121) 0 --> (1905) 0:ND4, NW4, *, PEGB6
			10'd4 : rdata = 48'b000110110000010001000000100000000000000011100000;
			// PEs: 9, 9 -> 15
			// srcs: (6, 5)(416) -1, (1201) 1 --> (1985) -1:ND5, NW5, *, PEGB7
			10'd5 : rdata = 48'b000110110000010101000000101000000000000011110000;
			// PEs: 9, 9 -> 14
			// srcs: (7, 6)(497) 0, (1282) 2 --> (2066) 0:ND6, NW6, *, PEGB6
			10'd6 : rdata = 48'b000110110000011001000000110000000000000011100000;
			// PEs: 9, 9 -> 9
			// srcs: (8, 7)(578) 1, (1363) 1 --> (2147) 1:ND7, NW7, *, NI0
			10'd7 : rdata = 48'b000110110000011101000000111100000000000000000000;
			// PEs: 9, 9 -> 9
			// srcs: (9, 8)(658) 1, (1443) 1 --> (2227) 1:ND8, NW8, *, NI1
			10'd8 : rdata = 48'b000110110000100001000001000100001000000000000000;
			// PEs: 9, 9 -> 9
			// srcs: (10, 9)(740) -3, (1525) -3 --> (2309) 9:ND9, NW9, *, NI2
			10'd9 : rdata = 48'b000110110000100101000001001100010000000000000000;
			// PEs: 9, 9 -> 9
			// srcs: (11, 10)(83) -3, (868) 0 --> (1652) 0:ND10, NW10, *, NI3
			10'd10 : rdata = 48'b000110110000101001000001010100011000000000000000;
			// PEs: 9, 9 -> 8
			// srcs: (12, 11)(267) -2, (1052) -3 --> (1836) 6:ND11, NW11, *, PEGB0
			10'd11 : rdata = 48'b000110110000101101000001011000000000000010000000;
			// PEs: 9, 9 -> 9
			// srcs: (13, 12)(451) 1, (1236) 1 --> (2020) 1:ND12, NW12, *, NI4
			10'd12 : rdata = 48'b000110110000110001000001100100100000000000000000;
			// PEs: 9, 9 -> 9
			// srcs: (14, 13)(631) -3, (1416) 1 --> (2200) -3:ND13, NW13, *, NI5
			10'd13 : rdata = 48'b000110110000110101000001101100101000000000000000;
			// PEs: 8 -> 
			// srcs: (40, 14)(1676) -6 --> (1676) -6:PENB, pass, 
			10'd14 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 8, 9 -> 8
			// srcs: (46, 15)(1675) 4, (1676) -6 --> (2457) -2:PENB, ALU, +, PEGB0
			10'd15 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 8 -> 
			// srcs: (58, 16)(1755) -4 --> (1755) -4:PENB, pass, 
			10'd16 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 8, 9 -> 8
			// srcs: (64, 17)(1754) 0, (1755) -4 --> (2533) -4:PENB, ALU, +, PEGB0
			10'd17 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 8 -> 
			// srcs: (71, 18)(1896) -3 --> (1896) -3:PENB, pass, 
			10'd18 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 8, 9 -> 9
			// srcs: (77, 19)(1895) -4, (1896) -3 --> (2675) -7:PENB, ALU, +, NI6
			10'd19 : rdata = 48'b000011101111111000111111111100110000000000000000;
			// PEs: 8 -> 
			// srcs: (79, 20)(1899) 0 --> (1899) 0:PENB, pass, 
			10'd20 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 8, 9 -> 8
			// srcs: (85, 21)(1898) 4, (1899) 0 --> (2678) 4:PENB, ALU, +, PEGB0
			10'd21 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 8 -> 
			// srcs: (87, 22)(1902) -6 --> (1902) -6:PENB, pass, 
			10'd22 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 8, 9 -> 8
			// srcs: (93, 23)(1901) -2, (1902) -6 --> (2680) -8:PENB, ALU, +, PEGB0
			10'd23 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 8 -> 
			// srcs: (95, 24)(1976) -3 --> (1976) -3:PENB, pass, 
			10'd24 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 8, 9 -> 8
			// srcs: (101, 25)(1975) -2, (1976) -3 --> (2756) -5:PENB, ALU, +, PEGB0
			10'd25 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 8 -> 
			// srcs: (103, 26)(1979) 0 --> (1979) 0:PENB, pass, 
			10'd26 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 8, 9 -> 8
			// srcs: (109, 27)(1978) 0, (1979) 0 --> (2760) 0:PENB, ALU, +, PEGB0
			10'd27 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 8 -> 
			// srcs: (111, 28)(1982) 0 --> (1982) 0:PENB, pass, 
			10'd28 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 8, 9 -> 8
			// srcs: (117, 29)(1981) -6, (1982) 0 --> (2762) -6:PENB, ALU, +, PEGB0
			10'd29 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 8 -> 
			// srcs: (119, 30)(2058) 0 --> (2058) 0:PENB, pass, 
			10'd30 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 8, 9 -> 9
			// srcs: (125, 31)(2057) 0, (2058) 0 --> (2836) 0:PENB, ALU, +, NI7
			10'd31 : rdata = 48'b000011101111111000111111111100111000000000000000;
			// PEs: 8 -> 
			// srcs: (127, 32)(2061) -2 --> (2061) -2:PENB, pass, 
			10'd32 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 8, 9 -> 9
			// srcs: (133, 33)(2060) -6, (2061) -2 --> (2838) -8:PENB, ALU, +, NI8
			10'd33 : rdata = 48'b000011101111111000111111111101000000000000000000;
			// PEs: 8 -> 
			// srcs: (135, 34)(2138) 0 --> (2138) 0:PENB, pass, 
			10'd34 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 8, 9 -> 9
			// srcs: (141, 35)(2137) 0, (2138) 0 --> (2917) 0:PENB, ALU, +, NI9
			10'd35 : rdata = 48'b000011101111111000111111111101001000000000000000;
			// PEs: 8 -> 
			// srcs: (143, 36)(2141) -2 --> (2141) -2:PENB, pass, 
			10'd36 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 8, 9 -> 9
			// srcs: (149, 37)(2140) 2, (2141) -2 --> (2919) 0:PENB, ALU, +, NI10
			10'd37 : rdata = 48'b000011101111111000111111111101010000000000000000;
			// PEs: 8 -> 9
			// srcs: (151, 38)(2144) 0 --> (2144) 0:PENB, pass, NI11
			10'd38 : rdata = 48'b110001101111111000000000000101011000000000000000;
			// PEs: 9 -> 8
			// srcs: (153, 72)(2020) 1 --> (2020) 1:NI4, pass, PEGB0
			10'd39 : rdata = 48'b110001010000010000000000000000000000000010000000;
			// PEs: 8, 9 -> 8
			// srcs: (157, 39)(2143) 0, (2144) 0 --> (2922) 0:PENB, NI11, +, PEGB0
			10'd40 : rdata = 48'b000011101111111010100001011000000000000010000000;
			// PEs: 8, 9 -> 9
			// srcs: (158, 40)(2146) -4, (2147) 1 --> (2924) -3:PENB, NI0, +, NI4
			10'd41 : rdata = 48'b000011101111111010100000000100100000000000000000;
			// PEs: 8, 9 -> 9
			// srcs: (159, 41)(2226) 0, (2227) 1 --> (3005) 1:PENB, NI1, +, NI0
			10'd42 : rdata = 48'b000011101111111010100000001100000000000000000000;
			// PEs: 9 -> 8
			// srcs: (252, 75)(2836) 0 --> (2836) 0:NI7, pass, PEGB0
			10'd43 : rdata = 48'b110001010000011100000000000000000000000010000000;
			// PEs: 9 -> 8
			// srcs: (253, 76)(2838) -8 --> (2838) -8:NI8, pass, PEGB0
			10'd44 : rdata = 48'b110001010000100000000000000000000000000010000000;
			// PEs: 9 -> 8
			// srcs: (254, 81)(2917) 0 --> (2917) 0:NI9, pass, PEGB0
			10'd45 : rdata = 48'b110001010000100100000000000000000000000010000000;
			// PEs: 9 -> 8
			// srcs: (255, 82)(2919) 0 --> (2919) 0:NI10, pass, PEGB0
			10'd46 : rdata = 48'b110001010000101000000000000000000000000010000000;
			// PEs: 9 -> 8
			// srcs: (266, 83)(2924) -3 --> (2924) -3:NI4, pass, PEGB0
			10'd47 : rdata = 48'b110001010000010000000000000000000000000010000000;
			// PEs: 9 -> 8
			// srcs: (267, 87)(3005) 1 --> (3005) 1:NI0, pass, PEGB0
			10'd48 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 8 -> 
			// srcs: (306, 42)(2064) -3 --> (2064) -3:PENB, pass, 
			10'd49 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 8, 9 -> 10
			// srcs: (312, 43)(2063) 0, (2064) -3 --> (2845) -3:PENB, ALU, +, PENB
			10'd50 : rdata = 48'b000011101111111000111111111000000000000100000000;
			// PEs: 8, 9 -> 13
			// srcs: (326, 44)(2308) 6, (2309) 9 --> (3088) 15:PENB, NI2, +, PEGB5
			10'd51 : rdata = 48'b000011101111111010100000010000000000000011010000;
			// PEs: 10, 8 -> 9
			// srcs: (327, 45)(2381) 2, (1600) -2 --> (2382) 0:PEGB2, PENB, +, NI0
			10'd52 : rdata = 48'b000011110000010011011111110100000000000000000000;
			// PEs: 11, 8 -> 10
			// srcs: (328, 46)(2383) 0, (1603) -3 --> (2384) -3:PEGB3, PENB, +, PENB
			10'd53 : rdata = 48'b000011110000011011011111110000000000000100000000;
			// PEs: 9 -> 10
			// srcs: (335, 95)(2382) 0 --> (2382) 0:NI0, pass, PENB
			10'd54 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 8 -> 
			// srcs: (338, 47)(1634) 3 --> (1634) 3:PENB, pass, 
			10'd55 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 8, 9 -> 8
			// srcs: (344, 48)(2413) -6, (1634) 3 --> (2414) -3:PENB, ALU, +, PEGB0
			10'd56 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 8, 9 -> 8
			// srcs: (345, 49)(2431) 7, (1652) 0 --> (2432) 7:PENB, NI3, +, PEGB0
			10'd57 : rdata = 48'b000011101111111010100000011000000000000010000000;
			// PEs: 8, 13 -> 8
			// srcs: (346, 50)(2442) -6, (1664) 6 --> (2443) 0:PENB, PEGB5, +, PEGB0
			10'd58 : rdata = 48'b000011101111111011100001010000000000000010000000;
			// PEs: 8 -> 
			// srcs: (369, 51)(1692) 0 --> (1692) 0:PENB, pass, 
			10'd59 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 8, 9 -> 8
			// srcs: (375, 52)(2471) 15, (1692) 0 --> (2472) 15:PENB, ALU, +, PEGB0
			10'd60 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 8 -> 
			// srcs: (377, 53)(1719) 6 --> (1719) 6:PENB, pass, 
			10'd61 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 8, 9 -> 9
			// srcs: (383, 54)(2496) 2, (1719) 6 --> (2497) 8:PENB, ALU, +, NI0
			10'd62 : rdata = 48'b000011101111111000111111111100000000000000000000;
			// PEs: 12, 8 -> 8
			// srcs: (384, 55)(2519) -1, (1741) 0 --> (2520) -1:PEGB4, PENB, +, PEGB0
			10'd63 : rdata = 48'b000011110000100011011111110000000000000010000000;
			// PEs: 8 -> 
			// srcs: (386, 56)(1753) -4 --> (1753) -4:PENB, pass, 
			10'd64 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 8, 9 -> 8
			// srcs: (392, 57)(2531) 2, (1753) -4 --> (2532) -2:PENB, ALU, +, PEGB0
			10'd65 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 8 -> 
			// srcs: (394, 58)(1814) -6 --> (1814) -6:PENB, pass, 
			10'd66 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 8, 9 -> 9
			// srcs: (400, 59)(2592) 5, (1814) -6 --> (2593) -1:PENB, ALU, +, NI1
			10'd67 : rdata = 48'b000011101111111000111111111100001000000000000000;
			// PEs: 13, 8 -> 10
			// srcs: (401, 60)(2594) -3, (1817) -1 --> (2595) -4:PEGB5, PENB, +, PENB
			10'd68 : rdata = 48'b000011110000101011011111110000000000000100000000;
			// PEs: 9 -> 10
			// srcs: (408, 101)(2593) -1 --> (2593) -1:NI1, pass, PENB
			10'd69 : rdata = 48'b110001010000000100000000000000000000000100000000;
			// PEs: 8, 13 -> 8
			// srcs: (409, 61)(2626) 0, (1848) 6 --> (2627) 6:PENB, PEGB5, +, PEGB0
			10'd70 : rdata = 48'b000011101111111011100001010000000000000010000000;
			// PEs: 8 -> 
			// srcs: (410, 62)(1873) 2 --> (1873) 2:PENB, pass, 
			10'd71 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 8, 9 -> 8
			// srcs: (415, 63)(2652) 3, (1873) 2 --> (2653) 5:PENB, ALU, +, PEGB0
			10'd72 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 9, 8 -> 8
			// srcs: (416, 64)(2675) -7, (1897) -2 --> (2676) -9:NI6, PENB, +, PEGB0
			10'd73 : rdata = 48'b000011010000011011011111110000000000000010000000;
			// PEs: 14, 8 -> 8
			// srcs: (417, 65)(2684) -2, (1906) 6 --> (2685) 4:PEGB6, PENB, +, PEGB0
			10'd74 : rdata = 48'b000011110000110011011111110000000000000010000000;
			// PEs: 8 -> 
			// srcs: (419, 66)(1971) -6 --> (1971) -6:PENB, pass, 
			10'd75 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 8, 9 -> 9
			// srcs: (425, 67)(2751) -4, (1971) -6 --> (2752) -10:PENB, ALU, +, NI1
			10'd76 : rdata = 48'b000011101111111000111111111100001000000000000000;
			// PEs: 8 -> 
			// srcs: (427, 68)(1998) 0 --> (1998) 0:PENB, pass, 
			10'd77 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 8, 9 -> 8
			// srcs: (433, 69)(2777) -3, (1998) 0 --> (2778) -3:PENB, ALU, +, PEGB0
			10'd78 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 8 -> 
			// srcs: (435, 70)(2004) -2 --> (2004) -2:PENB, pass, 
			10'd79 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 8, 9 -> 8
			// srcs: (441, 71)(2783) -2, (2004) -2 --> (2784) -4:PENB, ALU, +, PEGB0
			10'd80 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 8 -> 
			// srcs: (443, 73)(2050) 0 --> (2050) 0:PENB, pass, 
			10'd81 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 8, 9 -> 8
			// srcs: (449, 74)(2827) 1, (2050) 0 --> (2828) 1:PENB, ALU, +, PEGB0
			10'd82 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 8 -> 
			// srcs: (451, 77)(2124) -3 --> (2124) -3:PENB, pass, 
			10'd83 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 8, 9 -> 9
			// srcs: (457, 78)(2901) 6, (2124) -3 --> (2902) 3:PENB, ALU, +, NI2
			10'd84 : rdata = 48'b000011101111111000111111111100010000000000000000;
			// PEs: 8 -> 
			// srcs: (459, 79)(2130) -4 --> (2130) -4:PENB, pass, 
			10'd85 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 8, 9 -> 8
			// srcs: (465, 80)(2907) 2, (2130) -4 --> (2908) -2:PENB, ALU, +, PEGB0
			10'd86 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 8, 9 -> 8
			// srcs: (466, 84)(2978) -4, (2200) -3 --> (2979) -7:PENB, NI5, +, PEGB0
			10'd87 : rdata = 48'b000011101111111010100000101000000000000010000000;
			// PEs: 8, 14 -> 9
			// srcs: (503, 85)(2997) 1, (2219) 0 --> (2998) 1:PENB, PEGB6, +, NI3
			10'd88 : rdata = 48'b000011101111111011100001100100011000000000000000;
			// PEs: 8, 15 -> 10
			// srcs: (515, 86)(2999) 0, (2222) -4 --> (3000) -4:PENB, PEGB7, +, PENB
			10'd89 : rdata = 48'b000011101111111011100001110000000000000100000000;
			// PEs: 8 -> 9
			// srcs: (517, 88)(2295) 1 --> (2295) 1:PENB, pass, NI4
			10'd90 : rdata = 48'b110001101111111000000000000100100000000000000000;
			// PEs: 9 -> 10
			// srcs: (522, 112)(2998) 1 --> (2998) 1:NI3, pass, PENB
			10'd91 : rdata = 48'b110001010000001100000000000000000000000100000000;
			// PEs: 8, 9 -> 8
			// srcs: (523, 89)(3071) -1, (2295) 1 --> (3072) 0:PENB, NI4, +, PEGB0
			10'd92 : rdata = 48'b000011101111111010100000100000000000000010000000;
			// PEs: 14, 8 -> 15
			// srcs: (531, 90)(3091) 0, (2314) 4 --> (3092) 4:PEGB6, PENB, +, PEGB7
			10'd93 : rdata = 48'b000011110000110011011111110000000000000011110000;
			// PEs: 8 -> 
			// srcs: (534, 91)(2338) 0 --> (2338) 0:PENB, pass, 
			10'd94 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 8, 9 -> 8
			// srcs: (540, 92)(3114) 4, (2338) 0 --> (3115) 4:PENB, ALU, +, PEGB0
			10'd95 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 8 -> 
			// srcs: (550, 93)(2353) 1 --> (2353) 1:PENB, pass, 
			10'd96 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 8, 9 -> 8
			// srcs: (556, 94)(3128) 8, (2353) 1 --> (3129) 9:PENB, ALU, +, PEGB0
			10'd97 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 8 -> 
			// srcs: (558, 96)(2425) -5 --> (2425) -5:PENB, pass, 
			10'd98 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 8, 9 -> 8
			// srcs: (564, 97)(2423) -3, (2425) -5 --> (2426) -8:PENB, ALU, +, PEGB0
			10'd99 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 8 -> 
			// srcs: (566, 98)(2486) 17 --> (2486) 17:PENB, pass, 
			10'd100 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 8, 9 -> 8
			// srcs: (572, 99)(2484) -3, (2486) 17 --> (2487) 14:PENB, ALU, +, PEGB0
			10'd101 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 8, 9 -> 8
			// srcs: (573, 100)(2495) 5, (2497) 8 --> (2498) 13:PENB, NI0, +, PEGB0
			10'd102 : rdata = 48'b000011101111111010100000000000000000000010000000;
			// PEs: 8 -> 
			// srcs: (575, 102)(2632) 0 --> (2632) 0:PENB, pass, 
			10'd103 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 8, 9 -> 9
			// srcs: (581, 103)(2630) 3, (2632) 0 --> (2633) 3:PENB, ALU, +, NI0
			10'd104 : rdata = 48'b000011101111111000111111111100000000000000000000;
			// PEs: 8, 9 -> 9
			// srcs: (582, 104)(2750) -1, (2752) -10 --> (2753) -11:PENB, NI1, +, NI3
			10'd105 : rdata = 48'b000011101111111010100000001100011000000000000000;
			// PEs: 8 -> 
			// srcs: (597, 105)(2763) -4 --> (2763) -4:PENB, pass, 
			10'd106 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 8, 9 -> 8
			// srcs: (603, 106)(2761) 0, (2763) -4 --> (2764) -4:PENB, ALU, +, PEGB0
			10'd107 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 10, 8 -> 8
			// srcs: (630, 107)(2847) -3, (2849) -1 --> (2850) -4:PEGB2, PENB, +, PEGB0
			10'd108 : rdata = 48'b000011110000010011011111110000000000000010000000;
			// PEs: 8, 9 -> 9
			// srcs: (631, 108)(2900) 13, (2902) 3 --> (2903) 16:PENB, NI2, +, NI1
			10'd109 : rdata = 48'b000011101111111010100000010100001000000000000000;
			// PEs: 8 -> 
			// srcs: (632, 109)(2958) 0 --> (2958) 0:PENB, pass, 
			10'd110 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 8, 9 -> 8
			// srcs: (638, 110)(2956) 11, (2958) 0 --> (2959) 11:PENB, ALU, +, PEGB0
			10'd111 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 8, 11 -> 10
			// srcs: (639, 111)(2993) -2, (2995) -4 --> (2996) -6:PENB, PEGB3, +, PENB
			10'd112 : rdata = 48'b000011101111111011100000110000000000000100000000;
			// PEs: 8 -> 
			// srcs: (720, 113)(3120) -4 --> (3120) -4:PENB, pass, 
			10'd113 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 8, 9 -> 9
			// srcs: (726, 114)(3118) -5, (3120) -4 --> (3121) -9:PENB, ALU, +, NI2
			10'd114 : rdata = 48'b000011101111111000111111111100010000000000000000;
			// PEs: 8 -> 
			// srcs: (737, 115)(2449) 6 --> (2449) 6:PENB, pass, 
			10'd115 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 8, 9 -> 8
			// srcs: (743, 116)(2444) 2, (2449) 6 --> (2450) 8:PENB, ALU, +, PEGB0
			10'd116 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 8, 10 -> 9
			// srcs: (744, 117)(2591) 14, (2596) -5 --> (2597) 9:PENB, PEGB2, +, NI4
			10'd117 : rdata = 48'b000011101111111011100000100100100000000000000000;
			// PEs: 8, 9 -> 8
			// srcs: (970, 118)(2628) 16, (2633) 3 --> (2634) 19:PENB, NI0, +, PEGB0
			10'd118 : rdata = 48'b000011101111111010100000000000000000000010000000;
			// PEs: 9, 8 -> 8
			// srcs: (987, 119)(2753) -11, (2758) -7 --> (2759) -18:NI3, PENB, +, PEGB0
			10'd119 : rdata = 48'b000011010000001111011111110000000000000010000000;
			// PEs: 8, 9 -> 8
			// srcs: (988, 120)(2898) 11, (2903) 16 --> (2904) 27:PENB, NI1, +, PEGB0
			10'd120 : rdata = 48'b000011101111111010100000001000000000000010000000;
			// PEs: 8 -> 
			// srcs: (1121, 121)(2953) -4 --> (2953) -4:PENB, pass, 
			10'd121 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 8, 9 -> 8
			// srcs: (1127, 122)(2948) 10, (2953) -4 --> (2954) 6:PENB, ALU, +, PEGB0
			10'd122 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 15, 8 -> 8
			// srcs: (1128, 123)(3093) 16, (3098) -1 --> (3099) 15:PEGB7, PENB, +, PEGB0
			10'd123 : rdata = 48'b000011110000111011011111110000000000000010000000;
			// PEs: 8, 9 -> 9
			// srcs: (1129, 124)(3116) -2, (3121) -9 --> (3122) -11:PENB, NI2, +, NI0
			10'd124 : rdata = 48'b000011101111111010100000010100000000000000000000;
			// PEs: 8, 9 -> 9
			// srcs: (1176, 125)(2586) -24, (2597) 9 --> (2598) -15:PENB, NI4, +, NI1
			10'd125 : rdata = 48'b000011101111111010100000100100001000000000000000;
			// PEs: 8 -> 
			// srcs: (1399, 126)(2818) -3 --> (2818) -3:PENB, pass, 
			10'd126 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 8, 9 -> 8
			// srcs: (1406, 127)(2807) 6, (2818) -3 --> (2819) 3:PENB, ALU, +, PEGB0
			10'd127 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 9, 8 -> 9
			// srcs: (1407, 128)(3122) -11, (3133) 11 --> (3134) 0:NI0, PENB, +, NI2
			10'd128 : rdata = 48'b000011010000000011011111110100010000000000000000;
			// PEs: 8, 9 -> 8
			// srcs: (1408, 129)(2575) 19, (2598) -15 --> (2599) 4:PENB, NI1, +, PEGB0
			10'd129 : rdata = 48'b000011101111111010100000001000000000000010000000;
			// PEs: 8 -> 
			// srcs: (1410, 130)(2794) -1 --> (2794) -1:PENB, pass, 
			10'd130 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 8, 9 -> 8
			// srcs: (1416, 131)(2771) -20, (2794) -1 --> (2795) -21:PENB, ALU, +, PEGB0
			10'd131 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 8, 9 -> 
			// srcs: (1417, 132)(3111) 3, (3134) 0 --> (3135) 3:PENB, NI2, +, 
			10'd132 : rdata = 48'b000011101111111010100000010000000000000000000000;
			// PEs: 8, 9 -> 8
			// srcs: (1437, 133)(3087) -28, (3135) 3 --> (3136) -25:PENB, ALU, +, PEGB0
			10'd133 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 8 -> 
			// srcs: (1487, 134)(3138) -39 --> (3138) -39:PENB, pass, 
			10'd134 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 8, 9 -> 10
			// srcs: (1494, 135)(2747) 88, (3138) -39 --> (3139) 49:PENB, ALU, +, PENB
			10'd135 : rdata = 48'b000011101111111000111111111000000000000100000000;
			// PEs: 10, 9 -> 
			// srcs: (1513, 136)(3140) 47, (12) -1 --> (3149) -47:PEGB2, ND0, *, 
			10'd136 : rdata = 48'b000111110000010001100000000000000000000000000000;
			// PEs: 9, 9 -> 
			// srcs: (1516, 150)(3) 1, (3149) -47 --> (3933) -47:NM0, ALU, *, 
			10'd137 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 9, 9 -> 9
			// srcs: (1519, 164)(797) -1, (3933) -47 --> (4717) 46:NW0, ALU, -, NW0
			10'd138 : rdata = 48'b000100100000000000111111111000000100000000000000;
			// PEs: 10, 9 -> 
			// srcs: (1583, 137)(3140) 47, (83) -3 --> (3220) -141:PEGB2, ND10, *, 
			10'd139 : rdata = 48'b000111110000010001100001010000000000000000000000;
			// PEs: 9, 9 -> 
			// srcs: (1586, 151)(3) 1, (3220) -141 --> (4004) -141:NM0, ALU, *, 
			10'd140 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 9, 9 -> 9
			// srcs: (1589, 165)(868) 0, (4004) -141 --> (4788) 141:NW10, ALU, -, NW10
			10'd141 : rdata = 48'b000100100000101000111111111000000110100000000000;
			// PEs: 10, 9 -> 
			// srcs: (1594, 138)(3140) 47, (94) -3 --> (3231) -141:PEGB2, ND1, *, 
			10'd142 : rdata = 48'b000111110000010001100000001000000000000000000000;
			// PEs: 9, 9 -> 
			// srcs: (1597, 152)(3) 1, (3231) -141 --> (4015) -141:NM0, ALU, *, 
			10'd143 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 9, 9 -> 9
			// srcs: (1600, 166)(879) 1, (4015) -141 --> (4799) 142:NW1, ALU, -, NW1
			10'd144 : rdata = 48'b000100100000000100111111111000000100010000000000;
			// PEs: 10, 9 -> 
			// srcs: (1674, 139)(3140) 47, (174) -1 --> (3311) -47:PEGB2, ND2, *, 
			10'd145 : rdata = 48'b000111110000010001100000010000000000000000000000;
			// PEs: 9, 9 -> 
			// srcs: (1677, 153)(3) 1, (3311) -47 --> (4095) -47:NM0, ALU, *, 
			10'd146 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 9, 9 -> 9
			// srcs: (1680, 167)(959) -1, (4095) -47 --> (4879) 46:NW2, ALU, -, NW2
			10'd147 : rdata = 48'b000100100000001000111111111000000100100000000000;
			// PEs: 10, 9 -> 
			// srcs: (1754, 140)(3140) 47, (254) -1 --> (3391) -47:PEGB2, ND3, *, 
			10'd148 : rdata = 48'b000111110000010001100000011000000000000000000000;
			// PEs: 9, 9 -> 
			// srcs: (1757, 154)(3) 1, (3391) -47 --> (4175) -47:NM0, ALU, *, 
			10'd149 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 9, 9 -> 9
			// srcs: (1760, 168)(1039) 0, (4175) -47 --> (4959) 47:NW3, ALU, -, NW3
			10'd150 : rdata = 48'b000100100000001100111111111000000100110000000000;
			// PEs: 10, 9 -> 
			// srcs: (1767, 141)(3140) 47, (267) -2 --> (3404) -94:PEGB2, ND11, *, 
			10'd151 : rdata = 48'b000111110000010001100001011000000000000000000000;
			// PEs: 9, 9 -> 
			// srcs: (1770, 155)(3) 1, (3404) -94 --> (4188) -94:NM0, ALU, *, 
			10'd152 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 9, 9 -> 9
			// srcs: (1773, 169)(1052) -3, (4188) -94 --> (4972) 91:NW11, ALU, -, NW11
			10'd153 : rdata = 48'b000100100000101100111111111000000110110000000000;
			// PEs: 10, 9 -> 
			// srcs: (1836, 142)(3140) 47, (336) 1 --> (3473) 47:PEGB2, ND4, *, 
			10'd154 : rdata = 48'b000111110000010001100000100000000000000000000000;
			// PEs: 9, 9 -> 
			// srcs: (1839, 156)(3) 1, (3473) 47 --> (4257) 47:NM0, ALU, *, 
			10'd155 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 9, 9 -> 9
			// srcs: (1842, 170)(1121) 0, (4257) 47 --> (5041) -47:NW4, ALU, -, NW4
			10'd156 : rdata = 48'b000100100000010000111111111000000101000000000000;
			// PEs: 10, 9 -> 
			// srcs: (1916, 143)(3140) 47, (416) -1 --> (3553) -47:PEGB2, ND5, *, 
			10'd157 : rdata = 48'b000111110000010001100000101000000000000000000000;
			// PEs: 9, 9 -> 
			// srcs: (1919, 157)(3) 1, (3553) -47 --> (4337) -47:NM0, ALU, *, 
			10'd158 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 9, 9 -> 9
			// srcs: (1922, 171)(1201) 1, (4337) -47 --> (5121) 48:NW5, ALU, -, NW5
			10'd159 : rdata = 48'b000100100000010100111111111000000101010000000000;
			// PEs: 10, 9 -> 
			// srcs: (1951, 144)(3140) 47, (451) 1 --> (3588) 47:PEGB2, ND12, *, 
			10'd160 : rdata = 48'b000111110000010001100001100000000000000000000000;
			// PEs: 9, 9 -> 
			// srcs: (1954, 158)(3) 1, (3588) 47 --> (4372) 47:NM0, ALU, *, 
			10'd161 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 9, 9 -> 9
			// srcs: (1957, 172)(1236) 1, (4372) 47 --> (5156) -46:NW12, ALU, -, NW12
			10'd162 : rdata = 48'b000100100000110000111111111000000111000000000000;
			// PEs: 10, 9 -> 
			// srcs: (1997, 145)(3140) 47, (497) 0 --> (3634) 0:PEGB2, ND6, *, 
			10'd163 : rdata = 48'b000111110000010001100000110000000000000000000000;
			// PEs: 9, 9 -> 
			// srcs: (2000, 159)(3) 1, (3634) 0 --> (4418) 0:NM0, ALU, *, 
			10'd164 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 9, 9 -> 9
			// srcs: (2003, 173)(1282) 2, (4418) 0 --> (5202) 2:NW6, ALU, -, NW6
			10'd165 : rdata = 48'b000100100000011000111111111000000101100000000000;
			// PEs: 10, 9 -> 
			// srcs: (2078, 146)(3140) 47, (578) 1 --> (3715) 47:PEGB2, ND7, *, 
			10'd166 : rdata = 48'b000111110000010001100000111000000000000000000000;
			// PEs: 9, 9 -> 
			// srcs: (2081, 160)(3) 1, (3715) 47 --> (4499) 47:NM0, ALU, *, 
			10'd167 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 9, 9 -> 9
			// srcs: (2084, 174)(1363) 1, (4499) 47 --> (5283) -46:NW7, ALU, -, NW7
			10'd168 : rdata = 48'b000100100000011100111111111000000101110000000000;
			// PEs: 10, 9 -> 
			// srcs: (2131, 147)(3140) 47, (631) -3 --> (3768) -141:PEGB2, ND13, *, 
			10'd169 : rdata = 48'b000111110000010001100001101000000000000000000000;
			// PEs: 9, 9 -> 
			// srcs: (2134, 161)(3) 1, (3768) -141 --> (4552) -141:NM0, ALU, *, 
			10'd170 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 9, 9 -> 9
			// srcs: (2137, 175)(1416) 1, (4552) -141 --> (5336) 142:NW13, ALU, -, NW13
			10'd171 : rdata = 48'b000100100000110100111111111000000111010000000000;
			// PEs: 10, 9 -> 
			// srcs: (2158, 148)(3140) 47, (658) 1 --> (3795) 47:PEGB2, ND8, *, 
			10'd172 : rdata = 48'b000111110000010001100001000000000000000000000000;
			// PEs: 9, 9 -> 
			// srcs: (2161, 162)(3) 1, (3795) 47 --> (4579) 47:NM0, ALU, *, 
			10'd173 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 9, 9 -> 9
			// srcs: (2164, 176)(1443) 1, (4579) 47 --> (5363) -46:NW8, ALU, -, NW8
			10'd174 : rdata = 48'b000100100000100000111111111000000110000000000000;
			// PEs: 10, 9 -> 
			// srcs: (2240, 149)(3140) 47, (740) -3 --> (3877) -141:PEGB2, ND9, *, 
			10'd175 : rdata = 48'b000111110000010001100001001000000000000000000000;
			// PEs: 9, 9 -> 
			// srcs: (2243, 163)(3) 1, (3877) -141 --> (4661) -141:NM0, ALU, *, 
			10'd176 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 9, 9 -> 9
			// srcs: (2246, 177)(1525) -3, (4661) -141 --> (5445) 138:NW9, ALU, -, NW9
			10'd177 : rdata = 48'b000100100000100100111111111000000110010000000000;
			default : rdata = 48'b000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 10) begin
	always @(*) begin
		case(address)
			// PEs: 10, 10 -> 8
			// srcs: (1, 0)(14) 2, (799) -2 --> (1583) -4:ND0, NW0, *, PEGB0
			10'd0 : rdata = 48'b000110110000000001000000000000000000000010000000;
			// PEs: 10, 10 -> 8
			// srcs: (2, 1)(96) -1, (881) 1 --> (1665) -1:ND1, NW1, *, PEGB0
			10'd1 : rdata = 48'b000110110000000101000000001000000000000010000000;
			// PEs: 10, 10 -> 8
			// srcs: (3, 2)(176) -1, (961) -2 --> (1745) 2:ND2, NW2, *, PEGB0
			10'd2 : rdata = 48'b000110110000001001000000010000000000000010000000;
			// PEs: 10, 10 -> 8
			// srcs: (4, 3)(256) -1, (1041) -1 --> (1825) 1:ND3, NW3, *, PEGB0
			10'd3 : rdata = 48'b000110110000001101000000011000000000000010000000;
			// PEs: 10, 10 -> 8
			// srcs: (5, 4)(338) -2, (1123) 0 --> (1907) 0:ND4, NW4, *, PEGB0
			10'd4 : rdata = 48'b000110110000010001000000100000000000000010000000;
			// PEs: 10, 10 -> 8
			// srcs: (6, 5)(418) -2, (1203) -2 --> (1987) 4:ND5, NW5, *, PEGB0
			10'd5 : rdata = 48'b000110110000010101000000101000000000000010000000;
			// PEs: 10, 10 -> 8
			// srcs: (7, 6)(498) 1, (1283) -1 --> (2067) -1:ND6, NW6, *, PEGB0
			10'd6 : rdata = 48'b000110110000011001000000110000000000000010000000;
			// PEs: 10, 10 -> 8
			// srcs: (8, 7)(580) -2, (1365) -2 --> (2149) 4:ND7, NW7, *, PEGB0
			10'd7 : rdata = 48'b000110110000011101000000111000000000000010000000;
			// PEs: 10, 10 -> 10
			// srcs: (9, 8)(660) -3, (1445) 2 --> (2229) -6:ND8, NW8, *, NI0
			10'd8 : rdata = 48'b000110110000100001000001000100000000000000000000;
			// PEs: 10, 10 -> 12
			// srcs: (10, 9)(741) -3, (1526) 1 --> (2310) -3:ND9, NW9, *, PEGB4
			10'd9 : rdata = 48'b000110110000100101000001001000000000000011000000;
			// PEs: 10, 10 -> 8
			// srcs: (11, 10)(86) -3, (871) -2 --> (1655) 6:ND10, NW10, *, PEGB0
			10'd10 : rdata = 48'b000110110000101001000001010000000000000010000000;
			// PEs: 10, 10 -> 10
			// srcs: (12, 11)(270) 2, (1055) -3 --> (1839) -6:ND11, NW11, *, NI1
			10'd11 : rdata = 48'b000110110000101101000001011100001000000000000000;
			// PEs: 10, 10 -> 10
			// srcs: (13, 12)(454) 1, (1239) 1 --> (2023) 1:ND12, NW12, *, NI2
			10'd12 : rdata = 48'b000110110000110001000001100100010000000000000000;
			// PEs: 10, 10 -> 10
			// srcs: (14, 13)(634) 1, (1419) 1 --> (2203) 1:ND13, NW13, *, NI3
			10'd13 : rdata = 48'b000110110000110101000001101100011000000000000000;
			// PEs: 10, 11 -> 10
			// srcs: (15, 18)(2229) -6, (2230) -6 --> (3008) -12:NI0, PEGB3, +, NI4
			10'd14 : rdata = 48'b000011010000000011100000110100100000000000000000;
			// PEs: 8 -> 
			// srcs: (23, 14)(1599) -2 --> (1599) -2:PEGB0, pass, 
			10'd15 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 8, 10 -> 9
			// srcs: (32, 15)(1598) 4, (1599) -2 --> (2381) 2:PEGB0, ALU, +, PEGB1
			10'd16 : rdata = 48'b000011110000000000111111111000000000000010010000;
			// PEs: 8 -> 
			// srcs: (45, 16)(1734) -1 --> (1734) -1:PEGB0, pass, 
			10'd17 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 8, 10 -> 8
			// srcs: (54, 17)(1733) 4, (1734) -1 --> (2514) 3:PEGB0, ALU, +, PEGB0
			10'd18 : rdata = 48'b000011110000000000111111111000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (138, 21)(1839) -6 --> (1839) -6:NI1, pass, PEGB0
			10'd19 : rdata = 48'b110001010000000100000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (148, 22)(2023) 1 --> (2023) 1:NI2, pass, PEGB0
			10'd20 : rdata = 48'b110001010000001000000000000000000000000010000000;
			// PEs: 8 -> 
			// srcs: (247, 19)(1819) 9 --> (1819) 9:PEGB0, pass, 
			10'd21 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 8, 10 -> 11
			// srcs: (256, 20)(1818) 2, (1819) 9 --> (2600) 11:PEGB0, ALU, +, PENB
			10'd22 : rdata = 48'b000011110000000000111111111000000000000100000000;
			// PEs: 10 -> 8
			// srcs: (266, 24)(2203) 1 --> (2203) 1:NI3, pass, PEGB0
			10'd23 : rdata = 48'b110001010000001100000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (279, 25)(3008) -12 --> (3008) -12:NI4, pass, PEGB0
			10'd24 : rdata = 48'b110001010000010000000000000000000000000010000000;
			// PEs: 9, 14 -> 9
			// srcs: (330, 23)(2845) -3, (2846) 0 --> (2847) -3:PENB, PEGB6, +, PEGB1
			10'd25 : rdata = 48'b000011101111111011100001100000000000000010010000;
			// PEs: 9 -> 
			// srcs: (331, 26)(2384) -3 --> (2384) -3:PENB, pass, 
			10'd26 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 9, 10 -> 8
			// srcs: (337, 27)(2382) 0, (2384) -3 --> (2385) -3:PENB, ALU, +, PEGB0
			10'd27 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 9 -> 
			// srcs: (403, 28)(2595) -4 --> (2595) -4:PENB, pass, 
			10'd28 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 9, 10 -> 9
			// srcs: (410, 29)(2593) -1, (2595) -4 --> (2596) -5:PENB, ALU, +, PEGB1
			10'd29 : rdata = 48'b000011101111111000111111111000000000000010010000;
			// PEs: 9 -> 
			// srcs: (517, 30)(3000) -4 --> (3000) -4:PENB, pass, 
			10'd30 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 9, 10 -> 
			// srcs: (524, 31)(2998) 1, (3000) -4 --> (3001) -3:PENB, ALU, +, 
			10'd31 : rdata = 48'b000011101111111000111111111000000000000000000000;
			// PEs: 9, 10 -> 8
			// srcs: (642, 32)(2996) -6, (3001) -3 --> (3002) -9:PENB, ALU, +, PEGB0
			10'd32 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 9, 10 -> 11, 8, 10
			// srcs: (1497, 33)(3139) 49, (788) 2 --> (3140) 47:PENB, ND14, -, NI0, PENB, PEGB0
			10'd33 : rdata = 48'b000101101111111001100001110100000000000110000000;
			// PEs: 10 -> 8
			// srcs: (1499, 34)(3140) 49 --> (3140) 47:ALU, pass, PEGB0
			10'd34 : rdata = 48'b110000011111111100000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1500, 35)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd35 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1501, 36)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd36 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1502, 37)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd37 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1503, 38)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd38 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1504, 39)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd39 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1505, 40)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd40 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 9
			// srcs: (1506, 41)(3140) 47 --> (3140) 47:NI0, pass, PEGB1
			10'd41 : rdata = 48'b110001010000000000000000000000000000000010010000;
			// PEs: 10 -> 8
			// srcs: (1507, 42)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd42 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10, 10 -> 11
			// srcs: (1508, 43)(3140) 47, (14) 2 --> (3151) 94:NI0, ND0, *, PENB
			10'd43 : rdata = 48'b000111010000000001100000000000000000000100000000;
			// PEs: 10 -> 8
			// srcs: (1509, 44)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd44 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 12
			// srcs: (1510, 45)(3140) 47 --> (3140) 47:NI0, pass, PEGB4
			10'd45 : rdata = 48'b110001010000000000000000000000000000000011000000;
			// PEs: 10 -> 13
			// srcs: (1511, 46)(3140) 47 --> (3140) 47:NI0, pass, PEGB5
			10'd46 : rdata = 48'b110001010000000000000000000000000000000011010000;
			// PEs: 10 -> 8
			// srcs: (1512, 47)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd47 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 14
			// srcs: (1513, 48)(3140) 47 --> (3140) 47:NI0, pass, PEGB6
			10'd48 : rdata = 48'b110001010000000000000000000000000000000011100000;
			// PEs: 10 -> 15
			// srcs: (1514, 49)(3140) 47 --> (3140) 47:NI0, pass, PEGB7
			10'd49 : rdata = 48'b110001010000000000000000000000000000000011110000;
			// PEs: 10 -> 8
			// srcs: (1515, 50)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd50 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1516, 51)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd51 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1517, 52)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd52 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1518, 53)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd53 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1519, 54)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd54 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1520, 55)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd55 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1521, 56)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd56 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1522, 57)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd57 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1523, 58)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd58 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1524, 59)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd59 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1525, 60)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd60 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1526, 61)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd61 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1527, 62)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd62 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1528, 63)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd63 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1529, 64)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd64 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1530, 65)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd65 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1531, 66)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd66 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1532, 67)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd67 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1533, 68)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd68 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1534, 69)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd69 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1535, 70)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd70 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1536, 71)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd71 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1537, 72)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd72 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1538, 73)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd73 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1539, 74)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd74 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1540, 75)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd75 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1541, 76)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd76 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1542, 77)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd77 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1543, 78)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd78 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1544, 79)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd79 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1545, 80)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd80 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1546, 81)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd81 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1547, 82)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd82 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1548, 83)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd83 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1549, 84)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd84 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1550, 85)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd85 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1551, 86)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd86 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1552, 87)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd87 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1553, 88)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd88 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1554, 89)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd89 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1555, 90)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd90 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1556, 91)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd91 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1557, 92)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd92 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1558, 93)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd93 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1559, 94)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd94 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1560, 95)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd95 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1561, 96)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd96 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1562, 97)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd97 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1563, 98)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd98 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1564, 99)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd99 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1565, 100)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd100 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1566, 101)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd101 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1567, 102)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd102 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1568, 103)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd103 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1569, 104)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd104 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1570, 105)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd105 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1571, 106)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd106 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1572, 107)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd107 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1573, 108)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd108 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1574, 109)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd109 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1575, 110)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd110 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 9
			// srcs: (1576, 111)(3140) 47 --> (3140) 47:NI0, pass, PEGB1
			10'd111 : rdata = 48'b110001010000000000000000000000000000000010010000;
			// PEs: 10 -> 8
			// srcs: (1577, 112)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd112 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1578, 113)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd113 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10, 10 -> 11
			// srcs: (1579, 114)(3140) 47, (86) -3 --> (3223) -141:NI0, ND10, *, PENB
			10'd114 : rdata = 48'b000111010000000001100001010000000000000100000000;
			// PEs: 10 -> 8
			// srcs: (1580, 115)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd115 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1581, 116)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd116 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 11
			// srcs: (1582, 117)(3140) 47 --> (3140) 47:NI0, pass, PENB
			10'd117 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 10 -> 8
			// srcs: (1583, 118)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd118 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1584, 119)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd119 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 12
			// srcs: (1585, 120)(3140) 47 --> (3140) 47:NI0, pass, PEGB4
			10'd120 : rdata = 48'b110001010000000000000000000000000000000011000000;
			// PEs: 10 -> 8
			// srcs: (1586, 121)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd121 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 9
			// srcs: (1587, 122)(3140) 47 --> (3140) 47:NI0, pass, PEGB1
			10'd122 : rdata = 48'b110001010000000000000000000000000000000010010000;
			// PEs: 10 -> 13
			// srcs: (1588, 123)(3140) 47 --> (3140) 47:NI0, pass, PEGB5
			10'd123 : rdata = 48'b110001010000000000000000000000000000000011010000;
			// PEs: 10, 10 -> 11
			// srcs: (1589, 124)(3140) 47, (96) -1 --> (3233) -47:NI0, ND1, *, PENB
			10'd124 : rdata = 48'b000111010000000001100000001000000000000100000000;
			// PEs: 10 -> 11
			// srcs: (1590, 125)(3140) 47 --> (3140) 47:NI0, pass, PENB
			10'd125 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 10 -> 14
			// srcs: (1591, 126)(3140) 47 --> (3140) 47:NI0, pass, PEGB6
			10'd126 : rdata = 48'b110001010000000000000000000000000000000011100000;
			// PEs: 10 -> 12
			// srcs: (1592, 127)(3140) 47 --> (3140) 47:NI0, pass, PEGB4
			10'd127 : rdata = 48'b110001010000000000000000000000000000000011000000;
			// PEs: 10 -> 13
			// srcs: (1593, 128)(3140) 47 --> (3140) 47:NI0, pass, PEGB5
			10'd128 : rdata = 48'b110001010000000000000000000000000000000011010000;
			// PEs: 10 -> 15
			// srcs: (1594, 129)(3140) 47 --> (3140) 47:NI0, pass, PEGB7
			10'd129 : rdata = 48'b110001010000000000000000000000000000000011110000;
			// PEs: 10 -> 14
			// srcs: (1595, 130)(3140) 47 --> (3140) 47:NI0, pass, PEGB6
			10'd130 : rdata = 48'b110001010000000000000000000000000000000011100000;
			// PEs: 10 -> 15
			// srcs: (1596, 131)(3140) 47 --> (3140) 47:NI0, pass, PEGB7
			10'd131 : rdata = 48'b110001010000000000000000000000000000000011110000;
			// PEs: 10 -> 8
			// srcs: (1597, 132)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd132 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1598, 133)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd133 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1599, 134)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd134 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1600, 135)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd135 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1601, 136)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd136 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1602, 137)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd137 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1603, 138)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd138 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1604, 139)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd139 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1605, 140)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd140 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1606, 141)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd141 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1607, 142)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd142 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1608, 143)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd143 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1609, 144)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd144 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1610, 145)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd145 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1611, 146)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd146 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1612, 147)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd147 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1613, 148)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd148 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1614, 149)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd149 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1615, 150)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd150 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1616, 151)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd151 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1617, 152)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd152 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1618, 153)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd153 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1619, 154)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd154 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1620, 155)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd155 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1621, 156)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd156 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1622, 157)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd157 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1623, 158)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd158 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1624, 159)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd159 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1625, 160)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd160 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1626, 161)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd161 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1627, 162)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd162 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1628, 163)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd163 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1629, 164)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd164 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1630, 165)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd165 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1631, 166)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd166 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1632, 167)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd167 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1633, 168)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd168 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1634, 169)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd169 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1635, 170)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd170 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1636, 171)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd171 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1637, 172)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd172 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1638, 173)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd173 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1639, 174)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd174 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1640, 175)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd175 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1641, 176)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd176 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1642, 177)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd177 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1643, 178)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd178 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1644, 179)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd179 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1645, 180)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd180 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1646, 181)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd181 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1647, 182)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd182 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1648, 183)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd183 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1649, 184)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd184 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1650, 185)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd185 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1651, 186)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd186 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1652, 187)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd187 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1653, 188)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd188 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1654, 189)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd189 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1655, 190)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd190 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1656, 191)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd191 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1657, 192)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd192 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1658, 193)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd193 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1659, 194)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd194 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1660, 195)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd195 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1661, 196)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd196 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1662, 197)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd197 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1663, 198)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd198 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1664, 199)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd199 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1665, 200)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd200 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1666, 201)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd201 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 9
			// srcs: (1667, 202)(3140) 47 --> (3140) 47:NI0, pass, PEGB1
			10'd202 : rdata = 48'b110001010000000000000000000000000000000010010000;
			// PEs: 10 -> 8
			// srcs: (1668, 203)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd203 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10, 10 -> 11
			// srcs: (1669, 204)(3140) 47, (176) -1 --> (3313) -47:NI0, ND2, *, PENB
			10'd204 : rdata = 48'b000111010000000001100000010000000000000100000000;
			// PEs: 10 -> 11
			// srcs: (1670, 205)(3140) 47 --> (3140) 47:NI0, pass, PENB
			10'd205 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 10 -> 8
			// srcs: (1671, 206)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd206 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 12
			// srcs: (1672, 207)(3140) 47 --> (3140) 47:NI0, pass, PEGB4
			10'd207 : rdata = 48'b110001010000000000000000000000000000000011000000;
			// PEs: 10 -> 13
			// srcs: (1673, 208)(3140) 47 --> (3140) 47:NI0, pass, PEGB5
			10'd208 : rdata = 48'b110001010000000000000000000000000000000011010000;
			// PEs: 10 -> 8
			// srcs: (1674, 209)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd209 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 14
			// srcs: (1675, 210)(3140) 47 --> (3140) 47:NI0, pass, PEGB6
			10'd210 : rdata = 48'b110001010000000000000000000000000000000011100000;
			// PEs: 10 -> 15
			// srcs: (1676, 211)(3140) 47 --> (3140) 47:NI0, pass, PEGB7
			10'd211 : rdata = 48'b110001010000000000000000000000000000000011110000;
			// PEs: 10 -> 8
			// srcs: (1677, 212)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd212 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1678, 213)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd213 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1679, 214)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd214 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1680, 215)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd215 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1681, 216)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd216 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1682, 217)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd217 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1683, 218)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd218 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1684, 219)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd219 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1685, 220)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd220 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1686, 221)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd221 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1687, 222)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd222 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1688, 223)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd223 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1689, 224)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd224 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1690, 225)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd225 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1691, 226)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd226 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1692, 227)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd227 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1693, 228)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd228 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1694, 229)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd229 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1695, 230)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd230 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1696, 231)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd231 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1697, 232)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd232 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1698, 233)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd233 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1699, 234)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd234 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1700, 235)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd235 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1701, 236)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd236 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1702, 237)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd237 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1703, 238)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd238 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1704, 239)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd239 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1705, 240)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd240 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1706, 241)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd241 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1707, 242)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd242 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1708, 243)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd243 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1709, 244)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd244 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1710, 245)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd245 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1711, 246)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd246 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1712, 247)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd247 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1713, 248)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd248 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1714, 249)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd249 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1715, 250)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd250 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1716, 251)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd251 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1717, 252)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd252 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1718, 253)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd253 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1719, 254)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd254 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1720, 255)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd255 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1721, 256)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd256 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1722, 257)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd257 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1723, 258)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd258 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1724, 259)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd259 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1725, 260)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd260 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1726, 261)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd261 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1727, 262)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd262 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1728, 263)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd263 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1729, 264)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd264 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1730, 265)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd265 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1731, 266)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd266 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1732, 267)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd267 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1733, 268)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd268 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1734, 269)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd269 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1735, 270)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd270 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1736, 271)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd271 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1737, 272)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd272 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1738, 273)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd273 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1739, 274)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd274 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1740, 275)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd275 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1741, 276)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd276 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1742, 277)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd277 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1743, 278)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd278 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1744, 279)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd279 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1745, 280)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd280 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1746, 281)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd281 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 9
			// srcs: (1747, 282)(3140) 47 --> (3140) 47:NI0, pass, PEGB1
			10'd282 : rdata = 48'b110001010000000000000000000000000000000010010000;
			// PEs: 10 -> 8
			// srcs: (1748, 283)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd283 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10, 10 -> 11
			// srcs: (1749, 284)(3140) 47, (256) -1 --> (3393) -47:NI0, ND3, *, PENB
			10'd284 : rdata = 48'b000111010000000001100000011000000000000100000000;
			// PEs: 10 -> 11
			// srcs: (1750, 285)(3140) 47 --> (3140) 47:NI0, pass, PENB
			10'd285 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 10 -> 8
			// srcs: (1751, 286)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd286 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 12
			// srcs: (1752, 287)(3140) 47 --> (3140) 47:NI0, pass, PEGB4
			10'd287 : rdata = 48'b110001010000000000000000000000000000000011000000;
			// PEs: 10 -> 13
			// srcs: (1753, 288)(3140) 47 --> (3140) 47:NI0, pass, PEGB5
			10'd288 : rdata = 48'b110001010000000000000000000000000000000011010000;
			// PEs: 10 -> 8
			// srcs: (1754, 289)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd289 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 14
			// srcs: (1755, 290)(3140) 47 --> (3140) 47:NI0, pass, PEGB6
			10'd290 : rdata = 48'b110001010000000000000000000000000000000011100000;
			// PEs: 10 -> 15
			// srcs: (1756, 291)(3140) 47 --> (3140) 47:NI0, pass, PEGB7
			10'd291 : rdata = 48'b110001010000000000000000000000000000000011110000;
			// PEs: 10 -> 8
			// srcs: (1757, 292)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd292 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1758, 293)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd293 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1759, 294)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd294 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 9
			// srcs: (1760, 295)(3140) 47 --> (3140) 47:NI0, pass, PEGB1
			10'd295 : rdata = 48'b110001010000000000000000000000000000000010010000;
			// PEs: 10 -> 8
			// srcs: (1761, 296)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd296 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1762, 297)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd297 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10, 10 -> 11
			// srcs: (1763, 298)(3140) 47, (270) 2 --> (3407) 94:NI0, ND11, *, PENB
			10'd298 : rdata = 48'b000111010000000001100001011000000000000100000000;
			// PEs: 10 -> 8
			// srcs: (1764, 299)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd299 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1765, 300)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd300 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 11
			// srcs: (1766, 301)(3140) 47 --> (3140) 47:NI0, pass, PENB
			10'd301 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 10 -> 8
			// srcs: (1767, 302)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd302 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1768, 303)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd303 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 12
			// srcs: (1769, 304)(3140) 47 --> (3140) 47:NI0, pass, PEGB4
			10'd304 : rdata = 48'b110001010000000000000000000000000000000011000000;
			// PEs: 10 -> 8
			// srcs: (1770, 305)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd305 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1771, 306)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd306 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 13
			// srcs: (1772, 307)(3140) 47 --> (3140) 47:NI0, pass, PEGB5
			10'd307 : rdata = 48'b110001010000000000000000000000000000000011010000;
			// PEs: 10 -> 8
			// srcs: (1773, 308)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd308 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1774, 309)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd309 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 14
			// srcs: (1775, 310)(3140) 47 --> (3140) 47:NI0, pass, PEGB6
			10'd310 : rdata = 48'b110001010000000000000000000000000000000011100000;
			// PEs: 10 -> 8
			// srcs: (1776, 311)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd311 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1777, 312)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd312 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 15
			// srcs: (1778, 313)(3140) 47 --> (3140) 47:NI0, pass, PEGB7
			10'd313 : rdata = 48'b110001010000000000000000000000000000000011110000;
			// PEs: 10 -> 8
			// srcs: (1779, 314)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd314 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1780, 315)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd315 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1781, 316)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd316 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1782, 317)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd317 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1783, 318)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd318 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1784, 319)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd319 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1785, 320)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd320 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1786, 321)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd321 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1787, 322)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd322 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1788, 323)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd323 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1789, 324)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd324 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1790, 325)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd325 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1791, 326)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd326 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1792, 327)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd327 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1793, 328)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd328 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1794, 329)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd329 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1795, 330)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd330 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1796, 331)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd331 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1797, 332)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd332 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1798, 333)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd333 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1799, 334)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd334 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1800, 335)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd335 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1801, 336)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd336 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1802, 337)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd337 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1803, 338)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd338 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1804, 339)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd339 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1805, 340)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd340 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1806, 341)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd341 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1807, 342)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd342 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1808, 343)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd343 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1809, 344)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd344 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1810, 345)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd345 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1811, 346)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd346 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1812, 347)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd347 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1813, 348)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd348 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1814, 349)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd349 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1815, 350)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd350 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1816, 351)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd351 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1817, 352)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd352 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1818, 353)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd353 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1819, 354)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd354 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1820, 355)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd355 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1821, 356)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd356 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1822, 357)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd357 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1823, 358)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd358 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1824, 359)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd359 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1825, 360)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd360 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1826, 361)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd361 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1827, 362)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd362 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1828, 363)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd363 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 9
			// srcs: (1829, 364)(3140) 47 --> (3140) 47:NI0, pass, PEGB1
			10'd364 : rdata = 48'b110001010000000000000000000000000000000010010000;
			// PEs: 10 -> 8
			// srcs: (1830, 365)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd365 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10, 10 -> 11
			// srcs: (1831, 366)(3140) 47, (338) -2 --> (3475) -94:NI0, ND4, *, PENB
			10'd366 : rdata = 48'b000111010000000001100000100000000000000100000000;
			// PEs: 10 -> 11
			// srcs: (1832, 367)(3140) 47 --> (3140) 47:NI0, pass, PENB
			10'd367 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 10 -> 8
			// srcs: (1833, 368)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd368 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 12
			// srcs: (1834, 369)(3140) 47 --> (3140) 47:NI0, pass, PEGB4
			10'd369 : rdata = 48'b110001010000000000000000000000000000000011000000;
			// PEs: 10 -> 13
			// srcs: (1835, 370)(3140) 47 --> (3140) 47:NI0, pass, PEGB5
			10'd370 : rdata = 48'b110001010000000000000000000000000000000011010000;
			// PEs: 10 -> 8
			// srcs: (1836, 371)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd371 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 14
			// srcs: (1837, 372)(3140) 47 --> (3140) 47:NI0, pass, PEGB6
			10'd372 : rdata = 48'b110001010000000000000000000000000000000011100000;
			// PEs: 10 -> 15
			// srcs: (1838, 373)(3140) 47 --> (3140) 47:NI0, pass, PEGB7
			10'd373 : rdata = 48'b110001010000000000000000000000000000000011110000;
			// PEs: 10 -> 8
			// srcs: (1839, 374)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd374 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1840, 375)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd375 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1841, 376)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd376 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1842, 377)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd377 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1843, 378)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd378 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1844, 379)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd379 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1845, 380)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd380 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1846, 381)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd381 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1847, 382)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd382 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1848, 383)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd383 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1849, 384)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd384 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1850, 385)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd385 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1851, 386)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd386 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1852, 387)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd387 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1853, 388)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd388 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1854, 389)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd389 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1855, 390)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd390 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1856, 391)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd391 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1857, 392)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd392 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1858, 393)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd393 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1859, 394)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd394 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1860, 395)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd395 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1861, 396)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd396 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1862, 397)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd397 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1863, 398)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd398 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1864, 399)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd399 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1865, 400)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd400 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1866, 401)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd401 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1867, 402)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd402 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1868, 403)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd403 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1869, 404)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd404 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1870, 405)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd405 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1871, 406)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd406 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1872, 407)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd407 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1873, 408)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd408 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1874, 409)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd409 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1875, 410)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd410 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1876, 411)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd411 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1877, 412)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd412 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1878, 413)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd413 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1879, 414)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd414 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1880, 415)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd415 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1881, 416)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd416 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1882, 417)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd417 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1883, 418)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd418 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1884, 419)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd419 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1885, 420)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd420 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1886, 421)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd421 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1887, 422)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd422 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1888, 423)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd423 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1889, 424)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd424 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1890, 425)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd425 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1891, 426)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd426 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1892, 427)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd427 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1893, 428)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd428 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1894, 429)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd429 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1895, 430)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd430 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1896, 431)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd431 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1897, 432)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd432 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1898, 433)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd433 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1899, 434)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd434 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1900, 435)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd435 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1901, 436)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd436 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1902, 437)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd437 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1903, 438)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd438 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1904, 439)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd439 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1905, 440)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd440 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1906, 441)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd441 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1907, 442)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd442 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1908, 443)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd443 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 9
			// srcs: (1909, 444)(3140) 47 --> (3140) 47:NI0, pass, PEGB1
			10'd444 : rdata = 48'b110001010000000000000000000000000000000010010000;
			// PEs: 10 -> 8
			// srcs: (1910, 445)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd445 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10, 10 -> 11
			// srcs: (1911, 446)(3140) 47, (418) -2 --> (3555) -94:NI0, ND5, *, PENB
			10'd446 : rdata = 48'b000111010000000001100000101000000000000100000000;
			// PEs: 10 -> 11
			// srcs: (1912, 447)(3140) 47 --> (3140) 47:NI0, pass, PENB
			10'd447 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 10 -> 8
			// srcs: (1913, 448)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd448 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 12
			// srcs: (1914, 449)(3140) 47 --> (3140) 47:NI0, pass, PEGB4
			10'd449 : rdata = 48'b110001010000000000000000000000000000000011000000;
			// PEs: 10 -> 13
			// srcs: (1915, 450)(3140) 47 --> (3140) 47:NI0, pass, PEGB5
			10'd450 : rdata = 48'b110001010000000000000000000000000000000011010000;
			// PEs: 10 -> 8
			// srcs: (1916, 451)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd451 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 14
			// srcs: (1917, 452)(3140) 47 --> (3140) 47:NI0, pass, PEGB6
			10'd452 : rdata = 48'b110001010000000000000000000000000000000011100000;
			// PEs: 10 -> 15
			// srcs: (1918, 453)(3140) 47 --> (3140) 47:NI0, pass, PEGB7
			10'd453 : rdata = 48'b110001010000000000000000000000000000000011110000;
			// PEs: 10 -> 8
			// srcs: (1919, 454)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd454 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1920, 455)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd455 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1921, 456)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd456 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1922, 457)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd457 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1923, 458)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd458 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1924, 459)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd459 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1925, 460)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd460 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1926, 461)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd461 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1927, 462)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd462 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1928, 463)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd463 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1929, 464)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd464 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1930, 465)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd465 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1931, 466)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd466 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1932, 467)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd467 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1933, 468)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd468 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1934, 469)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd469 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1935, 470)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd470 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1936, 471)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd471 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1937, 472)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd472 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1938, 473)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd473 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1939, 474)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd474 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1940, 475)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd475 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1941, 476)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd476 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1942, 477)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd477 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1943, 478)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd478 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 9
			// srcs: (1944, 479)(3140) 47 --> (3140) 47:NI0, pass, PEGB1
			10'd479 : rdata = 48'b110001010000000000000000000000000000000010010000;
			// PEs: 10 -> 8
			// srcs: (1945, 480)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd480 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1946, 481)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd481 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10, 10 -> 11
			// srcs: (1947, 482)(3140) 47, (454) 1 --> (3591) 47:NI0, ND12, *, PENB
			10'd482 : rdata = 48'b000111010000000001100001100000000000000100000000;
			// PEs: 10 -> 8
			// srcs: (1948, 483)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd483 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1949, 484)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd484 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 11
			// srcs: (1950, 485)(3140) 47 --> (3140) 47:NI0, pass, PENB
			10'd485 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 10 -> 8
			// srcs: (1951, 486)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd486 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1952, 487)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd487 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 12
			// srcs: (1953, 488)(3140) 47 --> (3140) 47:NI0, pass, PEGB4
			10'd488 : rdata = 48'b110001010000000000000000000000000000000011000000;
			// PEs: 10 -> 8
			// srcs: (1954, 489)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd489 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1955, 490)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd490 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 13
			// srcs: (1956, 491)(3140) 47 --> (3140) 47:NI0, pass, PEGB5
			10'd491 : rdata = 48'b110001010000000000000000000000000000000011010000;
			// PEs: 10 -> 8
			// srcs: (1957, 492)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd492 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1958, 493)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd493 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 14
			// srcs: (1959, 494)(3140) 47 --> (3140) 47:NI0, pass, PEGB6
			10'd494 : rdata = 48'b110001010000000000000000000000000000000011100000;
			// PEs: 10 -> 8
			// srcs: (1960, 495)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd495 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1961, 496)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd496 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 15
			// srcs: (1962, 497)(3140) 47 --> (3140) 47:NI0, pass, PEGB7
			10'd497 : rdata = 48'b110001010000000000000000000000000000000011110000;
			// PEs: 10 -> 8
			// srcs: (1963, 498)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd498 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1964, 499)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd499 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1965, 500)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd500 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1966, 501)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd501 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1967, 502)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd502 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1968, 503)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd503 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1969, 504)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd504 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1970, 505)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd505 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1971, 506)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd506 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1972, 507)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd507 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1973, 508)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd508 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1974, 509)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd509 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1975, 510)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd510 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1976, 511)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd511 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1977, 512)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd512 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1978, 513)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd513 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1979, 514)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd514 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1980, 515)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd515 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1981, 516)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd516 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1982, 517)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd517 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1983, 518)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd518 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1984, 519)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd519 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1985, 520)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd520 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1986, 521)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd521 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1987, 522)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd522 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1988, 523)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd523 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (1989, 524)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd524 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 9
			// srcs: (1990, 525)(3140) 47 --> (3140) 47:NI0, pass, PEGB1
			10'd525 : rdata = 48'b110001010000000000000000000000000000000010010000;
			// PEs: 10, 10 -> 11
			// srcs: (1991, 526)(3140) 47, (498) 1 --> (3635) 47:NI0, ND6, *, PENB
			10'd526 : rdata = 48'b000111010000000001100000110000000000000100000000;
			// PEs: 10 -> 11
			// srcs: (1992, 527)(3140) 47 --> (3140) 47:NI0, pass, PENB
			10'd527 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 10 -> 8
			// srcs: (1993, 528)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd528 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 12
			// srcs: (1994, 529)(3140) 47 --> (3140) 47:NI0, pass, PEGB4
			10'd529 : rdata = 48'b110001010000000000000000000000000000000011000000;
			// PEs: 10 -> 13
			// srcs: (1995, 530)(3140) 47 --> (3140) 47:NI0, pass, PEGB5
			10'd530 : rdata = 48'b110001010000000000000000000000000000000011010000;
			// PEs: 10 -> 8
			// srcs: (1996, 531)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd531 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 14
			// srcs: (1997, 532)(3140) 47 --> (3140) 47:NI0, pass, PEGB6
			10'd532 : rdata = 48'b110001010000000000000000000000000000000011100000;
			// PEs: 10 -> 15
			// srcs: (1998, 533)(3140) 47 --> (3140) 47:NI0, pass, PEGB7
			10'd533 : rdata = 48'b110001010000000000000000000000000000000011110000;
			// PEs: 10 -> 8
			// srcs: (1999, 534)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd534 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2000, 535)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd535 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2001, 536)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd536 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2002, 537)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd537 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2003, 538)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd538 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2004, 539)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd539 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2005, 540)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd540 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2006, 541)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd541 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2007, 542)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd542 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2008, 543)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd543 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2009, 544)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd544 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2010, 545)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd545 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2011, 546)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd546 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2012, 547)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd547 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2013, 548)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd548 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2014, 549)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd549 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2015, 550)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd550 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2016, 551)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd551 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2017, 552)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd552 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2018, 553)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd553 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2019, 554)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd554 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2020, 555)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd555 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2021, 556)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd556 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2022, 557)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd557 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2023, 558)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd558 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2024, 559)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd559 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2025, 560)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd560 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2026, 561)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd561 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2027, 562)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd562 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2028, 563)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd563 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2029, 564)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd564 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2030, 565)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd565 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2031, 566)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd566 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2032, 567)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd567 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2033, 568)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd568 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2034, 569)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd569 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2035, 570)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd570 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2036, 571)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd571 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2037, 572)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd572 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2038, 573)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd573 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2039, 574)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd574 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2040, 575)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd575 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2041, 576)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd576 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2042, 577)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd577 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2043, 578)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd578 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2044, 579)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd579 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2045, 580)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd580 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2046, 581)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd581 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2047, 582)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd582 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2048, 583)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd583 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2049, 584)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd584 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2050, 585)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd585 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2051, 586)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd586 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2052, 587)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd587 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2053, 588)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd588 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2054, 589)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd589 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2055, 590)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd590 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2056, 591)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd591 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2057, 592)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd592 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2058, 593)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd593 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2059, 594)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd594 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2060, 595)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd595 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2061, 596)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd596 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2062, 597)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd597 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2063, 598)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd598 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2064, 599)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd599 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2065, 600)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd600 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2066, 601)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd601 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2067, 602)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd602 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2068, 603)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd603 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2069, 604)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd604 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2070, 605)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd605 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 9
			// srcs: (2071, 606)(3140) 47 --> (3140) 47:NI0, pass, PEGB1
			10'd606 : rdata = 48'b110001010000000000000000000000000000000010010000;
			// PEs: 10 -> 8
			// srcs: (2072, 607)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd607 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10, 10 -> 11
			// srcs: (2073, 608)(3140) 47, (580) -2 --> (3717) -94:NI0, ND7, *, PENB
			10'd608 : rdata = 48'b000111010000000001100000111000000000000100000000;
			// PEs: 10 -> 11
			// srcs: (2074, 609)(3140) 47 --> (3140) 47:NI0, pass, PENB
			10'd609 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 10 -> 8
			// srcs: (2075, 610)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd610 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 12
			// srcs: (2076, 611)(3140) 47 --> (3140) 47:NI0, pass, PEGB4
			10'd611 : rdata = 48'b110001010000000000000000000000000000000011000000;
			// PEs: 10 -> 13
			// srcs: (2077, 612)(3140) 47 --> (3140) 47:NI0, pass, PEGB5
			10'd612 : rdata = 48'b110001010000000000000000000000000000000011010000;
			// PEs: 10 -> 8
			// srcs: (2078, 613)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd613 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 14
			// srcs: (2079, 614)(3140) 47 --> (3140) 47:NI0, pass, PEGB6
			10'd614 : rdata = 48'b110001010000000000000000000000000000000011100000;
			// PEs: 10 -> 15
			// srcs: (2080, 615)(3140) 47 --> (3140) 47:NI0, pass, PEGB7
			10'd615 : rdata = 48'b110001010000000000000000000000000000000011110000;
			// PEs: 10 -> 8
			// srcs: (2081, 616)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd616 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2082, 617)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd617 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2083, 618)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd618 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2084, 619)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd619 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2085, 620)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd620 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2086, 621)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd621 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2087, 622)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd622 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2088, 623)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd623 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2089, 624)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd624 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2090, 625)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd625 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2091, 626)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd626 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2092, 627)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd627 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2093, 628)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd628 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2094, 629)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd629 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2095, 630)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd630 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2096, 631)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd631 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2097, 632)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd632 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2098, 633)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd633 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2099, 634)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd634 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2100, 635)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd635 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2101, 636)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd636 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2102, 637)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd637 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2103, 638)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd638 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2104, 639)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd639 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2105, 640)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd640 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2106, 641)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd641 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2107, 642)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd642 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2108, 643)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd643 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2109, 644)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd644 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2110, 645)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd645 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2111, 646)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd646 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2112, 647)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd647 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2113, 648)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd648 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2114, 649)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd649 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2115, 650)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd650 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2116, 651)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd651 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2117, 652)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd652 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2118, 653)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd653 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2119, 654)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd654 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2120, 655)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd655 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2121, 656)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd656 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2122, 657)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd657 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2123, 658)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd658 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 9
			// srcs: (2124, 659)(3140) 47 --> (3140) 47:NI0, pass, PEGB1
			10'd659 : rdata = 48'b110001010000000000000000000000000000000010010000;
			// PEs: 10 -> 8
			// srcs: (2125, 660)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd660 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2126, 661)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd661 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10, 10 -> 11
			// srcs: (2127, 662)(3140) 47, (634) 1 --> (3771) 47:NI0, ND13, *, PENB
			10'd662 : rdata = 48'b000111010000000001100001101000000000000100000000;
			// PEs: 10 -> 8
			// srcs: (2128, 663)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd663 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2129, 664)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd664 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 11
			// srcs: (2130, 665)(3140) 47 --> (3140) 47:NI0, pass, PENB
			10'd665 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 10 -> 8
			// srcs: (2131, 666)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd666 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2132, 667)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd667 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 12
			// srcs: (2133, 668)(3140) 47 --> (3140) 47:NI0, pass, PEGB4
			10'd668 : rdata = 48'b110001010000000000000000000000000000000011000000;
			// PEs: 10 -> 8
			// srcs: (2134, 669)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd669 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2135, 670)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd670 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2136, 671)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd671 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2137, 672)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd672 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2138, 673)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd673 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2139, 674)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd674 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 13
			// srcs: (2140, 675)(3140) 47 --> (3140) 47:NI0, pass, PEGB5
			10'd675 : rdata = 48'b110001010000000000000000000000000000000011010000;
			// PEs: 10 -> 8
			// srcs: (2141, 676)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd676 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2142, 677)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd677 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 14
			// srcs: (2143, 678)(3140) 47 --> (3140) 47:NI0, pass, PEGB6
			10'd678 : rdata = 48'b110001010000000000000000000000000000000011100000;
			// PEs: 10 -> 8
			// srcs: (2144, 679)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd679 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2145, 680)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd680 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 15
			// srcs: (2146, 681)(3140) 47 --> (3140) 47:NI0, pass, PEGB7
			10'd681 : rdata = 48'b110001010000000000000000000000000000000011110000;
			// PEs: 10 -> 8
			// srcs: (2147, 682)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd682 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2148, 683)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd683 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2149, 684)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd684 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2150, 685)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd685 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 9
			// srcs: (2151, 686)(3140) 47 --> (3140) 47:NI0, pass, PEGB1
			10'd686 : rdata = 48'b110001010000000000000000000000000000000010010000;
			// PEs: 10 -> 8
			// srcs: (2152, 687)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd687 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10, 10 -> 11
			// srcs: (2153, 688)(3140) 47, (660) -3 --> (3797) -141:NI0, ND8, *, PENB
			10'd688 : rdata = 48'b000111010000000001100001000000000000000100000000;
			// PEs: 10 -> 11
			// srcs: (2154, 689)(3140) 47 --> (3140) 47:NI0, pass, PENB
			10'd689 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 10 -> 8
			// srcs: (2155, 690)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd690 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 12
			// srcs: (2156, 691)(3140) 47 --> (3140) 47:NI0, pass, PEGB4
			10'd691 : rdata = 48'b110001010000000000000000000000000000000011000000;
			// PEs: 10 -> 13
			// srcs: (2157, 692)(3140) 47 --> (3140) 47:NI0, pass, PEGB5
			10'd692 : rdata = 48'b110001010000000000000000000000000000000011010000;
			// PEs: 10 -> 8
			// srcs: (2158, 693)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd693 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 14
			// srcs: (2159, 694)(3140) 47 --> (3140) 47:NI0, pass, PEGB6
			10'd694 : rdata = 48'b110001010000000000000000000000000000000011100000;
			// PEs: 10 -> 15
			// srcs: (2160, 695)(3140) 47 --> (3140) 47:NI0, pass, PEGB7
			10'd695 : rdata = 48'b110001010000000000000000000000000000000011110000;
			// PEs: 10 -> 8
			// srcs: (2161, 696)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd696 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2162, 697)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd697 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2163, 698)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd698 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2164, 699)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd699 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2165, 700)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd700 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2166, 701)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd701 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2167, 702)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd702 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2168, 703)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd703 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2169, 704)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd704 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2170, 705)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd705 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2171, 706)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd706 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2172, 707)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd707 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2173, 708)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd708 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2174, 709)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd709 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2175, 710)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd710 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2176, 711)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd711 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2177, 712)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd712 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2178, 713)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd713 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2179, 714)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd714 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2180, 715)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd715 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2181, 716)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd716 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2182, 717)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd717 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2183, 718)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd718 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2184, 719)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd719 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2185, 720)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd720 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2186, 721)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd721 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2187, 722)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd722 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2188, 723)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd723 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2189, 724)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd724 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2190, 725)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd725 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2191, 726)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd726 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2192, 727)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd727 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2193, 728)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd728 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2194, 729)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd729 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2195, 730)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd730 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2196, 731)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd731 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2197, 732)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd732 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2198, 733)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd733 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2199, 734)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd734 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2200, 735)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd735 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2201, 736)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd736 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2202, 737)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd737 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2203, 738)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd738 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2204, 739)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd739 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2205, 740)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd740 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2206, 741)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd741 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2207, 742)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd742 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2208, 743)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd743 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2209, 744)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd744 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2210, 745)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd745 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2211, 746)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd746 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2212, 747)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd747 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2213, 748)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd748 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2214, 749)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd749 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2215, 750)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd750 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2216, 751)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd751 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2217, 752)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd752 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2218, 753)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd753 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2219, 754)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd754 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2220, 755)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd755 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2221, 756)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd756 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2222, 757)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd757 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2223, 758)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd758 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2224, 759)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd759 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2225, 760)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd760 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2226, 761)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd761 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2227, 762)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd762 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2228, 763)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd763 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2229, 764)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd764 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2230, 765)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd765 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2231, 766)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd766 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2232, 767)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd767 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 9
			// srcs: (2233, 768)(3140) 47 --> (3140) 47:NI0, pass, PEGB1
			10'd768 : rdata = 48'b110001010000000000000000000000000000000010010000;
			// PEs: 10, 10 -> 11
			// srcs: (2234, 769)(3140) 47, (741) -3 --> (3878) -141:NI0, ND9, *, PENB
			10'd769 : rdata = 48'b000111010000000001100001001000000000000100000000;
			// PEs: 10 -> 11
			// srcs: (2235, 770)(3140) 47 --> (3140) 47:NI0, pass, PENB
			10'd770 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 10 -> 12
			// srcs: (2236, 771)(3140) 47 --> (3140) 47:NI0, pass, PEGB4
			10'd771 : rdata = 48'b110001010000000000000000000000000000000011000000;
			// PEs: 10 -> 13
			// srcs: (2237, 772)(3140) 47 --> (3140) 47:NI0, pass, PEGB5
			10'd772 : rdata = 48'b110001010000000000000000000000000000000011010000;
			// PEs: 10 -> 8
			// srcs: (2238, 773)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd773 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 14
			// srcs: (2239, 774)(3140) 47 --> (3140) 47:NI0, pass, PEGB6
			10'd774 : rdata = 48'b110001010000000000000000000000000000000011100000;
			// PEs: 10 -> 15
			// srcs: (2240, 775)(3140) 47 --> (3140) 47:NI0, pass, PEGB7
			10'd775 : rdata = 48'b110001010000000000000000000000000000000011110000;
			// PEs: 10 -> 8
			// srcs: (2241, 776)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd776 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2242, 777)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd777 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2243, 778)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd778 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2244, 779)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd779 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2245, 780)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd780 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2246, 781)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd781 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2247, 782)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd782 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2248, 783)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd783 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2249, 784)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd784 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2250, 785)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd785 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2251, 786)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd786 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2252, 787)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd787 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2253, 788)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd788 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2254, 789)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd789 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2255, 790)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd790 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2256, 791)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd791 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2257, 792)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd792 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2258, 793)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd793 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2259, 794)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd794 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2260, 795)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd795 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2261, 796)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd796 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2262, 797)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd797 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2263, 798)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd798 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2264, 799)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd799 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2265, 800)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd800 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2266, 801)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd801 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2267, 802)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd802 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2268, 803)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd803 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2269, 804)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd804 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2270, 805)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd805 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2271, 806)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd806 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2272, 807)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd807 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2273, 808)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd808 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2274, 809)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd809 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2275, 810)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd810 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2276, 811)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd811 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2277, 812)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd812 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2278, 813)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd813 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2279, 814)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd814 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10 -> 8
			// srcs: (2280, 815)(3140) 47 --> (3140) 47:NI0, pass, PEGB0
			10'd815 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 10, 11 -> 10
			// srcs: (2281, 816)(799) -2, (3935) 94 --> (4719) -96:NW0, PEGB3, -, NW0
			10'd816 : rdata = 48'b000100100000000011100000110000000100000000000000;
			// PEs: 10, 11 -> 10
			// srcs: (2282, 817)(871) -2, (4007) -141 --> (4791) 139:NW10, PEGB3, -, NW10
			10'd817 : rdata = 48'b000100100000101011100000110000000110100000000000;
			// PEs: 10, 11 -> 10
			// srcs: (2283, 818)(881) 1, (4017) -47 --> (4801) 48:NW1, PEGB3, -, NW1
			10'd818 : rdata = 48'b000100100000000111100000110000000100010000000000;
			// PEs: 10, 11 -> 10
			// srcs: (2284, 819)(961) -2, (4097) -47 --> (4881) 45:NW2, PEGB3, -, NW2
			10'd819 : rdata = 48'b000100100000001011100000110000000100100000000000;
			// PEs: 10, 11 -> 10
			// srcs: (2285, 820)(1041) -1, (4177) -47 --> (4961) 46:NW3, PEGB3, -, NW3
			10'd820 : rdata = 48'b000100100000001111100000110000000100110000000000;
			// PEs: 10, 11 -> 10
			// srcs: (2286, 821)(1055) -3, (4191) 94 --> (4975) -97:NW11, PEGB3, -, NW11
			10'd821 : rdata = 48'b000100100000101111100000110000000110110000000000;
			// PEs: 10, 11 -> 10
			// srcs: (2287, 822)(1123) 0, (4259) -94 --> (5043) 94:NW4, PEGB3, -, NW4
			10'd822 : rdata = 48'b000100100000010011100000110000000101000000000000;
			// PEs: 10, 11 -> 10
			// srcs: (2288, 823)(1203) -2, (4339) -94 --> (5123) 92:NW5, PEGB3, -, NW5
			10'd823 : rdata = 48'b000100100000010111100000110000000101010000000000;
			// PEs: 10, 11 -> 10
			// srcs: (2289, 824)(1239) 1, (4375) 47 --> (5159) -46:NW12, PEGB3, -, NW12
			10'd824 : rdata = 48'b000100100000110011100000110000000111000000000000;
			// PEs: 10, 11 -> 10
			// srcs: (2290, 825)(1283) -1, (4419) 47 --> (5203) -48:NW6, PEGB3, -, NW6
			10'd825 : rdata = 48'b000100100000011011100000110000000101100000000000;
			// PEs: 10, 11 -> 10
			// srcs: (2291, 826)(1365) -2, (4501) -94 --> (5285) 92:NW7, PEGB3, -, NW7
			10'd826 : rdata = 48'b000100100000011111100000110000000101110000000000;
			// PEs: 10, 11 -> 10
			// srcs: (2292, 827)(1419) 1, (4555) 47 --> (5339) -46:NW13, PEGB3, -, NW13
			10'd827 : rdata = 48'b000100100000110111100000110000000111010000000000;
			// PEs: 10, 11 -> 10
			// srcs: (2293, 828)(1445) 2, (4581) -141 --> (5365) 143:NW8, PEGB3, -, NW8
			10'd828 : rdata = 48'b000100100000100011100000110000000110000000000000;
			// PEs: 10, 11 -> 10
			// srcs: (2294, 829)(1526) 1, (4662) -141 --> (5446) 142:NW9, PEGB3, -, NW9
			10'd829 : rdata = 48'b000100100000100111100000110000000110010000000000;
			default : rdata = 48'b000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 11) begin
	always @(*) begin
		case(address)
			// PEs: 11, 11 -> 8
			// srcs: (1, 0)(15) 2, (800) -2 --> (1584) -4:ND0, NW0, *, PEGB0
			10'd0 : rdata = 48'b000110110000000001000000000000000000000010000000;
			// PEs: 11, 11 -> 8
			// srcs: (2, 1)(97) 2, (882) 0 --> (1666) 0:ND1, NW1, *, PEGB0
			10'd1 : rdata = 48'b000110110000000101000000001000000000000010000000;
			// PEs: 11, 11 -> 8
			// srcs: (3, 2)(177) 1, (962) -2 --> (1746) -2:ND2, NW2, *, PEGB0
			10'd2 : rdata = 48'b000110110000001001000000010000000000000010000000;
			// PEs: 11, 11 -> 8
			// srcs: (4, 3)(257) -1, (1042) 2 --> (1826) -2:ND3, NW3, *, PEGB0
			10'd3 : rdata = 48'b000110110000001101000000011000000000000010000000;
			// PEs: 11, 11 -> 8
			// srcs: (5, 4)(339) -3, (1124) 1 --> (1908) -3:ND4, NW4, *, PEGB0
			10'd4 : rdata = 48'b000110110000010001000000100000000000000010000000;
			// PEs: 11, 11 -> 8
			// srcs: (6, 5)(419) -2, (1204) 1 --> (1988) -2:ND5, NW5, *, PEGB0
			10'd5 : rdata = 48'b000110110000010101000000101000000000000010000000;
			// PEs: 11, 11 -> 8
			// srcs: (7, 6)(499) 0, (1284) -2 --> (2068) 0:ND6, NW6, *, PEGB0
			10'd6 : rdata = 48'b000110110000011001000000110000000000000010000000;
			// PEs: 11, 11 -> 8
			// srcs: (8, 7)(581) 1, (1366) 1 --> (2150) 1:ND7, NW7, *, PEGB0
			10'd7 : rdata = 48'b000110110000011101000000111000000000000010000000;
			// PEs: 11, 11 -> 10
			// srcs: (9, 8)(661) -3, (1446) 2 --> (2230) -6:ND8, NW8, *, PEGB2
			10'd8 : rdata = 48'b000110110000100001000001000000000000000010100000;
			// PEs: 11, 11 -> 12
			// srcs: (10, 9)(742) 0, (1527) -1 --> (2311) 0:ND9, NW9, *, PENB
			10'd9 : rdata = 48'b000110110000100101000001001000000000000100000000;
			// PEs: 11, 11 -> 8
			// srcs: (11, 10)(89) 2, (874) 2 --> (1658) 4:ND10, NW10, *, PEGB0
			10'd10 : rdata = 48'b000110110000101001000001010000000000000010000000;
			// PEs: 11, 11 -> 11
			// srcs: (12, 11)(273) -3, (1058) -1 --> (1842) 3:ND11, NW11, *, NI0
			10'd11 : rdata = 48'b000110110000101101000001011100000000000000000000;
			// PEs: 11, 11 -> 11
			// srcs: (13, 12)(457) 1, (1242) -1 --> (2026) -1:ND12, NW12, *, NI1
			10'd12 : rdata = 48'b000110110000110001000001100100001000000000000000;
			// PEs: 11, 11 -> 11
			// srcs: (14, 13)(637) -1, (1422) 2 --> (2206) -2:ND13, NW13, *, NI2
			10'd13 : rdata = 48'b000110110000110101000001101100010000000000000000;
			// PEs: 13 -> 
			// srcs: (15, 18)(2233) 0 --> (2233) 0:PEGB5, pass, 
			10'd14 : rdata = 48'b110001110000101000000000000000000000000000000000;
			// PEs: 12, 11 -> 11
			// srcs: (17, 19)(2232) -4, (2233) 0 --> (3010) -4:PEGB4, ALU, +, NI3
			10'd15 : rdata = 48'b000011110000100000111111111100011000000000000000;
			// PEs: 8 -> 
			// srcs: (24, 14)(1601) 4 --> (1601) 4:PEGB0, pass, 
			10'd16 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 11, 8 -> 9
			// srcs: (33, 15)(1601) 4, (1602) -4 --> (2383) 0:ALU, PEGB0, +, PEGB1
			10'd17 : rdata = 48'b000010011111111111100000000000000000000010010000;
			// PEs: 8 -> 
			// srcs: (47, 16)(1737) 0 --> (1737) 0:PEGB0, pass, 
			10'd18 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 8, 11 -> 8
			// srcs: (56, 17)(1736) -2, (1737) 0 --> (2516) -2:PEGB0, ALU, +, PEGB0
			10'd19 : rdata = 48'b000011110000000000111111111000000000000010000000;
			// PEs: 11 -> 8
			// srcs: (140, 22)(2026) -1 --> (2026) -1:NI1, pass, PEGB0
			10'd20 : rdata = 48'b110001010000000100000000000000000000000010000000;
			// PEs: 11 -> 8
			// srcs: (240, 21)(1842) 3 --> (1842) 3:NI0, pass, PEGB0
			10'd21 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 11 -> 8
			// srcs: (266, 23)(2206) -2 --> (2206) -2:NI2, pass, PEGB0
			10'd22 : rdata = 48'b110001010000001000000000000000000000000010000000;
			// PEs: 11 -> 8
			// srcs: (288, 26)(3010) -4 --> (3010) -4:NI3, pass, PEGB0
			10'd23 : rdata = 48'b110001010000001100000000000000000000000010000000;
			// PEs: 10, 13 -> 8
			// srcs: (295, 20)(2600) 11, (2601) 2 --> (2602) 13:PENB, PEGB5, +, PEGB0
			10'd24 : rdata = 48'b000011101111111011100001010000000000000010000000;
			// PEs: 8 -> 
			// srcs: (463, 24)(2994) -1 --> (2994) -1:PEGB0, pass, 
			10'd25 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 11, 13 -> 9
			// srcs: (472, 25)(2994) -1, (2216) -3 --> (2995) -4:ALU, PEGB5, +, PEGB1
			10'd26 : rdata = 48'b000010011111111111100001010000000000000010010000;
			// PEs: 10, 11 -> 12
			// srcs: (1500, 27)(3140) 47, (15) 2 --> (3152) 94:PENB, ND0, *, PENB
			10'd27 : rdata = 48'b000111101111111001100000000000000000000100000000;
			// PEs: 11, 12 -> 11
			// srcs: (1509, 58)(800) -2, (3936) 94 --> (4720) -96:NW0, PEGB4, -, NW0
			10'd28 : rdata = 48'b000100100000000011100001000000000100000000000000;
			// PEs: 11, 10 -> 10
			// srcs: (1511, 41)(3) 1, (3151) 94 --> (3935) 94:NM0, PENB, *, PEGB2
			10'd29 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 11, 10 -> 10
			// srcs: (1582, 42)(3) 1, (3223) -141 --> (4007) -141:NM0, PENB, *, PEGB2
			10'd30 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 10, 11 -> 12
			// srcs: (1586, 28)(3140) 47, (89) 2 --> (3226) 94:PENB, ND10, *, PENB
			10'd31 : rdata = 48'b000111101111111001100001010000000000000100000000;
			// PEs: 11, 10 -> 10
			// srcs: (1592, 43)(3) 1, (3233) -47 --> (4017) -47:NM0, PENB, *, PEGB2
			10'd32 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 10, 11 -> 11
			// srcs: (1594, 29)(3140) 47, (97) 2 --> (3234) 94:PENB, ND1, *, NI0
			10'd33 : rdata = 48'b000111101111111001100000001100000000000000000000;
			// PEs: 11, 12 -> 11
			// srcs: (1595, 59)(874) 2, (4010) 94 --> (4794) -92:NW10, PEGB4, -, NW10
			10'd34 : rdata = 48'b000100100000101011100001000000000110100000000000;
			// PEs: 11, 11 -> 
			// srcs: (1597, 44)(3) 1, (3234) 94 --> (4018) 94:NM0, NI0, *, 
			10'd35 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 11, 11 -> 11
			// srcs: (1600, 60)(882) 0, (4018) 94 --> (4802) -94:NW1, ALU, -, NW1
			10'd36 : rdata = 48'b000100100000000100111111111000000100010000000000;
			// PEs: 11, 10 -> 10
			// srcs: (1672, 45)(3) 1, (3313) -47 --> (4097) -47:NM0, PENB, *, PEGB2
			10'd37 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 10, 11 -> 12
			// srcs: (1674, 30)(3140) 47, (177) 1 --> (3314) 47:PENB, ND2, *, PENB
			10'd38 : rdata = 48'b000111101111111001100000010000000000000100000000;
			// PEs: 11, 12 -> 11
			// srcs: (1683, 61)(962) -2, (4098) 47 --> (4882) -49:NW2, PEGB4, -, NW2
			10'd39 : rdata = 48'b000100100000001011100001000000000100100000000000;
			// PEs: 11, 10 -> 10
			// srcs: (1752, 46)(3) 1, (3393) -47 --> (4177) -47:NM0, PENB, *, PEGB2
			10'd40 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 10, 11 -> 12
			// srcs: (1754, 31)(3140) 47, (257) -1 --> (3394) -47:PENB, ND3, *, PENB
			10'd41 : rdata = 48'b000111101111111001100000011000000000000100000000;
			// PEs: 11, 12 -> 11
			// srcs: (1763, 62)(1042) 2, (4178) -47 --> (4962) 49:NW3, PEGB4, -, NW3
			10'd42 : rdata = 48'b000100100000001111100001000000000100110000000000;
			// PEs: 11, 10 -> 10
			// srcs: (1766, 47)(3) 1, (3407) 94 --> (4191) 94:NM0, PENB, *, PEGB2
			10'd43 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 10, 11 -> 12
			// srcs: (1770, 32)(3140) 47, (273) -3 --> (3410) -141:PENB, ND11, *, PENB
			10'd44 : rdata = 48'b000111101111111001100001011000000000000100000000;
			// PEs: 11, 12 -> 11
			// srcs: (1779, 63)(1058) -1, (4194) -141 --> (4978) 140:NW11, PEGB4, -, NW11
			10'd45 : rdata = 48'b000100100000101111100001000000000110110000000000;
			// PEs: 11, 10 -> 10
			// srcs: (1834, 48)(3) 1, (3475) -94 --> (4259) -94:NM0, PENB, *, PEGB2
			10'd46 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 10, 11 -> 12
			// srcs: (1836, 33)(3140) 47, (339) -3 --> (3476) -141:PENB, ND4, *, PENB
			10'd47 : rdata = 48'b000111101111111001100000100000000000000100000000;
			// PEs: 11, 12 -> 11
			// srcs: (1845, 64)(1124) 1, (4260) -141 --> (5044) 142:NW4, PEGB4, -, NW4
			10'd48 : rdata = 48'b000100100000010011100001000000000101000000000000;
			// PEs: 11, 10 -> 10
			// srcs: (1914, 49)(3) 1, (3555) -94 --> (4339) -94:NM0, PENB, *, PEGB2
			10'd49 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 10, 11 -> 12
			// srcs: (1916, 34)(3140) 47, (419) -2 --> (3556) -94:PENB, ND5, *, PENB
			10'd50 : rdata = 48'b000111101111111001100000101000000000000100000000;
			// PEs: 11, 12 -> 11
			// srcs: (1925, 65)(1204) 1, (4340) -94 --> (5124) 95:NW5, PEGB4, -, NW5
			10'd51 : rdata = 48'b000100100000010111100001000000000101010000000000;
			// PEs: 11, 10 -> 10
			// srcs: (1950, 50)(3) 1, (3591) 47 --> (4375) 47:NM0, PENB, *, PEGB2
			10'd52 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 10, 11 -> 12
			// srcs: (1954, 35)(3140) 47, (457) 1 --> (3594) 47:PENB, ND12, *, PENB
			10'd53 : rdata = 48'b000111101111111001100001100000000000000100000000;
			// PEs: 11, 12 -> 11
			// srcs: (1963, 66)(1242) -1, (4378) 47 --> (5162) -48:NW12, PEGB4, -, NW12
			10'd54 : rdata = 48'b000100100000110011100001000000000111000000000000;
			// PEs: 11, 10 -> 10
			// srcs: (1994, 51)(3) 1, (3635) 47 --> (4419) 47:NM0, PENB, *, PEGB2
			10'd55 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 10, 11 -> 
			// srcs: (1996, 36)(3140) 47, (499) 0 --> (3636) 0:PENB, ND6, *, 
			10'd56 : rdata = 48'b000111101111111001100000110000000000000000000000;
			// PEs: 11, 11 -> 
			// srcs: (1999, 52)(3) 1, (3636) 0 --> (4420) 0:NM0, ALU, *, 
			10'd57 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 11, 11 -> 11
			// srcs: (2002, 67)(1284) -2, (4420) 0 --> (5204) -2:NW6, ALU, -, NW6
			10'd58 : rdata = 48'b000100100000011000111111111000000101100000000000;
			// PEs: 11, 10 -> 10
			// srcs: (2076, 53)(3) 1, (3717) -94 --> (4501) -94:NM0, PENB, *, PEGB2
			10'd59 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 10, 11 -> 12
			// srcs: (2078, 37)(3140) 47, (581) 1 --> (3718) 47:PENB, ND7, *, PENB
			10'd60 : rdata = 48'b000111101111111001100000111000000000000100000000;
			// PEs: 11, 12 -> 11
			// srcs: (2087, 68)(1366) 1, (4502) 47 --> (5286) -46:NW7, PEGB4, -, NW7
			10'd61 : rdata = 48'b000100100000011111100001000000000101110000000000;
			// PEs: 11, 10 -> 10
			// srcs: (2130, 54)(3) 1, (3771) 47 --> (4555) 47:NM0, PENB, *, PEGB2
			10'd62 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 10, 11 -> 12
			// srcs: (2134, 38)(3140) 47, (637) -1 --> (3774) -47:PENB, ND13, *, PENB
			10'd63 : rdata = 48'b000111101111111001100001101000000000000100000000;
			// PEs: 11, 12 -> 11
			// srcs: (2143, 69)(1422) 2, (4558) -47 --> (5342) 49:NW13, PEGB4, -, NW13
			10'd64 : rdata = 48'b000100100000110111100001000000000111010000000000;
			// PEs: 11, 10 -> 10
			// srcs: (2156, 55)(3) 1, (3797) -141 --> (4581) -141:NM0, PENB, *, PEGB2
			10'd65 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 10, 11 -> 12
			// srcs: (2158, 39)(3140) 47, (661) -3 --> (3798) -141:PENB, ND8, *, PENB
			10'd66 : rdata = 48'b000111101111111001100001000000000000000100000000;
			// PEs: 11, 12 -> 11
			// srcs: (2167, 70)(1446) 2, (4582) -141 --> (5366) 143:NW8, PEGB4, -, NW8
			10'd67 : rdata = 48'b000100100000100011100001000000000110000000000000;
			// PEs: 11, 10 -> 10
			// srcs: (2237, 56)(3) 1, (3878) -141 --> (4662) -141:NM0, PENB, *, PEGB2
			10'd68 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 10, 11 -> 
			// srcs: (2239, 40)(3140) 47, (742) 0 --> (3879) 0:PENB, ND9, *, 
			10'd69 : rdata = 48'b000111101111111001100001001000000000000000000000;
			// PEs: 11, 11 -> 
			// srcs: (2242, 57)(3) 1, (3879) 0 --> (4663) 0:NM0, ALU, *, 
			10'd70 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 11, 11 -> 11
			// srcs: (2245, 71)(1527) -1, (4663) 0 --> (5447) -1:NW9, ALU, -, NW9
			10'd71 : rdata = 48'b000100100000100100111111111000000110010000000000;
			default : rdata = 48'b000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 12) begin
	always @(*) begin
		case(address)
			// PEs: 12, 12 -> 8
			// srcs: (1, 0)(17) -2, (802) 2 --> (1586) -4:ND0, NW0, *, PEGB0
			10'd0 : rdata = 48'b000110110000000001000000000000000000000010000000;
			// PEs: 12, 12 -> 8
			// srcs: (2, 1)(99) -3, (884) -3 --> (1668) 9:ND1, NW1, *, PEGB0
			10'd1 : rdata = 48'b000110110000000101000000001000000000000010000000;
			// PEs: 12, 12 -> 8
			// srcs: (3, 2)(179) 1, (964) -3 --> (1748) -3:ND2, NW2, *, PEGB0
			10'd2 : rdata = 48'b000110110000001001000000010000000000000010000000;
			// PEs: 12, 12 -> 8
			// srcs: (4, 3)(259) 0, (1044) 0 --> (1828) 0:ND3, NW3, *, PEGB0
			10'd3 : rdata = 48'b000110110000001101000000011000000000000010000000;
			// PEs: 12, 12 -> 8
			// srcs: (5, 4)(341) -2, (1126) 1 --> (1910) -2:ND4, NW4, *, PEGB0
			10'd4 : rdata = 48'b000110110000010001000000100000000000000010000000;
			// PEs: 12, 12 -> 8
			// srcs: (6, 5)(421) -1, (1206) 2 --> (1990) -2:ND5, NW5, *, PEGB0
			10'd5 : rdata = 48'b000110110000010101000000101000000000000010000000;
			// PEs: 12, 12 -> 8
			// srcs: (7, 6)(501) 2, (1286) 2 --> (2070) 4:ND6, NW6, *, PEGB0
			10'd6 : rdata = 48'b000110110000011001000000110000000000000010000000;
			// PEs: 12, 12 -> 8
			// srcs: (8, 7)(583) 0, (1368) 1 --> (2152) 0:ND7, NW7, *, PEGB0
			10'd7 : rdata = 48'b000110110000011101000000111000000000000010000000;
			// PEs: 12, 12 -> 11
			// srcs: (9, 8)(663) 2, (1448) -2 --> (2232) -4:ND8, NW8, *, PEGB3
			10'd8 : rdata = 48'b000110110000100001000001000000000000000010110000;
			// PEs: 12, 12 -> 14
			// srcs: (10, 9)(743) -3, (1528) 0 --> (2312) 0:ND9, NW9, *, PEGB6
			10'd9 : rdata = 48'b000110110000100101000001001000000000000011100000;
			// PEs: 12, 12 -> 12
			// srcs: (11, 10)(92) 1, (877) 0 --> (1661) 0:ND10, NW10, *, NI0
			10'd10 : rdata = 48'b000110110000101001000001010100000000000000000000;
			// PEs: 12, 12 -> 12
			// srcs: (12, 11)(276) 0, (1061) -1 --> (1845) 0:ND11, NW11, *, NI1
			10'd11 : rdata = 48'b000110110000101101000001011100001000000000000000;
			// PEs: 12, 12 -> 12
			// srcs: (13, 12)(460) 2, (1245) 0 --> (2029) 0:ND12, NW12, *, NI2
			10'd12 : rdata = 48'b000110110000110001000001100100010000000000000000;
			// PEs: 12, 12 -> 12
			// srcs: (14, 13)(640) 1, (1425) 0 --> (2209) 0:ND13, NW13, *, NI3
			10'd13 : rdata = 48'b000110110000110101000001101100011000000000000000;
			// PEs: 15 -> 12
			// srcs: (15, 18)(2236) -4 --> (2236) -4:PEGB7, pass, NI4
			10'd14 : rdata = 48'b110001110000111000000000000100100000000000000000;
			// PEs: 10, 11 -> 13
			// srcs: (16, 20)(2310) -3, (2311) 0 --> (3089) -3:PEGB2, PENB, +, PENB
			10'd15 : rdata = 48'b000011110000010011011111110000000000000100000000;
			// PEs: 14, 12 -> 12
			// srcs: (17, 19)(2235) 1, (2236) -4 --> (3015) -3:PEGB6, NI4, +, NI5
			10'd16 : rdata = 48'b000011110000110010100000100100101000000000000000;
			// PEs: 8 -> 
			// srcs: (21, 14)(1605) -2 --> (1605) -2:PEGB0, pass, 
			10'd17 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 8, 12 -> 8
			// srcs: (30, 15)(1604) -1, (1605) -2 --> (2386) -3:PEGB0, ALU, +, PEGB0
			10'd18 : rdata = 48'b000011110000000000111111111000000000000010000000;
			// PEs: 8 -> 
			// srcs: (51, 16)(1740) 0 --> (1740) 0:PEGB0, pass, 
			10'd19 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 8, 12 -> 9
			// srcs: (60, 17)(1739) -1, (1740) 0 --> (2519) -1:PEGB0, ALU, +, PEGB1
			10'd20 : rdata = 48'b000011110000000000111111111000000000000010010000;
			// PEs: 12 -> 8
			// srcs: (122, 21)(1661) 0 --> (1661) 0:NI0, pass, PEGB0
			10'd21 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 12 -> 8
			// srcs: (124, 22)(1845) 0 --> (1845) 0:NI1, pass, PEGB0
			10'd22 : rdata = 48'b110001010000000100000000000000000000000010000000;
			// PEs: 12 -> 8
			// srcs: (252, 23)(2029) 0 --> (2029) 0:NI2, pass, PEGB0
			10'd23 : rdata = 48'b110001010000001000000000000000000000000010000000;
			// PEs: 12 -> 8
			// srcs: (266, 24)(2209) 0 --> (2209) 0:NI3, pass, PEGB0
			10'd24 : rdata = 48'b110001010000001100000000000000000000000010000000;
			// PEs: 12 -> 8
			// srcs: (296, 25)(3015) -3 --> (3015) -3:NI5, pass, PEGB0
			10'd25 : rdata = 48'b110001010000010100000000000000000000000010000000;
			// PEs: 12, 11 -> 11
			// srcs: (1503, 40)(3) 1, (3152) 94 --> (3936) 94:NM0, PENB, *, PEGB3
			10'd26 : rdata = 48'b000111000000000011011111110000000000000010110000;
			// PEs: 10, 12 -> 
			// srcs: (1517, 26)(3140) 47, (17) -2 --> (3154) -94:PEGB2, ND0, *, 
			10'd27 : rdata = 48'b000111110000010001100000000000000000000000000000;
			// PEs: 12, 12 -> 
			// srcs: (1520, 41)(3) 1, (3154) -94 --> (3938) -94:NM0, ALU, *, 
			10'd28 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 12, 12 -> 12
			// srcs: (1523, 57)(802) 2, (3938) -94 --> (4722) 96:NW0, ALU, -, NW0
			10'd29 : rdata = 48'b000100100000000000111111111000000100000000000000;
			// PEs: 12, 11 -> 11
			// srcs: (1589, 42)(3) 1, (3226) 94 --> (4010) 94:NM0, PENB, *, PEGB3
			10'd30 : rdata = 48'b000111000000000011011111110000000000000010110000;
			// PEs: 10, 12 -> 
			// srcs: (1592, 27)(3140) 47, (92) 1 --> (3229) 47:PEGB2, ND10, *, 
			10'd31 : rdata = 48'b000111110000010001100001010000000000000000000000;
			// PEs: 12, 12 -> 
			// srcs: (1595, 43)(3) 1, (3229) 47 --> (4013) 47:NM0, ALU, *, 
			10'd32 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 12, 12 -> 12
			// srcs: (1598, 58)(877) 0, (4013) 47 --> (4797) -47:NW10, ALU, -, NW10
			10'd33 : rdata = 48'b000100100000101000111111111000000110100000000000;
			// PEs: 10, 12 -> 13
			// srcs: (1599, 28)(3140) 47, (99) -3 --> (3236) -141:PEGB2, ND1, *, PENB
			10'd34 : rdata = 48'b000111110000010001100000001000000000000100000000;
			// PEs: 12, 13 -> 12
			// srcs: (1608, 59)(884) -3, (4020) -141 --> (4804) 138:NW1, PEGB5, -, NW1
			10'd35 : rdata = 48'b000100100000000111100001010000000100010000000000;
			// PEs: 12, 11 -> 11
			// srcs: (1677, 44)(3) 1, (3314) 47 --> (4098) 47:NM0, PENB, *, PEGB3
			10'd36 : rdata = 48'b000111000000000011011111110000000000000010110000;
			// PEs: 10, 12 -> 13
			// srcs: (1679, 29)(3140) 47, (179) 1 --> (3316) 47:PEGB2, ND2, *, PENB
			10'd37 : rdata = 48'b000111110000010001100000010000000000000100000000;
			// PEs: 12, 13 -> 12
			// srcs: (1688, 60)(964) -3, (4100) 47 --> (4884) -50:NW2, PEGB5, -, NW2
			10'd38 : rdata = 48'b000100100000001011100001010000000100100000000000;
			// PEs: 12, 11 -> 11
			// srcs: (1757, 45)(3) 1, (3394) -47 --> (4178) -47:NM0, PENB, *, PEGB3
			10'd39 : rdata = 48'b000111000000000011011111110000000000000010110000;
			// PEs: 10, 12 -> 13
			// srcs: (1759, 30)(3140) 47, (259) 0 --> (3396) 0:PEGB2, ND3, *, PENB
			10'd40 : rdata = 48'b000111110000010001100000011000000000000100000000;
			// PEs: 12, 13 -> 12
			// srcs: (1768, 61)(1044) 0, (4180) 0 --> (4964) 0:NW3, PEGB5, -, NW3
			10'd41 : rdata = 48'b000100100000001111100001010000000100110000000000;
			// PEs: 12, 11 -> 11
			// srcs: (1773, 46)(3) 1, (3410) -141 --> (4194) -141:NM0, PENB, *, PEGB3
			10'd42 : rdata = 48'b000111000000000011011111110000000000000010110000;
			// PEs: 10, 12 -> 
			// srcs: (1776, 31)(3140) 47, (276) 0 --> (3413) 0:PEGB2, ND11, *, 
			10'd43 : rdata = 48'b000111110000010001100001011000000000000000000000;
			// PEs: 12, 12 -> 
			// srcs: (1779, 47)(3) 1, (3413) 0 --> (4197) 0:NM0, ALU, *, 
			10'd44 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 12, 12 -> 12
			// srcs: (1782, 62)(1061) -1, (4197) 0 --> (4981) -1:NW11, ALU, -, NW11
			10'd45 : rdata = 48'b000100100000101100111111111000000110110000000000;
			// PEs: 12, 11 -> 11
			// srcs: (1839, 48)(3) 1, (3476) -141 --> (4260) -141:NM0, PENB, *, PEGB3
			10'd46 : rdata = 48'b000111000000000011011111110000000000000010110000;
			// PEs: 10, 12 -> 13
			// srcs: (1841, 32)(3140) 47, (341) -2 --> (3478) -94:PEGB2, ND4, *, PENB
			10'd47 : rdata = 48'b000111110000010001100000100000000000000100000000;
			// PEs: 12, 13 -> 12
			// srcs: (1850, 63)(1126) 1, (4262) -94 --> (5046) 95:NW4, PEGB5, -, NW4
			10'd48 : rdata = 48'b000100100000010011100001010000000101000000000000;
			// PEs: 12, 11 -> 11
			// srcs: (1919, 49)(3) 1, (3556) -94 --> (4340) -94:NM0, PENB, *, PEGB3
			10'd49 : rdata = 48'b000111000000000011011111110000000000000010110000;
			// PEs: 10, 12 -> 13
			// srcs: (1921, 33)(3140) 47, (421) -1 --> (3558) -47:PEGB2, ND5, *, PENB
			10'd50 : rdata = 48'b000111110000010001100000101000000000000100000000;
			// PEs: 12, 13 -> 12
			// srcs: (1930, 64)(1206) 2, (4342) -47 --> (5126) 49:NW5, PEGB5, -, NW5
			10'd51 : rdata = 48'b000100100000010111100001010000000101010000000000;
			// PEs: 12, 11 -> 11
			// srcs: (1957, 50)(3) 1, (3594) 47 --> (4378) 47:NM0, PENB, *, PEGB3
			10'd52 : rdata = 48'b000111000000000011011111110000000000000010110000;
			// PEs: 10, 12 -> 
			// srcs: (1960, 34)(3140) 47, (460) 2 --> (3597) 94:PEGB2, ND12, *, 
			10'd53 : rdata = 48'b000111110000010001100001100000000000000000000000;
			// PEs: 12, 12 -> 
			// srcs: (1963, 51)(3) 1, (3597) 94 --> (4381) 94:NM0, ALU, *, 
			10'd54 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 12, 12 -> 12
			// srcs: (1966, 65)(1245) 0, (4381) 94 --> (5165) -94:NW12, ALU, -, NW12
			10'd55 : rdata = 48'b000100100000110000111111111000000111000000000000;
			// PEs: 10, 12 -> 13
			// srcs: (2001, 35)(3140) 47, (501) 2 --> (3638) 94:PEGB2, ND6, *, PENB
			10'd56 : rdata = 48'b000111110000010001100000110000000000000100000000;
			// PEs: 12, 13 -> 12
			// srcs: (2010, 66)(1286) 2, (4422) 94 --> (5206) -92:NW6, PEGB5, -, NW6
			10'd57 : rdata = 48'b000100100000011011100001010000000101100000000000;
			// PEs: 12, 11 -> 11
			// srcs: (2081, 52)(3) 1, (3718) 47 --> (4502) 47:NM0, PENB, *, PEGB3
			10'd58 : rdata = 48'b000111000000000011011111110000000000000010110000;
			// PEs: 10, 12 -> 
			// srcs: (2083, 36)(3140) 47, (583) 0 --> (3720) 0:PEGB2, ND7, *, 
			10'd59 : rdata = 48'b000111110000010001100000111000000000000000000000;
			// PEs: 12, 12 -> 
			// srcs: (2086, 53)(3) 1, (3720) 0 --> (4504) 0:NM0, ALU, *, 
			10'd60 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 12, 12 -> 12
			// srcs: (2089, 67)(1368) 1, (4504) 0 --> (5288) 1:NW7, ALU, -, NW7
			10'd61 : rdata = 48'b000100100000011100111111111000000101110000000000;
			// PEs: 12, 11 -> 11
			// srcs: (2137, 54)(3) 1, (3774) -47 --> (4558) -47:NM0, PENB, *, PEGB3
			10'd62 : rdata = 48'b000111000000000011011111110000000000000010110000;
			// PEs: 10, 12 -> 13
			// srcs: (2140, 37)(3140) 47, (640) 1 --> (3777) 47:PEGB2, ND13, *, PENB
			10'd63 : rdata = 48'b000111110000010001100001101000000000000100000000;
			// PEs: 12, 13 -> 12
			// srcs: (2149, 68)(1425) 0, (4561) 47 --> (5345) -47:NW13, PEGB5, -, NW13
			10'd64 : rdata = 48'b000100100000110111100001010000000111010000000000;
			// PEs: 12, 11 -> 11
			// srcs: (2161, 55)(3) 1, (3798) -141 --> (4582) -141:NM0, PENB, *, PEGB3
			10'd65 : rdata = 48'b000111000000000011011111110000000000000010110000;
			// PEs: 10, 12 -> 
			// srcs: (2163, 38)(3140) 47, (663) 2 --> (3800) 94:PEGB2, ND8, *, 
			10'd66 : rdata = 48'b000111110000010001100001000000000000000000000000;
			// PEs: 12, 12 -> 
			// srcs: (2166, 56)(3) 1, (3800) 94 --> (4584) 94:NM0, ALU, *, 
			10'd67 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 12, 12 -> 12
			// srcs: (2169, 69)(1448) -2, (4584) 94 --> (5368) -96:NW8, ALU, -, NW8
			10'd68 : rdata = 48'b000100100000100000111111111000000110000000000000;
			// PEs: 10, 12 -> 13
			// srcs: (2243, 39)(3140) 47, (743) -3 --> (3880) -141:PEGB2, ND9, *, PENB
			10'd69 : rdata = 48'b000111110000010001100001001000000000000100000000;
			// PEs: 12, 13 -> 12
			// srcs: (2252, 70)(1528) 0, (4664) -141 --> (5448) 141:NW9, PEGB5, -, NW9
			10'd70 : rdata = 48'b000100100000100111100001010000000110010000000000;
			default : rdata = 48'b000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 13) begin
	always @(*) begin
		case(address)
			// PEs: 13, 13 -> 8
			// srcs: (1, 0)(18) -3, (803) -1 --> (1587) 3:ND0, NW0, *, PEGB0
			10'd0 : rdata = 48'b000110110000000001000000000000000000000010000000;
			// PEs: 13, 13 -> 8
			// srcs: (2, 1)(100) 0, (885) -2 --> (1669) 0:ND1, NW1, *, PEGB0
			10'd1 : rdata = 48'b000110110000000101000000001000000000000010000000;
			// PEs: 13, 13 -> 8
			// srcs: (3, 2)(180) 1, (965) 2 --> (1749) 2:ND2, NW2, *, PEGB0
			10'd2 : rdata = 48'b000110110000001001000000010000000000000010000000;
			// PEs: 13, 13 -> 8
			// srcs: (4, 3)(260) -3, (1045) 0 --> (1829) 0:ND3, NW3, *, PEGB0
			10'd3 : rdata = 48'b000110110000001101000000011000000000000010000000;
			// PEs: 13, 13 -> 8
			// srcs: (5, 4)(342) -3, (1127) 0 --> (1911) 0:ND4, NW4, *, PEGB0
			10'd4 : rdata = 48'b000110110000010001000000100000000000000010000000;
			// PEs: 13, 13 -> 8
			// srcs: (6, 5)(422) 1, (1207) 1 --> (1991) 1:ND5, NW5, *, PEGB0
			10'd5 : rdata = 48'b000110110000010101000000101000000000000010000000;
			// PEs: 13, 13 -> 8
			// srcs: (7, 6)(502) -1, (1287) -2 --> (2071) 2:ND6, NW6, *, PEGB0
			10'd6 : rdata = 48'b000110110000011001000000110000000000000010000000;
			// PEs: 13, 13 -> 8
			// srcs: (8, 7)(584) 2, (1369) 2 --> (2153) 4:ND7, NW7, *, PEGB0
			10'd7 : rdata = 48'b000110110000011101000000111000000000000010000000;
			// PEs: 13, 13 -> 11
			// srcs: (9, 8)(664) 1, (1449) 0 --> (2233) 0:ND8, NW8, *, PEGB3
			10'd8 : rdata = 48'b000110110000100001000001000000000000000010110000;
			// PEs: 13, 13 -> 14
			// srcs: (10, 9)(744) 0, (1529) 2 --> (2313) 0:ND9, NW9, *, PENB
			10'd9 : rdata = 48'b000110110000100101000001001000000000000100000000;
			// PEs: 13, 13 -> 9
			// srcs: (11, 10)(95) -3, (880) -2 --> (1664) 6:ND10, NW10, *, PEGB1
			10'd10 : rdata = 48'b000110110000101001000001010000000000000010010000;
			// PEs: 13, 13 -> 13
			// srcs: (12, 11)(279) -2, (1064) -3 --> (1848) 6:ND11, NW11, *, NI0
			10'd11 : rdata = 48'b000110110000101101000001011100000000000000000000;
			// PEs: 13, 13 -> 13
			// srcs: (13, 12)(463) 1, (1248) 0 --> (2032) 0:ND12, NW12, *, NI1
			10'd12 : rdata = 48'b000110110000110001000001100100001000000000000000;
			// PEs: 13, 13 -> 13
			// srcs: (14, 13)(647) 1, (1432) -3 --> (2216) -3:ND13, NW13, *, NI2
			10'd13 : rdata = 48'b000110110000110101000001101100010000000000000000;
			// PEs: 15 -> 
			// srcs: (15, 18)(2316) -4 --> (2316) -4:PEGB7, pass, 
			10'd14 : rdata = 48'b110001110000111000000000000000000000000000000000;
			// PEs: 14, 13 -> 13
			// srcs: (18, 19)(2315) 1, (2316) -4 --> (3094) -3:PEGB6, ALU, +, NI3
			10'd15 : rdata = 48'b000011110000110000111111111100011000000000000000;
			// PEs: 8 -> 
			// srcs: (25, 14)(1608) 0 --> (1608) 0:PEGB0, pass, 
			10'd16 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 8, 13 -> 8
			// srcs: (34, 15)(1607) -2, (1608) 0 --> (2388) -2:PEGB0, ALU, +, PEGB0
			10'd17 : rdata = 48'b000011110000000000111111111000000000000010000000;
			// PEs: 8 -> 
			// srcs: (63, 16)(1816) 0 --> (1816) 0:PEGB0, pass, 
			10'd18 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 8, 13 -> 9
			// srcs: (72, 17)(1815) -3, (1816) 0 --> (2594) -3:PEGB0, ALU, +, PEGB1
			10'd19 : rdata = 48'b000011110000000000111111111000000000000010010000;
			// PEs: 13 -> 8
			// srcs: (156, 23)(2032) 0 --> (2032) 0:NI1, pass, PEGB0
			10'd20 : rdata = 48'b110001010000000100000000000000000000000010000000;
			// PEs: 13 -> 8
			// srcs: (254, 26)(3094) -3 --> (3094) -3:NI3, pass, PEGB0
			10'd21 : rdata = 48'b110001010000001100000000000000000000000010000000;
			// PEs: 8 -> 
			// srcs: (280, 20)(1821) 0 --> (1821) 0:PEGB0, pass, 
			10'd22 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 8, 13 -> 11
			// srcs: (289, 21)(1820) 2, (1821) 0 --> (2601) 2:PEGB0, ALU, +, PEGB3
			10'd23 : rdata = 48'b000011110000000000111111111000000000000010110000;
			// PEs: 9, 12 -> 15
			// srcs: (332, 25)(3088) 15, (3089) -3 --> (3090) 12:PEGB1, PENB, +, PEGB7
			10'd24 : rdata = 48'b000011110000001011011111110000000000000011110000;
			// PEs: 13 -> 9
			// srcs: (404, 22)(1848) 6 --> (1848) 6:NI0, pass, PEGB1
			10'd25 : rdata = 48'b110001010000000000000000000000000000000010010000;
			// PEs: 13 -> 11
			// srcs: (467, 24)(2216) -3 --> (2216) -3:NI2, pass, PEGB3
			10'd26 : rdata = 48'b110001010000001000000000000000000000000010110000;
			// PEs: 10, 13 -> 
			// srcs: (1518, 27)(3140) 47, (18) -3 --> (3155) -141:PEGB2, ND0, *, 
			10'd27 : rdata = 48'b000111110000010001100000000000000000000000000000;
			// PEs: 13, 13 -> 
			// srcs: (1521, 41)(3) 1, (3155) -141 --> (3939) -141:NM0, ALU, *, 
			10'd28 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 13, 13 -> 13
			// srcs: (1524, 57)(803) -1, (3939) -141 --> (4723) 140:NW0, ALU, -, NW0
			10'd29 : rdata = 48'b000100100000000000111111111000000100000000000000;
			// PEs: 10, 13 -> 
			// srcs: (1595, 28)(3140) 47, (95) -3 --> (3232) -141:PEGB2, ND10, *, 
			10'd30 : rdata = 48'b000111110000010001100001010000000000000000000000;
			// PEs: 13, 13 -> 13
			// srcs: (1598, 42)(3) 1, (3232) -141 --> (4016) -141:NM0, ALU, *, NI0
			10'd31 : rdata = 48'b000111000000000000111111111100000000000000000000;
			// PEs: 10, 13 -> 14
			// srcs: (1600, 29)(3140) 47, (100) 0 --> (3237) 0:PEGB2, ND1, *, PENB
			10'd32 : rdata = 48'b000111110000010001100000001000000000000100000000;
			// PEs: 13, 13 -> 13
			// srcs: (1601, 58)(880) -2, (4016) -141 --> (4800) 139:NW10, NI0, -, NW10
			10'd33 : rdata = 48'b000100100000101010100000000000000110100000000000;
			// PEs: 13, 12 -> 12
			// srcs: (1602, 43)(3) 1, (3236) -141 --> (4020) -141:NM0, PENB, *, PEGB4
			10'd34 : rdata = 48'b000111000000000011011111110000000000000011000000;
			// PEs: 13, 14 -> 13
			// srcs: (1609, 59)(885) -2, (4021) 0 --> (4805) -2:NW1, PEGB6, -, NW1
			10'd35 : rdata = 48'b000100100000000111100001100000000100010000000000;
			// PEs: 10, 13 -> 14
			// srcs: (1680, 30)(3140) 47, (180) 1 --> (3317) 47:PEGB2, ND2, *, PENB
			10'd36 : rdata = 48'b000111110000010001100000010000000000000100000000;
			// PEs: 13, 12 -> 12
			// srcs: (1682, 44)(3) 1, (3316) 47 --> (4100) 47:NM0, PENB, *, PEGB4
			10'd37 : rdata = 48'b000111000000000011011111110000000000000011000000;
			// PEs: 13, 14 -> 13
			// srcs: (1689, 60)(965) 2, (4101) 47 --> (4885) -45:NW2, PEGB6, -, NW2
			10'd38 : rdata = 48'b000100100000001011100001100000000100100000000000;
			// PEs: 10, 13 -> 13
			// srcs: (1760, 31)(3140) 47, (260) -3 --> (3397) -141:PEGB2, ND3, *, NI0
			10'd39 : rdata = 48'b000111110000010001100000011100000000000000000000;
			// PEs: 13, 12 -> 12
			// srcs: (1762, 45)(3) 1, (3396) 0 --> (4180) 0:NM0, PENB, *, PEGB4
			10'd40 : rdata = 48'b000111000000000011011111110000000000000011000000;
			// PEs: 13, 13 -> 
			// srcs: (1763, 46)(3) 1, (3397) -141 --> (4181) -141:NM0, NI0, *, 
			10'd41 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 13, 13 -> 13
			// srcs: (1766, 61)(1045) 0, (4181) -141 --> (4965) 141:NW3, ALU, -, NW3
			10'd42 : rdata = 48'b000100100000001100111111111000000100110000000000;
			// PEs: 10, 13 -> 
			// srcs: (1779, 32)(3140) 47, (279) -2 --> (3416) -94:PEGB2, ND11, *, 
			10'd43 : rdata = 48'b000111110000010001100001011000000000000000000000;
			// PEs: 13, 13 -> 
			// srcs: (1782, 47)(3) 1, (3416) -94 --> (4200) -94:NM0, ALU, *, 
			10'd44 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 13, 13 -> 13
			// srcs: (1785, 62)(1064) -3, (4200) -94 --> (4984) 91:NW11, ALU, -, NW11
			10'd45 : rdata = 48'b000100100000101100111111111000000110110000000000;
			// PEs: 10, 13 -> 14
			// srcs: (1842, 33)(3140) 47, (342) -3 --> (3479) -141:PEGB2, ND4, *, PENB
			10'd46 : rdata = 48'b000111110000010001100000100000000000000100000000;
			// PEs: 13, 12 -> 12
			// srcs: (1844, 48)(3) 1, (3478) -94 --> (4262) -94:NM0, PENB, *, PEGB4
			10'd47 : rdata = 48'b000111000000000011011111110000000000000011000000;
			// PEs: 13, 14 -> 13
			// srcs: (1851, 63)(1127) 0, (4263) -141 --> (5047) 141:NW4, PEGB6, -, NW4
			10'd48 : rdata = 48'b000100100000010011100001100000000101000000000000;
			// PEs: 10, 13 -> 14
			// srcs: (1922, 34)(3140) 47, (422) 1 --> (3559) 47:PEGB2, ND5, *, PENB
			10'd49 : rdata = 48'b000111110000010001100000101000000000000100000000;
			// PEs: 13, 12 -> 12
			// srcs: (1924, 49)(3) 1, (3558) -47 --> (4342) -47:NM0, PENB, *, PEGB4
			10'd50 : rdata = 48'b000111000000000011011111110000000000000011000000;
			// PEs: 13, 14 -> 13
			// srcs: (1931, 64)(1207) 1, (4343) 47 --> (5127) -46:NW5, PEGB6, -, NW5
			10'd51 : rdata = 48'b000100100000010111100001100000000101010000000000;
			// PEs: 10, 13 -> 
			// srcs: (1963, 35)(3140) 47, (463) 1 --> (3600) 47:PEGB2, ND12, *, 
			10'd52 : rdata = 48'b000111110000010001100001100000000000000000000000;
			// PEs: 13, 13 -> 
			// srcs: (1966, 50)(3) 1, (3600) 47 --> (4384) 47:NM0, ALU, *, 
			10'd53 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 13, 13 -> 13
			// srcs: (1969, 65)(1248) 0, (4384) 47 --> (5168) -47:NW12, ALU, -, NW12
			10'd54 : rdata = 48'b000100100000110000111111111000000111000000000000;
			// PEs: 10, 13 -> 13
			// srcs: (2002, 36)(3140) 47, (502) -1 --> (3639) -47:PEGB2, ND6, *, NI0
			10'd55 : rdata = 48'b000111110000010001100000110100000000000000000000;
			// PEs: 13, 12 -> 12
			// srcs: (2004, 51)(3) 1, (3638) 94 --> (4422) 94:NM0, PENB, *, PEGB4
			10'd56 : rdata = 48'b000111000000000011011111110000000000000011000000;
			// PEs: 13, 13 -> 
			// srcs: (2005, 52)(3) 1, (3639) -47 --> (4423) -47:NM0, NI0, *, 
			10'd57 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 13, 13 -> 13
			// srcs: (2008, 66)(1287) -2, (4423) -47 --> (5207) 45:NW6, ALU, -, NW6
			10'd58 : rdata = 48'b000100100000011000111111111000000101100000000000;
			// PEs: 10, 13 -> 
			// srcs: (2084, 37)(3140) 47, (584) 2 --> (3721) 94:PEGB2, ND7, *, 
			10'd59 : rdata = 48'b000111110000010001100000111000000000000000000000;
			// PEs: 13, 13 -> 
			// srcs: (2087, 53)(3) 1, (3721) 94 --> (4505) 94:NM0, ALU, *, 
			10'd60 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 13, 13 -> 13
			// srcs: (2090, 67)(1369) 2, (4505) 94 --> (5289) -92:NW7, ALU, -, NW7
			10'd61 : rdata = 48'b000100100000011100111111111000000101110000000000;
			// PEs: 13, 12 -> 12
			// srcs: (2143, 54)(3) 1, (3777) 47 --> (4561) 47:NM0, PENB, *, PEGB4
			10'd62 : rdata = 48'b000111000000000011011111110000000000000011000000;
			// PEs: 10, 13 -> 
			// srcs: (2147, 38)(3140) 47, (647) 1 --> (3784) 47:PEGB2, ND13, *, 
			10'd63 : rdata = 48'b000111110000010001100001101000000000000000000000;
			// PEs: 13, 13 -> 
			// srcs: (2150, 55)(3) 1, (3784) 47 --> (4568) 47:NM0, ALU, *, 
			10'd64 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 13, 13 -> 13
			// srcs: (2153, 68)(1432) -3, (4568) 47 --> (5352) -50:NW13, ALU, -, NW13
			10'd65 : rdata = 48'b000100100000110100111111111000000111010000000000;
			// PEs: 10, 13 -> 14
			// srcs: (2164, 39)(3140) 47, (664) 1 --> (3801) 47:PEGB2, ND8, *, PENB
			10'd66 : rdata = 48'b000111110000010001100001000000000000000100000000;
			// PEs: 13, 14 -> 13
			// srcs: (2173, 69)(1449) 0, (4585) 47 --> (5369) -47:NW8, PEGB6, -, NW8
			10'd67 : rdata = 48'b000100100000100011100001100000000110000000000000;
			// PEs: 10, 13 -> 14
			// srcs: (2244, 40)(3140) 47, (744) 0 --> (3881) 0:PEGB2, ND9, *, PENB
			10'd68 : rdata = 48'b000111110000010001100001001000000000000100000000;
			// PEs: 13, 12 -> 12
			// srcs: (2246, 56)(3) 1, (3880) -141 --> (4664) -141:NM0, PENB, *, PEGB4
			10'd69 : rdata = 48'b000111000000000011011111110000000000000011000000;
			// PEs: 13, 14 -> 13
			// srcs: (2253, 70)(1529) 2, (4665) 0 --> (5449) 2:NW9, PEGB6, -, NW9
			10'd70 : rdata = 48'b000100100000100111100001100000000110010000000000;
			default : rdata = 48'b000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 14) begin
	always @(*) begin
		case(address)
			// PEs: 14, 14 -> 8
			// srcs: (1, 0)(20) -2, (805) -3 --> (1589) 6:ND0, NW0, *, PEGB0
			10'd0 : rdata = 48'b000110110000000001000000000000000000000010000000;
			// PEs: 14, 14 -> 14
			// srcs: (2, 1)(102) 2, (887) 1 --> (1671) 2:ND1, NW1, *, NI0
			10'd1 : rdata = 48'b000110110000000101000000001100000000000000000000;
			// PEs: 14, 14 -> 8
			// srcs: (3, 2)(182) -3, (967) 0 --> (1751) 0:ND2, NW2, *, PEGB0
			10'd2 : rdata = 48'b000110110000001001000000010000000000000010000000;
			// PEs: 14, 14 -> 8
			// srcs: (4, 3)(262) 1, (1047) -3 --> (1831) -3:ND3, NW3, *, PEGB0
			10'd3 : rdata = 48'b000110110000001101000000011000000000000010000000;
			// PEs: 14, 14 -> 8
			// srcs: (5, 4)(344) -2, (1129) -1 --> (1913) 2:ND4, NW4, *, PEGB0
			10'd4 : rdata = 48'b000110110000010001000000100000000000000010000000;
			// PEs: 14, 14 -> 8
			// srcs: (6, 5)(424) 0, (1209) 0 --> (1993) 0:ND5, NW5, *, PEGB0
			10'd5 : rdata = 48'b000110110000010101000000101000000000000010000000;
			// PEs: 14, 14 -> 8
			// srcs: (7, 6)(504) 1, (1289) 2 --> (2073) 2:ND6, NW6, *, PEGB0
			10'd6 : rdata = 48'b000110110000011001000000110000000000000010000000;
			// PEs: 14, 14 -> 8
			// srcs: (8, 7)(586) 1, (1371) 2 --> (2155) 2:ND7, NW7, *, PEGB0
			10'd7 : rdata = 48'b000110110000011101000000111000000000000010000000;
			// PEs: 14, 14 -> 12
			// srcs: (9, 8)(666) -1, (1451) -1 --> (2235) 1:ND8, NW8, *, PEGB4
			10'd8 : rdata = 48'b000110110000100001000001000000000000000011000000;
			// PEs: 14, 14 -> 13
			// srcs: (10, 9)(746) 1, (1531) 1 --> (2315) 1:ND9, NW9, *, PEGB5
			10'd9 : rdata = 48'b000110110000100101000001001000000000000011010000;
			// PEs: 14, 14 -> 14
			// srcs: (11, 10)(98) 2, (883) 2 --> (1667) 4:ND10, NW10, *, NI1
			10'd10 : rdata = 48'b000110110000101001000001010100001000000000000000;
			// PEs: 14, 14 -> 14
			// srcs: (12, 11)(282) 2, (1067) 0 --> (1851) 0:ND11, NW11, *, NI2
			10'd11 : rdata = 48'b000110110000101101000001011100010000000000000000;
			// PEs: 14, 14 -> 14
			// srcs: (13, 12)(466) -1, (1251) 1 --> (2035) -1:ND12, NW12, *, NI3
			10'd12 : rdata = 48'b000110110000110001000001100100011000000000000000;
			// PEs: 14, 14 -> 14
			// srcs: (14, 13)(650) 0, (1435) 2 --> (2219) 0:ND13, NW13, *, NI4
			10'd13 : rdata = 48'b000110110000110101000001101100100000000000000000;
			// PEs: 12, 13 -> 14
			// srcs: (16, 18)(2312) 0, (2313) 0 --> (3091) 0:PEGB4, PENB, +, NI5
			10'd14 : rdata = 48'b000011110000100011011111110100101000000000000000;
			// PEs: 8 -> 
			// srcs: (27, 14)(1611) -2 --> (1611) -2:PEGB0, pass, 
			10'd15 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 8, 14 -> 8
			// srcs: (36, 15)(1610) -6, (1611) -2 --> (2392) -8:PEGB0, ALU, +, PEGB0
			10'd16 : rdata = 48'b000011110000000000111111111000000000000010000000;
			// PEs: 8 -> 
			// srcs: (91, 16)(1904) -2 --> (1904) -2:PEGB0, pass, 
			10'd17 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 14, 9 -> 9
			// srcs: (93, 17)(1904) -2, (1905) 0 --> (2684) -2:ALU, PEGB1, +, PEGB1
			10'd18 : rdata = 48'b000010011111111111100000010000000000000010010000;
			// PEs: 14 -> 8
			// srcs: (113, 19)(1671) 2 --> (1671) 2:NI0, pass, PEGB0
			10'd19 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 14 -> 8
			// srcs: (124, 23)(1851) 0 --> (1851) 0:NI2, pass, PEGB0
			10'd20 : rdata = 48'b110001010000001000000000000000000000000010000000;
			// PEs: 14 -> 8
			// srcs: (153, 24)(2035) -1 --> (2035) -1:NI3, pass, PEGB0
			10'd21 : rdata = 48'b110001010000001100000000000000000000000010000000;
			// PEs: 14 -> 8
			// srcs: (232, 22)(1667) 4 --> (1667) 4:NI1, pass, PEGB0
			10'd22 : rdata = 48'b110001010000000100000000000000000000000010000000;
			// PEs: 8 -> 
			// srcs: (322, 20)(2065) 0 --> (2065) 0:PEGB0, pass, 
			10'd23 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 14, 9 -> 10
			// srcs: (324, 21)(2065) 0, (2066) 0 --> (2846) 0:ALU, PEGB1, +, PEGB2
			10'd24 : rdata = 48'b000010011111111111100000010000000000000010100000;
			// PEs: 14 -> 9
			// srcs: (498, 25)(2219) 0 --> (2219) 0:NI4, pass, PEGB1
			10'd25 : rdata = 48'b110001010000010000000000000000000000000010010000;
			// PEs: 14 -> 9
			// srcs: (526, 26)(3091) 0 --> (3091) 0:NI5, pass, PEGB1
			10'd26 : rdata = 48'b110001010000010100000000000000000000000010010000;
			// PEs: 10, 14 -> 
			// srcs: (1520, 27)(3140) 47, (20) -2 --> (3157) -94:PEGB2, ND0, *, 
			10'd27 : rdata = 48'b000111110000010001100000000000000000000000000000;
			// PEs: 14, 14 -> 
			// srcs: (1523, 41)(3) 1, (3157) -94 --> (3941) -94:NM0, ALU, *, 
			10'd28 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 14, 14 -> 14
			// srcs: (1526, 58)(805) -3, (3941) -94 --> (4725) 91:NW0, ALU, -, NW0
			10'd29 : rdata = 48'b000100100000000000111111111000000100000000000000;
			// PEs: 10, 14 -> 
			// srcs: (1598, 28)(3140) 47, (98) 2 --> (3235) 94:PEGB2, ND10, *, 
			10'd30 : rdata = 48'b000111110000010001100001010000000000000000000000;
			// PEs: 14, 14 -> 14
			// srcs: (1601, 42)(3) 1, (3235) 94 --> (4019) 94:NM0, ALU, *, NI0
			10'd31 : rdata = 48'b000111000000000000111111111100000000000000000000;
			// PEs: 10, 14 -> 15
			// srcs: (1602, 29)(3140) 47, (102) 2 --> (3239) 94:PEGB2, ND1, *, PENB
			10'd32 : rdata = 48'b000111110000010001100000001000000000000100000000;
			// PEs: 14, 13 -> 13
			// srcs: (1603, 43)(3) 1, (3237) 0 --> (4021) 0:NM0, PENB, *, PEGB5
			10'd33 : rdata = 48'b000111000000000011011111110000000000000011010000;
			// PEs: 14, 14 -> 14
			// srcs: (1604, 59)(883) 2, (4019) 94 --> (4803) -92:NW10, NI0, -, NW10
			10'd34 : rdata = 48'b000100100000101010100000000000000110100000000000;
			// PEs: 14, 15 -> 14
			// srcs: (1611, 60)(887) 1, (4023) 94 --> (4807) -93:NW1, PEGB7, -, NW1
			10'd35 : rdata = 48'b000100100000000111100001110000000100010000000000;
			// PEs: 10, 14 -> 14
			// srcs: (1682, 30)(3140) 47, (182) -3 --> (3319) -141:PEGB2, ND2, *, NI0
			10'd36 : rdata = 48'b000111110000010001100000010100000000000000000000;
			// PEs: 14, 13 -> 13
			// srcs: (1683, 44)(3) 1, (3317) 47 --> (4101) 47:NM0, PENB, *, PEGB5
			10'd37 : rdata = 48'b000111000000000011011111110000000000000011010000;
			// PEs: 14, 14 -> 
			// srcs: (1685, 45)(3) 1, (3319) -141 --> (4103) -141:NM0, NI0, *, 
			10'd38 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 14, 14 -> 14
			// srcs: (1688, 61)(967) 0, (4103) -141 --> (4887) 141:NW2, ALU, -, NW2
			10'd39 : rdata = 48'b000100100000001000111111111000000100100000000000;
			// PEs: 10, 14 -> 
			// srcs: (1762, 31)(3140) 47, (262) 1 --> (3399) 47:PEGB2, ND3, *, 
			10'd40 : rdata = 48'b000111110000010001100000011000000000000000000000;
			// PEs: 14, 14 -> 
			// srcs: (1765, 46)(3) 1, (3399) 47 --> (4183) 47:NM0, ALU, *, 
			10'd41 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 14, 14 -> 14
			// srcs: (1768, 62)(1047) -3, (4183) 47 --> (4967) -50:NW3, ALU, -, NW3
			10'd42 : rdata = 48'b000100100000001100111111111000000100110000000000;
			// PEs: 10, 14 -> 
			// srcs: (1782, 32)(3140) 47, (282) 2 --> (3419) 94:PEGB2, ND11, *, 
			10'd43 : rdata = 48'b000111110000010001100001011000000000000000000000;
			// PEs: 14, 14 -> 
			// srcs: (1785, 47)(3) 1, (3419) 94 --> (4203) 94:NM0, ALU, *, 
			10'd44 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 14, 14 -> 14
			// srcs: (1788, 63)(1067) 0, (4203) 94 --> (4987) -94:NW11, ALU, -, NW11
			10'd45 : rdata = 48'b000100100000101100111111111000000110110000000000;
			// PEs: 10, 14 -> 15
			// srcs: (1844, 33)(3140) 47, (344) -2 --> (3481) -94:PEGB2, ND4, *, PENB
			10'd46 : rdata = 48'b000111110000010001100000100000000000000100000000;
			// PEs: 14, 13 -> 13
			// srcs: (1845, 48)(3) 1, (3479) -141 --> (4263) -141:NM0, PENB, *, PEGB5
			10'd47 : rdata = 48'b000111000000000011011111110000000000000011010000;
			// PEs: 14, 15 -> 14
			// srcs: (1853, 64)(1129) -1, (4265) -94 --> (5049) 93:NW4, PEGB7, -, NW4
			10'd48 : rdata = 48'b000100100000010011100001110000000101000000000000;
			// PEs: 10, 14 -> 14
			// srcs: (1924, 34)(3140) 47, (424) 0 --> (3561) 0:PEGB2, ND5, *, NI0
			10'd49 : rdata = 48'b000111110000010001100000101100000000000000000000;
			// PEs: 14, 13 -> 13
			// srcs: (1925, 49)(3) 1, (3559) 47 --> (4343) 47:NM0, PENB, *, PEGB5
			10'd50 : rdata = 48'b000111000000000011011111110000000000000011010000;
			// PEs: 14, 14 -> 
			// srcs: (1927, 50)(3) 1, (3561) 0 --> (4345) 0:NM0, NI0, *, 
			10'd51 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 14, 14 -> 14
			// srcs: (1930, 65)(1209) 0, (4345) 0 --> (5129) 0:NW5, ALU, -, NW5
			10'd52 : rdata = 48'b000100100000010100111111111000000101010000000000;
			// PEs: 10, 14 -> 
			// srcs: (1966, 35)(3140) 47, (466) -1 --> (3603) -47:PEGB2, ND12, *, 
			10'd53 : rdata = 48'b000111110000010001100001100000000000000000000000;
			// PEs: 14, 14 -> 
			// srcs: (1969, 51)(3) 1, (3603) -47 --> (4387) -47:NM0, ALU, *, 
			10'd54 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 14, 14 -> 14
			// srcs: (1972, 66)(1251) 1, (4387) -47 --> (5171) 48:NW12, ALU, -, NW12
			10'd55 : rdata = 48'b000100100000110000111111111000000111000000000000;
			// PEs: 10, 14 -> 
			// srcs: (2004, 36)(3140) 47, (504) 1 --> (3641) 47:PEGB2, ND6, *, 
			10'd56 : rdata = 48'b000111110000010001100000110000000000000000000000;
			// PEs: 14, 14 -> 
			// srcs: (2007, 52)(3) 1, (3641) 47 --> (4425) 47:NM0, ALU, *, 
			10'd57 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 14, 14 -> 14
			// srcs: (2010, 67)(1289) 2, (4425) 47 --> (5209) -45:NW6, ALU, -, NW6
			10'd58 : rdata = 48'b000100100000011000111111111000000101100000000000;
			// PEs: 10, 14 -> 
			// srcs: (2086, 37)(3140) 47, (586) 1 --> (3723) 47:PEGB2, ND7, *, 
			10'd59 : rdata = 48'b000111110000010001100000111000000000000000000000;
			// PEs: 14, 14 -> 
			// srcs: (2089, 53)(3) 1, (3723) 47 --> (4507) 47:NM0, ALU, *, 
			10'd60 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 14, 14 -> 14
			// srcs: (2092, 68)(1371) 2, (4507) 47 --> (5291) -45:NW7, ALU, -, NW7
			10'd61 : rdata = 48'b000100100000011100111111111000000101110000000000;
			// PEs: 10, 14 -> 
			// srcs: (2150, 38)(3140) 47, (650) 0 --> (3787) 0:PEGB2, ND13, *, 
			10'd62 : rdata = 48'b000111110000010001100001101000000000000000000000;
			// PEs: 14, 14 -> 
			// srcs: (2153, 54)(3) 1, (3787) 0 --> (4571) 0:NM0, ALU, *, 
			10'd63 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 14, 14 -> 14
			// srcs: (2156, 69)(1435) 2, (4571) 0 --> (5355) 2:NW13, ALU, -, NW13
			10'd64 : rdata = 48'b000100100000110100111111111000000111010000000000;
			// PEs: 10, 14 -> 15
			// srcs: (2166, 39)(3140) 47, (666) -1 --> (3803) -47:PEGB2, ND8, *, PENB
			10'd65 : rdata = 48'b000111110000010001100001000000000000000100000000;
			// PEs: 14, 13 -> 13
			// srcs: (2167, 55)(3) 1, (3801) 47 --> (4585) 47:NM0, PENB, *, PEGB5
			10'd66 : rdata = 48'b000111000000000011011111110000000000000011010000;
			// PEs: 14, 15 -> 14
			// srcs: (2175, 70)(1451) -1, (4587) -47 --> (5371) 46:NW8, PEGB7, -, NW8
			10'd67 : rdata = 48'b000100100000100011100001110000000110000000000000;
			// PEs: 10, 14 -> 14
			// srcs: (2246, 40)(3140) 47, (746) 1 --> (3883) 47:PEGB2, ND9, *, NI0
			10'd68 : rdata = 48'b000111110000010001100001001100000000000000000000;
			// PEs: 14, 13 -> 13
			// srcs: (2247, 56)(3) 1, (3881) 0 --> (4665) 0:NM0, PENB, *, PEGB5
			10'd69 : rdata = 48'b000111000000000011011111110000000000000011010000;
			// PEs: 14, 14 -> 
			// srcs: (2249, 57)(3) 1, (3883) 47 --> (4667) 47:NM0, NI0, *, 
			10'd70 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 14, 14 -> 14
			// srcs: (2252, 71)(1531) 1, (4667) 47 --> (5451) -46:NW9, ALU, -, NW9
			10'd71 : rdata = 48'b000100100000100100111111111000000110010000000000;
			default : rdata = 48'b000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 15) begin
	always @(*) begin
		case(address)
			// PEs: 15, 15 -> 8
			// srcs: (1, 0)(21) -1, (806) -3 --> (1590) 3:ND0, NW0, *, PENB
			10'd0 : rdata = 48'b000110110000000001000000000000000000000100000000;
			// PEs: 15, 15 -> 15
			// srcs: (2, 1)(103) -1, (888) -1 --> (1672) 1:ND1, NW1, *, NI0
			10'd1 : rdata = 48'b000110110000000101000000001100000000000000000000;
			// PEs: 15, 15 -> 8
			// srcs: (3, 2)(183) 1, (968) 2 --> (1752) 2:ND2, NW2, *, PENB
			10'd2 : rdata = 48'b000110110000001001000000010000000000000100000000;
			// PEs: 15, 15 -> 8
			// srcs: (4, 3)(263) -3, (1048) -3 --> (1832) 9:ND3, NW3, *, PENB
			10'd3 : rdata = 48'b000110110000001101000000011000000000000100000000;
			// PEs: 15, 15 -> 8
			// srcs: (5, 4)(345) 2, (1130) -2 --> (1914) -4:ND4, NW4, *, PENB
			10'd4 : rdata = 48'b000110110000010001000000100000000000000100000000;
			// PEs: 15, 15 -> 8
			// srcs: (6, 5)(425) -3, (1210) 0 --> (1994) 0:ND5, NW5, *, PENB
			10'd5 : rdata = 48'b000110110000010101000000101000000000000100000000;
			// PEs: 15, 15 -> 8
			// srcs: (7, 6)(505) -2, (1290) -2 --> (2074) 4:ND6, NW6, *, PENB
			10'd6 : rdata = 48'b000110110000011001000000110000000000000100000000;
			// PEs: 15, 15 -> 8
			// srcs: (8, 7)(587) -2, (1372) -1 --> (2156) 2:ND7, NW7, *, PENB
			10'd7 : rdata = 48'b000110110000011101000000111000000000000100000000;
			// PEs: 15, 15 -> 12
			// srcs: (9, 8)(667) -2, (1452) 2 --> (2236) -4:ND8, NW8, *, PEGB4
			10'd8 : rdata = 48'b000110110000100001000001000000000000000011000000;
			// PEs: 15, 15 -> 13
			// srcs: (10, 9)(747) 2, (1532) -2 --> (2316) -4:ND9, NW9, *, PEGB5
			10'd9 : rdata = 48'b000110110000100101000001001000000000000011010000;
			// PEs: 15, 15 -> 15
			// srcs: (11, 10)(101) -3, (886) 2 --> (1670) -6:ND10, NW10, *, NI1
			10'd10 : rdata = 48'b000110110000101001000001010100001000000000000000;
			// PEs: 15, 15 -> 15
			// srcs: (12, 11)(285) 0, (1070) -1 --> (1854) 0:ND11, NW11, *, NI2
			10'd11 : rdata = 48'b000110110000101101000001011100010000000000000000;
			// PEs: 15, 15 -> 15
			// srcs: (13, 12)(469) -2, (1254) 1 --> (2038) -2:ND12, NW12, *, NI3
			10'd12 : rdata = 48'b000110110000110001000001100100011000000000000000;
			// PEs: 15, 15 -> 9
			// srcs: (14, 13)(653) 2, (1438) -2 --> (2222) -4:ND13, NW13, *, PEGB1
			10'd13 : rdata = 48'b000110110000110101000001101000000000000010010000;
			// PEs: 8 -> 
			// srcs: (29, 14)(1614) 6 --> (1614) 6:PEGB0, pass, 
			10'd14 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 8, 15 -> 8
			// srcs: (38, 15)(1613) 0, (1614) 6 --> (2394) 6:PEGB0, ALU, +, PENB
			10'd15 : rdata = 48'b000011110000000000111111111000000000000100000000;
			// PEs: 8 -> 
			// srcs: (115, 16)(1984) -3 --> (1984) -3:PEGB0, pass, 
			10'd16 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 15, 9 -> 15
			// srcs: (117, 17)(1984) -3, (1985) -1 --> (2765) -4:ALU, PEGB1, +, NI4
			10'd17 : rdata = 48'b000010011111111111100000010100100000000000000000;
			// PEs: 15 -> 8
			// srcs: (121, 20)(1672) 1 --> (1672) 1:NI0, pass, PENB
			10'd18 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 15 -> 8
			// srcs: (131, 21)(1670) -6 --> (1670) -6:NI1, pass, PENB
			10'd19 : rdata = 48'b110001010000000100000000000000000000000100000000;
			// PEs: 15 -> 8
			// srcs: (140, 22)(1854) 0 --> (1854) 0:NI2, pass, PENB
			10'd20 : rdata = 48'b110001010000001000000000000000000000000100000000;
			// PEs: 15 -> 8
			// srcs: (148, 23)(2765) -4 --> (2765) -4:NI4, pass, PENB
			10'd21 : rdata = 48'b110001010000010000000000000000000000000100000000;
			// PEs: 8 -> 
			// srcs: (218, 18)(1625) 4 --> (1625) 4:PEGB0, pass, 
			10'd22 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 8, 15 -> 8
			// srcs: (227, 19)(1624) 0, (1625) 4 --> (2406) 4:PEGB0, ALU, +, PENB
			10'd23 : rdata = 48'b000011110000000000111111111000000000000100000000;
			// PEs: 15 -> 8
			// srcs: (260, 24)(2038) -2 --> (2038) -2:NI3, pass, PENB
			10'd24 : rdata = 48'b110001010000001100000000000000000000000100000000;
			// PEs: 9 -> 
			// srcs: (536, 25)(3092) 4 --> (3092) 4:PEGB1, pass, 
			10'd25 : rdata = 48'b110001110000001000000000000000000000000000000000;
			// PEs: 13, 15 -> 9
			// srcs: (539, 26)(3090) 12, (3092) 4 --> (3093) 16:PEGB5, ALU, +, PEGB1
			10'd26 : rdata = 48'b000011110000101000111111111000000000000010010000;
			// PEs: 10, 15 -> 
			// srcs: (1521, 27)(3140) 47, (21) -1 --> (3158) -47:PEGB2, ND0, *, 
			10'd27 : rdata = 48'b000111110000010001100000000000000000000000000000;
			// PEs: 15, 15 -> 
			// srcs: (1524, 41)(3) 1, (3158) -47 --> (3942) -47:NM0, ALU, *, 
			10'd28 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 15, 15 -> 15
			// srcs: (1527, 58)(806) -3, (3942) -47 --> (4726) 44:NW0, ALU, -, NW0
			10'd29 : rdata = 48'b000100100000000000111111111000000100000000000000;
			// PEs: 10, 15 -> 15
			// srcs: (1601, 28)(3140) 47, (101) -3 --> (3238) -141:PEGB2, ND10, *, NI0
			10'd30 : rdata = 48'b000111110000010001100001010100000000000000000000;
			// PEs: 10, 15 -> 15
			// srcs: (1603, 29)(3140) 47, (103) -1 --> (3240) -47:PEGB2, ND1, *, NI1
			10'd31 : rdata = 48'b000111110000010001100000001100001000000000000000;
			// PEs: 15, 15 -> 15
			// srcs: (1604, 42)(3) 1, (3238) -141 --> (4022) -141:NM0, NI0, *, NI2
			10'd32 : rdata = 48'b000111000000000010100000000100010000000000000000;
			// PEs: 15, 14 -> 14
			// srcs: (1605, 43)(3) 1, (3239) 94 --> (4023) 94:NM0, PENB, *, PEGB6
			10'd33 : rdata = 48'b000111000000000011011111110000000000000011100000;
			// PEs: 15, 15 -> 15
			// srcs: (1606, 44)(3) 1, (3240) -47 --> (4024) -47:NM0, NI1, *, NI0
			10'd34 : rdata = 48'b000111000000000010100000001100000000000000000000;
			// PEs: 15, 15 -> 15
			// srcs: (1607, 59)(886) 2, (4022) -141 --> (4806) 143:NW10, NI2, -, NW10
			10'd35 : rdata = 48'b000100100000101010100000010000000110100000000000;
			// PEs: 15, 15 -> 15
			// srcs: (1609, 60)(888) -1, (4024) -47 --> (4808) 46:NW1, NI0, -, NW1
			10'd36 : rdata = 48'b000100100000000110100000000000000100010000000000;
			// PEs: 10, 15 -> 
			// srcs: (1683, 30)(3140) 47, (183) 1 --> (3320) 47:PEGB2, ND2, *, 
			10'd37 : rdata = 48'b000111110000010001100000010000000000000000000000;
			// PEs: 15, 15 -> 
			// srcs: (1686, 45)(3) 1, (3320) 47 --> (4104) 47:NM0, ALU, *, 
			10'd38 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 15, 15 -> 15
			// srcs: (1689, 61)(968) 2, (4104) 47 --> (4888) -45:NW2, ALU, -, NW2
			10'd39 : rdata = 48'b000100100000001000111111111000000100100000000000;
			// PEs: 10, 15 -> 
			// srcs: (1763, 31)(3140) 47, (263) -3 --> (3400) -141:PEGB2, ND3, *, 
			10'd40 : rdata = 48'b000111110000010001100000011000000000000000000000;
			// PEs: 15, 15 -> 
			// srcs: (1766, 46)(3) 1, (3400) -141 --> (4184) -141:NM0, ALU, *, 
			10'd41 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 15, 15 -> 15
			// srcs: (1769, 62)(1048) -3, (4184) -141 --> (4968) 138:NW3, ALU, -, NW3
			10'd42 : rdata = 48'b000100100000001100111111111000000100110000000000;
			// PEs: 10, 15 -> 
			// srcs: (1785, 32)(3140) 47, (285) 0 --> (3422) 0:PEGB2, ND11, *, 
			10'd43 : rdata = 48'b000111110000010001100001011000000000000000000000;
			// PEs: 15, 15 -> 
			// srcs: (1788, 47)(3) 1, (3422) 0 --> (4206) 0:NM0, ALU, *, 
			10'd44 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 15, 15 -> 15
			// srcs: (1791, 63)(1070) -1, (4206) 0 --> (4990) -1:NW11, ALU, -, NW11
			10'd45 : rdata = 48'b000100100000101100111111111000000110110000000000;
			// PEs: 10, 15 -> 15
			// srcs: (1845, 33)(3140) 47, (345) 2 --> (3482) 94:PEGB2, ND4, *, NI0
			10'd46 : rdata = 48'b000111110000010001100000100100000000000000000000;
			// PEs: 15, 14 -> 14
			// srcs: (1847, 48)(3) 1, (3481) -94 --> (4265) -94:NM0, PENB, *, PEGB6
			10'd47 : rdata = 48'b000111000000000011011111110000000000000011100000;
			// PEs: 15, 15 -> 
			// srcs: (1848, 49)(3) 1, (3482) 94 --> (4266) 94:NM0, NI0, *, 
			10'd48 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 15, 15 -> 15
			// srcs: (1851, 64)(1130) -2, (4266) 94 --> (5050) -96:NW4, ALU, -, NW4
			10'd49 : rdata = 48'b000100100000010000111111111000000101000000000000;
			// PEs: 10, 15 -> 
			// srcs: (1925, 34)(3140) 47, (425) -3 --> (3562) -141:PEGB2, ND5, *, 
			10'd50 : rdata = 48'b000111110000010001100000101000000000000000000000;
			// PEs: 15, 15 -> 
			// srcs: (1928, 50)(3) 1, (3562) -141 --> (4346) -141:NM0, ALU, *, 
			10'd51 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 15, 15 -> 15
			// srcs: (1931, 65)(1210) 0, (4346) -141 --> (5130) 141:NW5, ALU, -, NW5
			10'd52 : rdata = 48'b000100100000010100111111111000000101010000000000;
			// PEs: 10, 15 -> 
			// srcs: (1969, 35)(3140) 47, (469) -2 --> (3606) -94:PEGB2, ND12, *, 
			10'd53 : rdata = 48'b000111110000010001100001100000000000000000000000;
			// PEs: 15, 15 -> 
			// srcs: (1972, 51)(3) 1, (3606) -94 --> (4390) -94:NM0, ALU, *, 
			10'd54 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 15, 15 -> 15
			// srcs: (1975, 66)(1254) 1, (4390) -94 --> (5174) 95:NW12, ALU, -, NW12
			10'd55 : rdata = 48'b000100100000110000111111111000000111000000000000;
			// PEs: 10, 15 -> 
			// srcs: (2005, 36)(3140) 47, (505) -2 --> (3642) -94:PEGB2, ND6, *, 
			10'd56 : rdata = 48'b000111110000010001100000110000000000000000000000;
			// PEs: 15, 15 -> 
			// srcs: (2008, 52)(3) 1, (3642) -94 --> (4426) -94:NM0, ALU, *, 
			10'd57 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 15, 15 -> 15
			// srcs: (2011, 67)(1290) -2, (4426) -94 --> (5210) 92:NW6, ALU, -, NW6
			10'd58 : rdata = 48'b000100100000011000111111111000000101100000000000;
			// PEs: 10, 15 -> 
			// srcs: (2087, 37)(3140) 47, (587) -2 --> (3724) -94:PEGB2, ND7, *, 
			10'd59 : rdata = 48'b000111110000010001100000111000000000000000000000;
			// PEs: 15, 15 -> 
			// srcs: (2090, 53)(3) 1, (3724) -94 --> (4508) -94:NM0, ALU, *, 
			10'd60 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 15, 15 -> 15
			// srcs: (2093, 68)(1372) -1, (4508) -94 --> (5292) 93:NW7, ALU, -, NW7
			10'd61 : rdata = 48'b000100100000011100111111111000000101110000000000;
			// PEs: 10, 15 -> 
			// srcs: (2153, 38)(3140) 47, (653) 2 --> (3790) 94:PEGB2, ND13, *, 
			10'd62 : rdata = 48'b000111110000010001100001101000000000000000000000;
			// PEs: 15, 15 -> 
			// srcs: (2156, 54)(3) 1, (3790) 94 --> (4574) 94:NM0, ALU, *, 
			10'd63 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 15, 15 -> 15
			// srcs: (2159, 69)(1438) -2, (4574) 94 --> (5358) -96:NW13, ALU, -, NW13
			10'd64 : rdata = 48'b000100100000110100111111111000000111010000000000;
			// PEs: 10, 15 -> 15
			// srcs: (2167, 39)(3140) 47, (667) -2 --> (3804) -94:PEGB2, ND8, *, NI0
			10'd65 : rdata = 48'b000111110000010001100001000100000000000000000000;
			// PEs: 15, 14 -> 14
			// srcs: (2169, 55)(3) 1, (3803) -47 --> (4587) -47:NM0, PENB, *, PEGB6
			10'd66 : rdata = 48'b000111000000000011011111110000000000000011100000;
			// PEs: 15, 15 -> 
			// srcs: (2170, 56)(3) 1, (3804) -94 --> (4588) -94:NM0, NI0, *, 
			10'd67 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 15, 15 -> 15
			// srcs: (2173, 70)(1452) 2, (4588) -94 --> (5372) 96:NW8, ALU, -, NW8
			10'd68 : rdata = 48'b000100100000100000111111111000000110000000000000;
			// PEs: 10, 15 -> 
			// srcs: (2247, 40)(3140) 47, (747) 2 --> (3884) 94:PEGB2, ND9, *, 
			10'd69 : rdata = 48'b000111110000010001100001001000000000000000000000;
			// PEs: 15, 15 -> 
			// srcs: (2250, 57)(3) 1, (3884) 94 --> (4668) 94:NM0, ALU, *, 
			10'd70 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 15, 15 -> 15
			// srcs: (2253, 71)(1532) -2, (4668) 94 --> (5452) -96:NW9, ALU, -, NW9
			10'd71 : rdata = 48'b000100100000100100111111111000000110010000000000;
			default : rdata = 48'b000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 16) begin
	always @(*) begin
		case(address)
			// PEs: 17 -> 0
			// srcs: (6, 3)(1592) 9 --> (1592) 9:PEGB1, pass, PUGB0
			10'd0 : rdata = 48'b110001110000001000000000000000000000000000001000;
			// PEs: 18 -> 0
			// srcs: (7, 4)(1593) -3 --> (1593) -3:PEGB2, pass, PUGB0
			10'd1 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 19 -> 0
			// srcs: (8, 5)(1595) 0 --> (1595) 0:PEGB3, pass, PUGB0
			10'd2 : rdata = 48'b110001110000011000000000000000000000000000001000;
			// PEs: 20 -> 0
			// srcs: (9, 6)(1596) -6 --> (1596) -6:PEGB4, pass, PUGB0
			10'd3 : rdata = 48'b110001110000100000000000000000000000000000001000;
			// PEs: 21 -> 8
			// srcs: (10, 7)(1598) 4 --> (1598) 4:PEGB5, pass, PUGB1
			10'd4 : rdata = 48'b110001110000101000000000000000000000000000001001;
			// PEs: 0 -> 16
			// srcs: (11, 0)(1577) -4 --> (1577) -4:PUGB0, pass, NI0
			10'd5 : rdata = 48'b110001110000000100000000000100000000000000000000;
			// PEs: 0 -> 18
			// srcs: (12, 1)(1578) -6 --> (1578) -6:PUGB0, pass, PEGB2
			10'd6 : rdata = 48'b110001110000000100000000000000000000000010100000;
			// PEs: 22 -> 8
			// srcs: (13, 8)(1599) -2 --> (1599) -2:PEGB6, pass, PUGB1
			10'd7 : rdata = 48'b110001110000110000000000000000000000000000001001;
			// PEs: 23 -> 8
			// srcs: (14, 9)(1601) 4 --> (1601) 4:PENB, pass, PUGB1
			10'd8 : rdata = 48'b110001101111111000000000000000000000000000001001;
			// PEs: 32 -> 16
			// srcs: (15, 10)(1616) 0 --> (1616) 0:PUGB4, pass, NI1
			10'd9 : rdata = 48'b110001110000100100000000000100001000000000000000;
			// PEs: 32 -> 19
			// srcs: (16, 11)(1617) -4 --> (1617) -4:PUGB4, pass, PEGB3
			10'd10 : rdata = 48'b110001110000100100000000000000000000000010110000;
			// PEs: 32 -> 16
			// srcs: (17, 13)(1619) 0 --> (1619) 0:PUGB4, pass, NI2
			10'd11 : rdata = 48'b110001110000100100000000000100010000000000000000;
			// PEs: 32 -> 20
			// srcs: (18, 14)(1620) 0 --> (1620) 0:PUGB4, pass, PEGB4
			10'd12 : rdata = 48'b110001110000100100000000000000000000000011000000;
			// PEs: 40 -> 16
			// srcs: (19, 16)(1626) 0 --> (1626) 0:PUGB5, pass, NI3
			10'd13 : rdata = 48'b110001110000101100000000000100011000000000000000;
			// PEs: 40 -> 21
			// srcs: (20, 17)(1627) 6 --> (1627) 6:PUGB5, pass, PEGB5
			10'd14 : rdata = 48'b110001110000101100000000000000000000000011010000;
			// PEs: 16 -> 18
			// srcs: (21, 2)(1577) -4 --> (1577) -4:NI0, pass, PEGB2
			10'd15 : rdata = 48'b110001010000000000000000000000000000000010100000;
			// PEs: 40 -> 16
			// srcs: (22, 19)(1629) 2 --> (1629) 2:PUGB5, pass, NI0
			10'd16 : rdata = 48'b110001110000101100000000000100000000000000000000;
			// PEs: 40 -> 22
			// srcs: (23, 20)(1630) -2 --> (1630) -2:PUGB5, pass, PEGB6
			10'd17 : rdata = 48'b110001110000101100000000000000000000000011100000;
			// PEs: 48 -> 16
			// srcs: (24, 22)(1632) 0 --> (1632) 0:PUGB6, pass, NI4
			10'd18 : rdata = 48'b110001110000110100000000000100100000000000000000;
			// PEs: 16 -> 19
			// srcs: (25, 12)(1616) 0 --> (1616) 0:NI1, pass, PEGB3
			10'd19 : rdata = 48'b110001010000000100000000000000000000000010110000;
			// PEs: 48 -> 23
			// srcs: (26, 23)(1633) -6 --> (1633) -6:PUGB6, pass, PEGB7
			10'd20 : rdata = 48'b110001110000110100000000000000000000000011110000;
			// PEs: 16 -> 20
			// srcs: (27, 15)(1619) 0 --> (1619) 0:NI2, pass, PEGB4
			10'd21 : rdata = 48'b110001010000001000000000000000000000000011000000;
			// PEs: 0 -> 16
			// srcs: (28, 25)(1653) 0 --> (1653) 0:PUGB0, pass, NI1
			10'd22 : rdata = 48'b110001110000000100000000000100001000000000000000;
			// PEs: 16 -> 21
			// srcs: (29, 18)(1626) 0 --> (1626) 0:NI3, pass, PEGB5
			10'd23 : rdata = 48'b110001010000001100000000000000000000000011010000;
			// PEs: 0 -> 17
			// srcs: (30, 26)(1654) -4 --> (1654) -4:PUGB0, pass, PENB
			10'd24 : rdata = 48'b110001110000000100000000000000000000000100000000;
			// PEs: 19 -> 8
			// srcs: (31, 28)(1675) 4 --> (1675) 4:PEGB3, pass, PUGB1
			10'd25 : rdata = 48'b110001110000011000000000000000000000000000001001;
			// PEs: 16 -> 22
			// srcs: (32, 21)(1629) 2 --> (1629) 2:NI0, pass, PEGB6
			10'd26 : rdata = 48'b110001010000000000000000000000000000000011100000;
			// PEs: 20 -> 8
			// srcs: (33, 29)(1676) -6 --> (1676) -6:PEGB4, pass, PUGB1
			10'd27 : rdata = 48'b110001110000100000000000000000000000000000001001;
			// PEs: 21 -> 56
			// srcs: (34, 30)(1678) -1 --> (1678) -1:PEGB5, pass, PUGB7
			10'd28 : rdata = 48'b110001110000101000000000000000000000000000001111;
			// PEs: 16 -> 23
			// srcs: (35, 24)(1632) 0 --> (1632) 0:NI4, pass, PEGB7
			10'd29 : rdata = 48'b110001010000010000000000000000000000000011110000;
			// PEs: 16 -> 17
			// srcs: (36, 27)(1653) 0 --> (1653) 0:NI1, pass, PENB
			10'd30 : rdata = 48'b110001010000000100000000000000000000000100000000;
			// PEs: 22 -> 56
			// srcs: (37, 31)(1679) -4 --> (1679) -4:PEGB6, pass, PUGB7
			10'd31 : rdata = 48'b110001110000110000000000000000000000000000001111;
			// PEs: 23 -> 32
			// srcs: (38, 32)(1681) 3 --> (1681) 3:PENB, pass, PUGB4
			10'd32 : rdata = 48'b110001101111111000000000000000000000000000001100;
			// PEs: 17 -> 8
			// srcs: (39, 39)(1754) 0 --> (1754) 0:PEGB1, pass, PUGB1
			10'd33 : rdata = 48'b110001110000001000000000000000000000000000001001;
			// PEs: 18 -> 8
			// srcs: (40, 40)(1755) -4 --> (1755) -4:PEGB2, pass, PUGB1
			10'd34 : rdata = 48'b110001110000010000000000000000000000000000001001;
			// PEs: 19 -> 24
			// srcs: (41, 41)(1757) -4 --> (1757) -4:PEGB3, pass, PUNB
			10'd35 : rdata = 48'b110001110000011000000000000000000000001000000000;
			// PEs: 20 -> 24
			// srcs: (42, 42)(1758) 0 --> (1758) 0:PEGB4, pass, PUNB
			10'd36 : rdata = 48'b110001110000100000000000000000000000001000000000;
			// PEs: 21 -> 24
			// srcs: (43, 43)(1760) -4 --> (1760) -4:PEGB5, pass, PUNB
			10'd37 : rdata = 48'b110001110000101000000000000000000000001000000000;
			// PEs: 22 -> 24
			// srcs: (44, 44)(1761) -1 --> (1761) -1:PEGB6, pass, PUNB
			10'd38 : rdata = 48'b110001110000110000000000000000000000001000000000;
			// PEs: 23 -> 32
			// srcs: (45, 45)(1763) 0 --> (1763) 0:PENB, pass, PUGB4
			10'd39 : rdata = 48'b110001101111111000000000000000000000000000001100;
			// PEs: 40 -> 16
			// srcs: (46, 46)(1788) 3 --> (1788) 3:PUGB5, pass, NI0
			10'd40 : rdata = 48'b110001110000101100000000000100000000000000000000;
			// PEs: 40 -> 17
			// srcs: (47, 47)(1789) 4 --> (1789) 4:PUGB5, pass, PENB
			10'd41 : rdata = 48'b110001110000101100000000000000000000000100000000;
			// PEs: 17 -> 24
			// srcs: (48, 61)(1834) 0 --> (1834) 0:PEGB1, pass, PUNB
			10'd42 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 18 -> 24
			// srcs: (49, 62)(1835) -2 --> (1835) -2:PEGB2, pass, PUNB
			10'd43 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 8 -> 16
			// srcs: (50, 33)(1748) -3 --> (1748) -3:PUNB, pass, NI1
			10'd44 : rdata = 48'b110001101111111100000000000100001000000000000000;
			// PEs: 19 -> 24
			// srcs: (51, 63)(1837) 1 --> (1837) 1:PEGB3, pass, PUNB
			10'd45 : rdata = 48'b110001110000011000000000000000000000001000000000;
			// PEs: 8 -> 18
			// srcs: (52, 34)(1749) 2 --> (1749) 2:PUNB, pass, PEGB2
			10'd46 : rdata = 48'b110001101111111100000000000000000000000010100000;
			// PEs: 16 -> 17
			// srcs: (53, 48)(1788) 3 --> (1788) 3:NI0, pass, PENB
			10'd47 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 8 -> 16
			// srcs: (54, 36)(1751) 0 --> (1751) 0:PUNB, pass, NI0
			10'd48 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 8 -> 19
			// srcs: (55, 37)(1752) 2 --> (1752) 2:PUNB, pass, PEGB3
			10'd49 : rdata = 48'b110001101111111100000000000000000000000010110000;
			// PEs: 20 -> 24
			// srcs: (56, 64)(1838) 3 --> (1838) 3:PEGB4, pass, PUNB
			10'd50 : rdata = 48'b110001110000100000000000000000000000001000000000;
			// PEs: 21 -> 24
			// srcs: (57, 65)(1840) -1 --> (1840) -1:PEGB5, pass, PUNB
			10'd51 : rdata = 48'b110001110000101000000000000000000000001000000000;
			// PEs: 22 -> 24
			// srcs: (58, 66)(1841) -1 --> (1841) -1:PEGB6, pass, PUNB
			10'd52 : rdata = 48'b110001110000110000000000000000000000001000000000;
			// PEs: 23 -> 32
			// srcs: (59, 67)(1843) 1 --> (1843) 1:PENB, pass, PUGB4
			10'd53 : rdata = 48'b110001101111111000000000000000000000000000001100;
			// PEs: 21 -> 24
			// srcs: (60, 77)(1920) 6 --> (1920) 6:PEGB5, pass, PUNB
			10'd54 : rdata = 48'b110001110000101000000000000000000000001000000000;
			// PEs: 16 -> 18
			// srcs: (61, 35)(1748) -3 --> (1748) -3:NI1, pass, PEGB2
			10'd55 : rdata = 48'b110001010000000100000000000000000000000010100000;
			// PEs: 0 -> 16
			// srcs: (62, 49)(1822) 0 --> (1822) 0:PUGB0, pass, NI1
			10'd56 : rdata = 48'b110001110000000100000000000100001000000000000000;
			// PEs: 8 -> 20
			// srcs: (63, 50)(1823) 0 --> (1823) 0:PUNB, pass, PEGB4
			10'd57 : rdata = 48'b110001101111111100000000000000000000000011000000;
			// PEs: 16 -> 19
			// srcs: (64, 38)(1751) 0 --> (1751) 0:NI0, pass, PEGB3
			10'd58 : rdata = 48'b110001010000000000000000000000000000000010110000;
			// PEs: 8 -> 16
			// srcs: (65, 52)(1825) 1 --> (1825) 1:PUNB, pass, NI0
			10'd59 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 8 -> 21
			// srcs: (66, 53)(1826) -2 --> (1826) -2:PUNB, pass, PEGB5
			10'd60 : rdata = 48'b110001101111111100000000000000000000000011010000;
			// PEs: 8 -> 16
			// srcs: (67, 55)(1828) 0 --> (1828) 0:PUNB, pass, NI2
			10'd61 : rdata = 48'b110001101111111100000000000100010000000000000000;
			// PEs: 8 -> 22
			// srcs: (68, 56)(1829) 0 --> (1829) 0:PUNB, pass, PEGB6
			10'd62 : rdata = 48'b110001101111111100000000000000000000000011100000;
			// PEs: 8 -> 16
			// srcs: (69, 58)(1831) -3 --> (1831) -3:PUNB, pass, NI3
			10'd63 : rdata = 48'b110001101111111100000000000100011000000000000000;
			// PEs: 8 -> 23
			// srcs: (70, 59)(1832) 9 --> (1832) 9:PUNB, pass, PEGB7
			10'd64 : rdata = 48'b110001101111111100000000000000000000000011110000;
			// PEs: 22 -> 24
			// srcs: (71, 78)(1921) -6 --> (1921) -6:PEGB6, pass, PUNB
			10'd65 : rdata = 48'b110001110000110000000000000000000000001000000000;
			// PEs: 16 -> 20
			// srcs: (72, 51)(1822) 0 --> (1822) 0:NI1, pass, PEGB4
			10'd66 : rdata = 48'b110001010000000100000000000000000000000011000000;
			// PEs: 8 -> 16
			// srcs: (73, 68)(1907) 0 --> (1907) 0:PUNB, pass, NI1
			10'd67 : rdata = 48'b110001101111111100000000000100001000000000000000;
			// PEs: 8 -> 17
			// srcs: (74, 69)(1908) -3 --> (1908) -3:PUNB, pass, PENB
			10'd68 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 16 -> 21
			// srcs: (75, 54)(1825) 1 --> (1825) 1:NI0, pass, PEGB5
			10'd69 : rdata = 48'b110001010000000000000000000000000000000011010000;
			// PEs: 23 -> 24
			// srcs: (76, 79)(1923) -6 --> (1923) -6:PENB, pass, PUNB
			10'd70 : rdata = 48'b110001101111111000000000000000000000001000000000;
			// PEs: 16 -> 22
			// srcs: (77, 57)(1828) 0 --> (1828) 0:NI2, pass, PEGB6
			10'd71 : rdata = 48'b110001010000001000000000000000000000000011100000;
			// PEs: 17 -> 24
			// srcs: (78, 89)(1996) 3 --> (1996) 3:PEGB1, pass, PUNB
			10'd72 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 16 -> 23
			// srcs: (79, 60)(1831) -3 --> (1831) -3:NI3, pass, PEGB7
			10'd73 : rdata = 48'b110001010000001100000000000000000000000011110000;
			// PEs: 16 -> 17
			// srcs: (80, 70)(1907) 0 --> (1907) 0:NI1, pass, PENB
			10'd74 : rdata = 48'b110001010000000100000000000000000000000100000000;
			// PEs: 8 -> 16
			// srcs: (81, 71)(1910) -2 --> (1910) -2:PUNB, pass, NI0
			10'd75 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 8 -> 17
			// srcs: (82, 72)(1911) 0 --> (1911) 0:PUNB, pass, PENB
			10'd76 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 18 -> 24
			// srcs: (83, 90)(1997) -6 --> (1997) -6:PEGB2, pass, PUNB
			10'd77 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 19 -> 24
			// srcs: (84, 91)(1999) 2 --> (1999) 2:PEGB3, pass, PUNB
			10'd78 : rdata = 48'b110001110000011000000000000000000000001000000000;
			// PEs: 20 -> 24
			// srcs: (85, 92)(2000) 6 --> (2000) 6:PEGB4, pass, PUNB
			10'd79 : rdata = 48'b110001110000100000000000000000000000001000000000;
			// PEs: 21 -> 24
			// srcs: (86, 93)(2002) -4 --> (2002) -4:PEGB5, pass, PUNB
			10'd80 : rdata = 48'b110001110000101000000000000000000000001000000000;
			// PEs: 22 -> 24
			// srcs: (87, 94)(2003) 2 --> (2003) 2:PEGB6, pass, PUNB
			10'd81 : rdata = 48'b110001110000110000000000000000000000001000000000;
			// PEs: 16 -> 17
			// srcs: (88, 73)(1910) -2 --> (1910) -2:NI0, pass, PENB
			10'd82 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 8 -> 16
			// srcs: (89, 74)(1913) 2 --> (1913) 2:PUNB, pass, NI0
			10'd83 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 8 -> 17
			// srcs: (90, 75)(1914) -4 --> (1914) -4:PUNB, pass, PENB
			10'd84 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 23 -> 24
			// srcs: (91, 95)(2005) 1 --> (2005) 1:PENB, pass, PUNB
			10'd85 : rdata = 48'b110001101111111000000000000000000000001000000000;
			// PEs: 17 -> 24
			// srcs: (92, 105)(2076) 0 --> (2076) 0:PEGB1, pass, PUNB
			10'd86 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 18 -> 24
			// srcs: (93, 106)(2077) 1 --> (2077) 1:PEGB2, pass, PUNB
			10'd87 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 19 -> 24
			// srcs: (94, 107)(2079) 0 --> (2079) 0:PEGB3, pass, PUNB
			10'd88 : rdata = 48'b110001110000011000000000000000000000001000000000;
			// PEs: 20 -> 24
			// srcs: (95, 108)(2080) 0 --> (2080) 0:PEGB4, pass, PUNB
			10'd89 : rdata = 48'b110001110000100000000000000000000000001000000000;
			// PEs: 16 -> 17
			// srcs: (96, 76)(1913) 2 --> (1913) 2:NI0, pass, PENB
			10'd90 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 8 -> 16
			// srcs: (97, 80)(1987) 4 --> (1987) 4:PUNB, pass, NI0
			10'd91 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 8 -> 17
			// srcs: (98, 81)(1988) -2 --> (1988) -2:PUNB, pass, PENB
			10'd92 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 21 -> 24
			// srcs: (99, 109)(2082) 2 --> (2082) 2:PEGB5, pass, PUNB
			10'd93 : rdata = 48'b110001110000101000000000000000000000001000000000;
			// PEs: 22 -> 24
			// srcs: (100, 110)(2083) 0 --> (2083) 0:PEGB6, pass, PUNB
			10'd94 : rdata = 48'b110001110000110000000000000000000000001000000000;
			// PEs: 23 -> 24
			// srcs: (101, 111)(2085) 0 --> (2085) 0:PENB, pass, PUNB
			10'd95 : rdata = 48'b110001101111111000000000000000000000001000000000;
			// PEs: 17 -> 24
			// srcs: (102, 121)(2158) 0 --> (2158) 0:PEGB1, pass, PUNB
			10'd96 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 18 -> 24
			// srcs: (103, 122)(2159) -3 --> (2159) -3:PEGB2, pass, PUNB
			10'd97 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 16 -> 17
			// srcs: (104, 82)(1987) 4 --> (1987) 4:NI0, pass, PENB
			10'd98 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 8 -> 16
			// srcs: (105, 83)(1990) -2 --> (1990) -2:PUNB, pass, NI0
			10'd99 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 8 -> 17
			// srcs: (106, 84)(1991) 1 --> (1991) 1:PUNB, pass, PENB
			10'd100 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 23 -> 24
			// srcs: (107, 123)(2165) 0 --> (2165) 0:PENB, pass, PUNB
			10'd101 : rdata = 48'b110001101111111000000000000000000000001000000000;
			// PEs: 23 -> 24
			// srcs: (108, 124)(2247) -2 --> (2247) -2:PENB, pass, PUNB
			10'd102 : rdata = 48'b110001101111111000000000000000000000001000000000;
			// PEs: 23 -> 24
			// srcs: (109, 125)(2327) 0 --> (2327) 0:PENB, pass, PUNB
			10'd103 : rdata = 48'b110001101111111000000000000000000000001000000000;
			// PEs: 18 -> 0
			// srcs: (110, 139)(2360) -10 --> (2360) -10:PEGB2, pass, PUGB0
			10'd104 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 20 -> 48
			// srcs: (111, 144)(2399) 0 --> (2399) 0:PEGB4, pass, PUGB6
			10'd105 : rdata = 48'b110001110000100000000000000000000000000000001110;
			// PEs: 16 -> 17
			// srcs: (112, 85)(1990) -2 --> (1990) -2:NI0, pass, PENB
			10'd106 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 8 -> 16
			// srcs: (113, 86)(1993) 0 --> (1993) 0:PUNB, pass, NI0
			10'd107 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 8 -> 17
			// srcs: (114, 87)(1994) 0 --> (1994) 0:PUNB, pass, PENB
			10'd108 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 23 -> 8
			// srcs: (115, 147)(2413) -6 --> (2413) -6:PENB, pass, PUGB1
			10'd109 : rdata = 48'b110001101111111000000000000000000000000000001001;
			// PEs: 19 -> 0
			// srcs: (116, 155)(1683) 1 --> (1683) 1:PEGB3, pass, PUGB0
			10'd110 : rdata = 48'b110001110000011000000000000000000000000000001000;
			// PEs: 17 -> 24
			// srcs: (117, 129)(1673) 0 --> (1673) 0:PEGB1, pass, PUNB
			10'd111 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 16 -> 17
			// srcs: (120, 88)(1993) 0 --> (1993) 0:NI0, pass, PENB
			10'd112 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 8 -> 16
			// srcs: (121, 96)(2067) -1 --> (2067) -1:PUNB, pass, NI0
			10'd113 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 8 -> 17
			// srcs: (122, 97)(2068) 0 --> (2068) 0:PUNB, pass, PENB
			10'd114 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 18 -> 32
			// srcs: (123, 154)(1680) 3 --> (1680) 3:PEGB2, pass, PUGB4
			10'd115 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 23 -> 48
			// srcs: (124, 159)(1695) 3 --> (1695) 3:PENB, pass, PUGB6
			10'd116 : rdata = 48'b110001101111111000000000000000000000000000001110;
			// PEs: 18 -> 24
			// srcs: (125, 130)(1674) 0 --> (1674) 0:PEGB2, pass, PUNB
			10'd117 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 16 -> 17
			// srcs: (128, 98)(2067) -1 --> (2067) -1:NI0, pass, PENB
			10'd118 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 8 -> 16
			// srcs: (129, 99)(2070) 4 --> (2070) 4:PUNB, pass, NI0
			10'd119 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 8 -> 17
			// srcs: (130, 100)(2071) 2 --> (2071) 2:PUNB, pass, PENB
			10'd120 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 17 -> 24
			// srcs: (133, 131)(1916) 2 --> (1916) 2:PEGB1, pass, PUNB
			10'd121 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 18 -> 32
			// srcs: (134, 166)(2528) -1 --> (2528) -1:PEGB2, pass, PUGB4
			10'd122 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 18 -> 48
			// srcs: (135, 180)(1860) 0 --> (1860) 0:PEGB2, pass, PUGB6
			10'd123 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 16 -> 17
			// srcs: (136, 101)(2070) 4 --> (2070) 4:NI0, pass, PENB
			10'd124 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 8 -> 16
			// srcs: (137, 102)(2073) 2 --> (2073) 2:PUNB, pass, NI0
			10'd125 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 8 -> 17
			// srcs: (138, 103)(2074) 4 --> (2074) 4:PUNB, pass, PENB
			10'd126 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 18 -> 24
			// srcs: (141, 132)(1917) 0 --> (1917) 0:PEGB2, pass, PUNB
			10'd127 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 23 -> 48
			// srcs: (143, 185)(1879) 4 --> (1879) 4:PENB, pass, PUGB6
			10'd128 : rdata = 48'b110001101111111000000000000000000000000000001110;
			// PEs: 16 -> 17
			// srcs: (144, 104)(2073) 2 --> (2073) 2:NI0, pass, PENB
			10'd129 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 8 -> 16
			// srcs: (145, 112)(2149) 4 --> (2149) 4:PUNB, pass, NI0
			10'd130 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 8 -> 17
			// srcs: (146, 113)(2150) 1 --> (2150) 1:PUNB, pass, PENB
			10'd131 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 19 -> 24
			// srcs: (149, 133)(1918) 1 --> (1918) 1:PEGB3, pass, PUNB
			10'd132 : rdata = 48'b110001110000011000000000000000000000001000000000;
			// PEs: 16 -> 17
			// srcs: (152, 114)(2149) 4 --> (2149) 4:NI0, pass, PENB
			10'd133 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 8 -> 16
			// srcs: (153, 115)(2152) 0 --> (2152) 0:PUNB, pass, NI0
			10'd134 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 8 -> 17
			// srcs: (154, 116)(2153) 4 --> (2153) 4:PUNB, pass, PENB
			10'd135 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 17 -> 48
			// srcs: (155, 191)(2691) -2 --> (2691) -2:PEGB1, pass, PUGB6
			10'd136 : rdata = 48'b110001110000001000000000000000000000000000001110;
			// PEs: 20 -> 24
			// srcs: (157, 134)(1919) 4 --> (1919) 4:PEGB4, pass, PUNB
			10'd137 : rdata = 48'b110001110000100000000000000000000000001000000000;
			// PEs: 16 -> 17
			// srcs: (160, 117)(2152) 0 --> (2152) 0:NI0, pass, PENB
			10'd138 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 8 -> 16
			// srcs: (161, 118)(2155) 2 --> (2155) 2:PUNB, pass, NI0
			10'd139 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 8 -> 17
			// srcs: (162, 119)(2156) 2 --> (2156) 2:PUNB, pass, PENB
			10'd140 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 17 -> 48
			// srcs: (163, 192)(2767) 2 --> (2767) 2:PEGB1, pass, PUGB6
			10'd141 : rdata = 48'b110001110000001000000000000000000000000000001110;
			// PEs: 19 -> 24
			// srcs: (165, 135)(2161) 0 --> (2161) 0:PEGB3, pass, PUNB
			10'd142 : rdata = 48'b110001110000011000000000000000000000001000000000;
			// PEs: 16 -> 17
			// srcs: (168, 120)(2155) 2 --> (2155) 2:NI0, pass, PENB
			10'd143 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 0 -> 16
			// srcs: (169, 140)(2365) -8 --> (2365) -8:PUGB0, pass, NI0
			10'd144 : rdata = 48'b110001110000000100000000000100000000000000000000;
			// PEs: 48 -> 17
			// srcs: (170, 141)(1585) -3 --> (1585) -3:PUGB6, pass, PENB
			10'd145 : rdata = 48'b110001110000110100000000000000000000000100000000;
			// PEs: 20 -> 24
			// srcs: (173, 136)(2162) 4 --> (2162) 4:PEGB4, pass, PUNB
			10'd146 : rdata = 48'b110001110000100000000000000000000000001000000000;
			// PEs: 21 -> 24
			// srcs: (174, 137)(2163) 3 --> (2163) 3:PEGB5, pass, PUNB
			10'd147 : rdata = 48'b110001110000101000000000000000000000001000000000;
			// PEs: 22 -> 24
			// srcs: (175, 138)(2164) 4 --> (2164) 4:PEGB6, pass, PUNB
			10'd148 : rdata = 48'b110001110000110000000000000000000000001000000000;
			// PEs: 16 -> 17
			// srcs: (176, 142)(2365) -8 --> (2365) -8:NI0, pass, PENB
			10'd149 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 56 -> 17
			// srcs: (177, 143)(1618) -6 --> (1618) -6:PUGB7, pass, PENB
			10'd150 : rdata = 48'b110001110000111100000000000000000000000100000000;
			// PEs: 56 -> 17
			// srcs: (178, 145)(1628) 2 --> (1628) 2:PUGB7, pass, PENB
			10'd151 : rdata = 48'b110001110000111100000000000000000000000100000000;
			// PEs: 22 -> 40
			// srcs: (179, 146)(2411) 0 --> (2411) 0:PEGB6, pass, PUGB5
			10'd152 : rdata = 48'b110001110000110000000000000000000000000000001101;
			// PEs: 24 -> 16
			// srcs: (180, 148)(2424) -5 --> (2424) -5:PUGB3, pass, NI0
			10'd153 : rdata = 48'b110001110000011100000000000100000000000000000000;
			// PEs: 0 -> 17
			// srcs: (181, 149)(1646) 0 --> (1646) 0:PUGB0, pass, PENB
			10'd154 : rdata = 48'b110001110000000100000000000000000000000100000000;
			// PEs: 21 -> 56
			// srcs: (182, 157)(1689) 0 --> (1689) 0:PEGB5, pass, PUGB7
			10'd155 : rdata = 48'b110001110000101000000000000000000000000000001111;
			// PEs: 22 -> 32
			// srcs: (183, 174)(2608) 0 --> (2608) 0:PEGB6, pass, PUGB4
			10'd156 : rdata = 48'b110001110000110000000000000000000000000000001100;
			// PEs: 17 -> 48
			// srcs: (184, 232)(2366) -11 --> (2366) -11:PEGB1, pass, PUGB6
			10'd157 : rdata = 48'b110001110000001000000000000000000000000000001110;
			// PEs: 16 -> 17
			// srcs: (187, 150)(2424) -5 --> (2424) -5:NI0, pass, PENB
			10'd158 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 22 -> 8
			// srcs: (190, 158)(1692) 0 --> (1692) 0:PEGB6, pass, PUGB1
			10'd159 : rdata = 48'b110001110000110000000000000000000000000000001001;
			// PEs: 17 -> 56
			// srcs: (191, 171)(2569) 7 --> (2569) 7:PEGB1, pass, PUGB7
			10'd160 : rdata = 48'b110001110000001000000000000000000000000000001111;
			// PEs: 17 -> 40
			// srcs: (192, 179)(1857) -2 --> (1857) -2:PEGB1, pass, PUGB5
			10'd161 : rdata = 48'b110001110000001000000000000000000000000000001101;
			// PEs: 17 -> 32
			// srcs: (193, 189)(2686) -3 --> (2686) -3:PEGB1, pass, PUGB4
			10'd162 : rdata = 48'b110001110000001000000000000000000000000000001100;
			// PEs: 19 -> 8
			// srcs: (198, 167)(2531) 2 --> (2531) 2:PEGB3, pass, PUGB1
			10'd163 : rdata = 48'b110001110000011000000000000000000000000000001001;
			// PEs: 20 -> 56
			// srcs: (199, 172)(2603) 0 --> (2603) 0:PEGB4, pass, PUGB7
			10'd164 : rdata = 48'b110001110000100000000000000000000000000000001111;
			// PEs: 21 -> 8
			// srcs: (200, 183)(1873) 2 --> (1873) 2:PEGB5, pass, PUGB1
			10'd165 : rdata = 48'b110001110000101000000000000000000000000000001001;
			// PEs: 17 -> 40
			// srcs: (201, 190)(2689) -2 --> (2689) -2:PEGB1, pass, PUGB5
			10'd166 : rdata = 48'b110001110000001000000000000000000000000000001101;
			// PEs: 17 -> 32
			// srcs: (202, 194)(2774) 0 --> (2774) 0:PEGB1, pass, PUGB4
			10'd167 : rdata = 48'b110001110000001000000000000000000000000000001100;
			// PEs: 20 -> 56
			// srcs: (207, 182)(1866) -3 --> (1866) -3:PEGB4, pass, PUGB7
			10'd168 : rdata = 48'b110001110000100000000000000000000000000000001111;
			// PEs: 20 -> 8
			// srcs: (210, 204)(2050) 0 --> (2050) 0:PEGB4, pass, PUGB1
			10'd169 : rdata = 48'b110001110000100000000000000000000000000000001001;
			// PEs: 17 -> 40
			// srcs: (211, 213)(2933) 4 --> (2933) 4:PEGB1, pass, PUGB5
			10'd170 : rdata = 48'b110001110000001000000000000000000000000000001101;
			// PEs: 22 -> 32
			// srcs: (212, 224)(3100) 2 --> (3100) 2:PEGB6, pass, PUGB4
			10'd171 : rdata = 48'b110001110000110000000000000000000000000000001100;
			// PEs: 18 -> 56
			// srcs: (215, 202)(2044) 0 --> (2044) 0:PEGB2, pass, PUGB7
			10'd172 : rdata = 48'b110001110000010000000000000000000000000000001111;
			// PEs: 17 -> 40
			// srcs: (220, 233)(2398) -10 --> (2398) -10:PEGB1, pass, PUGB5
			10'd173 : rdata = 48'b110001110000001000000000000000000000000000001101;
			// PEs: 17 -> 8
			// srcs: (221, 235)(2425) -5 --> (2425) -5:PEGB1, pass, PUGB1
			10'd174 : rdata = 48'b110001110000001000000000000000000000000000001001;
			// PEs: 19 -> 56
			// srcs: (223, 203)(2047) -4 --> (2047) -4:PEGB3, pass, PUGB7
			10'd175 : rdata = 48'b110001110000011000000000000000000000000000001111;
			// PEs: 8 -> 16
			// srcs: (229, 126)(1671) 2 --> (1671) 2:PUNB, pass, NI0
			10'd176 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 22 -> 56
			// srcs: (231, 206)(2056) 0 --> (2056) 0:PEGB6, pass, PUGB7
			10'd177 : rdata = 48'b110001110000110000000000000000000000000000001111;
			// PEs: 17 -> 56
			// srcs: (239, 212)(2930) 4 --> (2930) 4:PEGB1, pass, PUGB7
			10'd178 : rdata = 48'b110001110000001000000000000000000000000000001111;
			// PEs: 23 -> 56
			// srcs: (244, 225)(3102) 0 --> (3102) 0:PENB, pass, PUGB7
			10'd179 : rdata = 48'b110001101111111000000000000000000000000000001111;
			// PEs: 8 -> 23
			// srcs: (245, 127)(1672) 1 --> (1672) 1:PUNB, pass, PEGB7
			10'd180 : rdata = 48'b110001101111111100000000000000000000000011110000;
			// PEs: 8 -> 17
			// srcs: (246, 151)(1655) 6 --> (1655) 6:PUNB, pass, PENB
			10'd181 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 8 -> 17
			// srcs: (247, 153)(2457) -2 --> (2457) -2:PUNB, pass, PENB
			10'd182 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 48 -> 16
			// srcs: (248, 160)(2485) 8 --> (2485) 8:PUGB6, pass, NI1
			10'd183 : rdata = 48'b110001110000110100000000000100001000000000000000;
			// PEs: 24 -> 17
			// srcs: (249, 161)(1707) 9 --> (1707) 9:PUGB3, pass, PENB
			10'd184 : rdata = 48'b110001110000011100000000000000000000000100000000;
			// PEs: 17 -> 32
			// srcs: (253, 236)(2435) 2 --> (2435) 2:PEGB1, pass, PUGB4
			10'd185 : rdata = 48'b110001110000001000000000000000000000000000001100;
			// PEs: 16 -> 23
			// srcs: (254, 128)(1671) 2 --> (1671) 2:NI0, pass, PEGB7
			10'd186 : rdata = 48'b110001010000000000000000000000000000000011110000;
			// PEs: 16 -> 17
			// srcs: (255, 162)(2485) 8 --> (2485) 8:NI1, pass, PENB
			10'd187 : rdata = 48'b110001010000000100000000000000000000000100000000;
			// PEs: 0 -> 16
			// srcs: (256, 163)(2510) -2 --> (2510) -2:PUGB0, pass, NI0
			10'd188 : rdata = 48'b110001110000000100000000000100000000000000000000;
			// PEs: 32 -> 17
			// srcs: (257, 164)(1732) 0 --> (1732) 0:PUGB4, pass, PENB
			10'd189 : rdata = 48'b110001110000100100000000000000000000000100000000;
			// PEs: 23 -> 24
			// srcs: (261, 152)(2454) 3 --> (2454) 3:PENB, pass, PUNB
			10'd190 : rdata = 48'b110001101111111000000000000000000000001000000000;
			// PEs: 17 -> 8
			// srcs: (262, 238)(2486) 17 --> (2486) 17:PEGB1, pass, PUGB1
			10'd191 : rdata = 48'b110001110000001000000000000000000000000000001001;
			// PEs: 16 -> 17
			// srcs: (263, 165)(2510) -2 --> (2510) -2:NI0, pass, PENB
			10'd192 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 24 -> 16
			// srcs: (264, 168)(2537) -4 --> (2537) -4:PUGB3, pass, NI0
			10'd193 : rdata = 48'b110001110000011100000000000100000000000000000000;
			// PEs: 40 -> 17
			// srcs: (265, 169)(1759) 2 --> (1759) 2:PUGB5, pass, PENB
			10'd194 : rdata = 48'b110001110000101100000000000000000000000100000000;
			// PEs: 20 -> 24
			// srcs: (269, 156)(1686) -1 --> (1686) -1:PEGB4, pass, PUNB
			10'd195 : rdata = 48'b110001110000100000000000000000000000001000000000;
			// PEs: 17 -> 56
			// srcs: (270, 239)(2511) -2 --> (2511) -2:PEGB1, pass, PUGB7
			10'd196 : rdata = 48'b110001110000001000000000000000000000000000001111;
			// PEs: 16 -> 17
			// srcs: (271, 170)(2537) -4 --> (2537) -4:NI0, pass, PENB
			10'd197 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 23 -> 24
			// srcs: (274, 175)(2612) 6 --> (2612) 6:PENB, pass, PUNB
			10'd198 : rdata = 48'b110001101111111000000000000000000000001000000000;
			// PEs: 19 -> 24
			// srcs: (282, 181)(1863) 6 --> (1863) 6:PEGB3, pass, PUNB
			10'd199 : rdata = 48'b110001110000011000000000000000000000001000000000;
			// PEs: 0 -> 17
			// srcs: (290, 173)(1827) 3 --> (1827) 3:PUGB0, pass, PENB
			10'd200 : rdata = 48'b110001110000000100000000000000000000000100000000;
			// PEs: 24 -> 16
			// srcs: (291, 176)(2617) 4 --> (2617) 4:PUGB3, pass, NI0
			10'd201 : rdata = 48'b110001110000011100000000000100000000000000000000;
			// PEs: 8 -> 17
			// srcs: (292, 177)(1839) -6 --> (1839) -6:PUNB, pass, PENB
			10'd202 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 17 -> 24
			// srcs: (293, 193)(2772) -1 --> (2772) -1:PEGB1, pass, PUNB
			10'd203 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 17 -> 32
			// srcs: (297, 244)(2607) 2 --> (2607) 2:PEGB1, pass, PUGB4
			10'd204 : rdata = 48'b110001110000001000000000000000000000000000001100;
			// PEs: 16 -> 17
			// srcs: (298, 178)(2617) 4 --> (2617) 4:NI0, pass, PENB
			10'd205 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 56 -> 17
			// srcs: (299, 184)(2655) -2 --> (2655) -2:PUGB7, pass, PENB
			10'd206 : rdata = 48'b110001110000111100000000000000000000000100000000;
			// PEs: 8 -> 16
			// srcs: (300, 186)(2678) 4 --> (2678) 4:PUNB, pass, NI0
			10'd207 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 24 -> 17
			// srcs: (301, 187)(1900) 0 --> (1900) 0:PUGB3, pass, PENB
			10'd208 : rdata = 48'b110001110000011100000000000000000000000100000000;
			// PEs: 17 -> 24
			// srcs: (302, 201)(2041) 2 --> (2041) 2:PEGB1, pass, PUNB
			10'd209 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 21 -> 24
			// srcs: (303, 205)(2053) 4 --> (2053) 4:PEGB5, pass, PUNB
			10'd210 : rdata = 48'b110001110000101000000000000000000000001000000000;
			// PEs: 21 -> 0
			// srcs: (304, 223)(3096) 2 --> (3096) 2:PEGB5, pass, PUGB0
			10'd211 : rdata = 48'b110001110000101000000000000000000000000000001000;
			// PEs: 17 -> 48
			// srcs: (305, 245)(2618) -2 --> (2618) -2:PEGB1, pass, PUGB6
			10'd212 : rdata = 48'b110001110000001000000000000000000000000000001110;
			// PEs: 17 -> 32
			// srcs: (306, 249)(2656) -4 --> (2656) -4:PEGB1, pass, PUGB4
			10'd213 : rdata = 48'b110001110000001000000000000000000000000000001100;
			// PEs: 16 -> 17
			// srcs: (307, 188)(2678) 4 --> (2678) 4:NI0, pass, PENB
			10'd214 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 40 -> 16
			// srcs: (308, 195)(2802) 2 --> (2802) 2:PUGB5, pass, NI0
			10'd215 : rdata = 48'b110001110000101100000000000100000000000000000000;
			// PEs: 8 -> 17
			// srcs: (309, 196)(2023) 1 --> (2023) 1:PUNB, pass, PENB
			10'd216 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 17 -> 24
			// srcs: (311, 208)(2848) -1 --> (2848) -1:PEGB1, pass, PUNB
			10'd217 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 17 -> 48
			// srcs: (314, 250)(2679) 4 --> (2679) 4:PEGB1, pass, PUGB6
			10'd218 : rdata = 48'b110001110000001000000000000000000000000000001110;
			// PEs: 16 -> 17
			// srcs: (315, 197)(2802) 2 --> (2802) 2:NI0, pass, PENB
			10'd219 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 48 -> 16
			// srcs: (316, 198)(2810) -3 --> (2810) -3:PUGB6, pass, NI0
			10'd220 : rdata = 48'b110001110000110100000000000100000000000000000000;
			// PEs: 8 -> 17
			// srcs: (317, 199)(2032) 0 --> (2032) 0:PUNB, pass, PENB
			10'd221 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 17 -> 24
			// srcs: (319, 209)(2851) 6 --> (2851) 6:PEGB1, pass, PUNB
			10'd222 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 17 -> 48
			// srcs: (322, 257)(2803) 3 --> (2803) 3:PEGB1, pass, PUGB6
			10'd223 : rdata = 48'b110001110000001000000000000000000000000000001110;
			// PEs: 16 -> 17
			// srcs: (323, 200)(2810) -3 --> (2810) -3:NI0, pass, PENB
			10'd224 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 17 -> 24
			// srcs: (327, 210)(2853) 6 --> (2853) 6:PEGB1, pass, PUNB
			10'd225 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 17 -> 40
			// srcs: (330, 258)(2811) -3 --> (2811) -3:PEGB1, pass, PUGB5
			10'd226 : rdata = 48'b110001110000001000000000000000000000000000001101;
			// PEs: 17 -> 24
			// srcs: (335, 211)(2928) 5 --> (2928) 5:PEGB1, pass, PUNB
			10'd227 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 20 -> 24
			// srcs: (343, 222)(3022) -2 --> (3022) -2:PEGB4, pass, PUNB
			10'd228 : rdata = 48'b110001110000100000000000000000000000001000000000;
			// PEs: 17 -> 24
			// srcs: (351, 234)(2409) 8 --> (2409) 8:PEGB1, pass, PUNB
			10'd229 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 17 -> 24
			// srcs: (359, 237)(2458) -2 --> (2458) -2:PEGB1, pass, PUNB
			10'd230 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 17 -> 24
			// srcs: (367, 243)(2538) -2 --> (2538) -2:PEGB1, pass, PUNB
			10'd231 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 8 -> 17
			// srcs: (385, 207)(2836) 0 --> (2836) 0:PUNB, pass, PENB
			10'd232 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 48 -> 16
			// srcs: (386, 214)(2972) -9 --> (2972) -9:PUGB6, pass, NI0
			10'd233 : rdata = 48'b110001110000110100000000000100000000000000000000;
			// PEs: 0 -> 17
			// srcs: (387, 215)(2194) -1 --> (2194) -1:PUGB0, pass, PENB
			10'd234 : rdata = 48'b110001110000000100000000000000000000000100000000;
			// PEs: 17 -> 24
			// srcs: (392, 259)(2837) 0 --> (2837) 0:PEGB1, pass, PUNB
			10'd235 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 16 -> 17
			// srcs: (393, 216)(2972) -9 --> (2972) -9:NI0, pass, PENB
			10'd236 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 0 -> 17
			// srcs: (394, 217)(3003) 0 --> (3003) 0:PUGB0, pass, PENB
			10'd237 : rdata = 48'b110001110000000100000000000000000000000100000000;
			// PEs: 8 -> 17
			// srcs: (395, 218)(3005) 1 --> (3005) 1:PUNB, pass, PENB
			10'd238 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 17 -> 32
			// srcs: (400, 263)(2973) -10 --> (2973) -10:PEGB1, pass, PUGB4
			10'd239 : rdata = 48'b110001110000001000000000000000000000000000001100;
			// PEs: 22 -> 24
			// srcs: (403, 267)(3021) -1 --> (3021) -1:PEGB6, pass, PUNB
			10'd240 : rdata = 48'b110001110000110000000000000000000000001000000000;
			// PEs: 8 -> 17
			// srcs: (549, 219)(3008) -12 --> (3008) -12:PUNB, pass, PENB
			10'd241 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 8 -> 17
			// srcs: (564, 220)(3010) -4 --> (3010) -4:PUNB, pass, PENB
			10'd242 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 8 -> 17
			// srcs: (580, 221)(3015) -3 --> (3015) -3:PUNB, pass, PENB
			10'd243 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 24 -> 16
			// srcs: (581, 226)(3105) -1 --> (3105) -1:PUGB3, pass, NI0
			10'd244 : rdata = 48'b110001110000011100000000000100000000000000000000;
			// PEs: 48 -> 17
			// srcs: (582, 227)(2329) -4 --> (2329) -4:PUGB6, pass, PENB
			10'd245 : rdata = 48'b110001110000110100000000000000000000000100000000;
			// PEs: 16 -> 17
			// srcs: (593, 228)(3105) -1 --> (3105) -1:NI0, pass, PENB
			10'd246 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 48 -> 16
			// srcs: (594, 229)(2359) 9 --> (2359) 9:PUGB6, pass, NI0
			10'd247 : rdata = 48'b110001110000110100000000000100000000000000000000;
			// PEs: 0 -> 17
			// srcs: (595, 230)(2361) -16 --> (2361) -16:PUGB0, pass, PENB
			10'd248 : rdata = 48'b110001110000000100000000000000000000000100000000;
			// PEs: 17 -> 56
			// srcs: (600, 268)(3106) -5 --> (3106) -5:PEGB1, pass, PUGB7
			10'd249 : rdata = 48'b110001110000001000000000000000000000000000001111;
			// PEs: 16 -> 17
			// srcs: (601, 231)(2359) 9 --> (2359) 9:NI0, pass, PENB
			10'd250 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 8 -> 16
			// srcs: (602, 240)(2532) -2 --> (2532) -2:PUNB, pass, NI0
			10'd251 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 48 -> 17
			// srcs: (603, 241)(2534) -6 --> (2534) -6:PUGB6, pass, PENB
			10'd252 : rdata = 48'b110001110000110100000000000000000000000100000000;
			// PEs: 17 -> 40
			// srcs: (608, 269)(2362) -7 --> (2362) -7:PEGB1, pass, PUGB5
			10'd253 : rdata = 48'b110001110000001000000000000000000000000000001101;
			// PEs: 16 -> 17
			// srcs: (609, 242)(2532) -2 --> (2532) -2:NI0, pass, PENB
			10'd254 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 48 -> 16
			// srcs: (610, 246)(2651) 5 --> (2651) 5:PUGB6, pass, NI0
			10'd255 : rdata = 48'b110001110000110100000000000100000000000000000000;
			// PEs: 8 -> 17
			// srcs: (611, 247)(2653) 5 --> (2653) 5:PUNB, pass, PENB
			10'd256 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 17 -> 24
			// srcs: (616, 276)(2535) -8 --> (2535) -8:PEGB1, pass, PUNB
			10'd257 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 16 -> 17
			// srcs: (617, 248)(2651) 5 --> (2651) 5:NI0, pass, PENB
			10'd258 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 0 -> 16
			// srcs: (618, 251)(2766) -4 --> (2766) -4:PUGB0, pass, NI0
			10'd259 : rdata = 48'b110001110000000100000000000100000000000000000000;
			// PEs: 48 -> 17
			// srcs: (619, 252)(2768) 6 --> (2768) 6:PUGB6, pass, PENB
			10'd260 : rdata = 48'b110001110000110100000000000000000000000100000000;
			// PEs: 17 -> 40
			// srcs: (624, 277)(2654) 10 --> (2654) 10:PEGB1, pass, PUGB5
			10'd261 : rdata = 48'b110001110000001000000000000000000000000000001101;
			// PEs: 16 -> 17
			// srcs: (625, 253)(2766) -4 --> (2766) -4:NI0, pass, PENB
			10'd262 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 40 -> 16
			// srcs: (626, 254)(2798) 5 --> (2798) 5:PUGB5, pass, NI0
			10'd263 : rdata = 48'b110001110000101100000000000100000000000000000000;
			// PEs: 0 -> 17
			// srcs: (627, 255)(2800) -1 --> (2800) -1:PUGB0, pass, PENB
			10'd264 : rdata = 48'b110001110000000100000000000000000000000100000000;
			// PEs: 16 -> 17
			// srcs: (633, 256)(2798) 5 --> (2798) 5:NI0, pass, PENB
			10'd265 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 56 -> 16
			// srcs: (634, 260)(2906) 0 --> (2906) 0:PUGB7, pass, NI0
			10'd266 : rdata = 48'b110001110000111100000000000100000000000000000000;
			// PEs: 8 -> 17
			// srcs: (635, 261)(2908) -2 --> (2908) -2:PUNB, pass, PENB
			10'd267 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 8 -> 21
			// srcs: (636, 281)(2764) -4 --> (2764) -4:PUNB, pass, PEGB5
			10'd268 : rdata = 48'b110001101111111100000000000000000000000011010000;
			// PEs: 17 -> 24
			// srcs: (640, 282)(2801) 4 --> (2801) 4:PEGB1, pass, PUNB
			10'd269 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 16 -> 17
			// srcs: (641, 262)(2906) 0 --> (2906) 0:NI0, pass, PENB
			10'd270 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 21 -> 24
			// srcs: (642, 288)(3019) -11 --> (3019) -11:PEGB5, pass, PUNB
			10'd271 : rdata = 48'b110001110000101000000000000000000000001000000000;
			// PEs: 24 -> 16
			// srcs: (650, 264)(2984) -3 --> (2984) -3:PUGB3, pass, NI0
			10'd272 : rdata = 48'b110001110000011100000000000100000000000000000000;
			// PEs: 0 -> 17
			// srcs: (651, 265)(2986) -2 --> (2986) -2:PUGB0, pass, PENB
			10'd273 : rdata = 48'b110001110000000100000000000000000000000100000000;
			// PEs: 16 -> 17
			// srcs: (657, 266)(2984) -3 --> (2984) -3:NI0, pass, PENB
			10'd274 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 0 -> 16
			// srcs: (658, 270)(2396) -2 --> (2396) -2:PUGB0, pass, NI0
			10'd275 : rdata = 48'b110001110000000100000000000100000000000000000000;
			// PEs: 17 -> 0
			// srcs: (664, 287)(2987) -5 --> (2987) -5:PEGB1, pass, PUGB0
			10'd276 : rdata = 48'b110001110000001000000000000000000000000000001000;
			// PEs: 40 -> 17
			// srcs: (726, 271)(2401) -8 --> (2401) -8:PUGB5, pass, PENB
			10'd277 : rdata = 48'b110001110000101100000000000000000000000100000000;
			// PEs: 16 -> 17
			// srcs: (733, 272)(2396) -2 --> (2396) -2:NI0, pass, PENB
			10'd278 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 32 -> 16
			// srcs: (734, 273)(2507) 15 --> (2507) 15:PUGB4, pass, NI0
			10'd279 : rdata = 48'b110001110000100100000000000100000000000000000000;
			// PEs: 56 -> 17
			// srcs: (735, 274)(2512) 1 --> (2512) 1:PUGB7, pass, PENB
			10'd280 : rdata = 48'b110001110000111100000000000000000000000100000000;
			// PEs: 17 -> 32
			// srcs: (740, 292)(2402) -10 --> (2402) -10:PEGB1, pass, PUGB4
			10'd281 : rdata = 48'b110001110000001000000000000000000000000000001100;
			// PEs: 16 -> 17
			// srcs: (741, 275)(2507) 15 --> (2507) 15:NI0, pass, PENB
			10'd282 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 17 -> 24
			// srcs: (748, 293)(2513) 16 --> (2513) 16:PEGB1, pass, PUNB
			10'd283 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 0 -> 16
			// srcs: (978, 278)(2688) -3 --> (2688) -3:PUGB0, pass, NI0
			10'd284 : rdata = 48'b110001110000000100000000000100000000000000000000;
			// PEs: 48 -> 17
			// srcs: (979, 279)(2693) -1 --> (2693) -1:PUGB6, pass, PENB
			10'd285 : rdata = 48'b110001110000110100000000000000000000000100000000;
			// PEs: 16 -> 17
			// srcs: (985, 280)(2688) -3 --> (2688) -3:NI0, pass, PENB
			10'd286 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 48 -> 17
			// srcs: (986, 283)(2914) -9 --> (2914) -9:PUGB6, pass, PENB
			10'd287 : rdata = 48'b110001110000110100000000000000000000000100000000;
			// PEs: 8 -> 16
			// srcs: (987, 284)(2959) 11 --> (2959) 11:PUNB, pass, NI0
			10'd288 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 24 -> 17
			// srcs: (988, 285)(2964) -8 --> (2964) -8:PUGB3, pass, PENB
			10'd289 : rdata = 48'b110001110000011100000000000000000000000100000000;
			// PEs: 17 -> 48
			// srcs: (992, 297)(2694) -4 --> (2694) -4:PEGB1, pass, PUGB6
			10'd290 : rdata = 48'b110001110000001000000000000000000000000000001110;
			// PEs: 16 -> 17
			// srcs: (994, 286)(2959) 11 --> (2959) 11:NI0, pass, PENB
			10'd291 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 40 -> 16
			// srcs: (995, 289)(2368) -29 --> (2368) -29:PUGB5, pass, NI0
			10'd292 : rdata = 48'b110001110000101100000000000100000000000000000000;
			// PEs: 0 -> 17
			// srcs: (1017, 290)(2379) 11 --> (2379) 11:PUGB0, pass, PENB
			10'd293 : rdata = 48'b110001110000000100000000000000000000000100000000;
			// PEs: 16 -> 17
			// srcs: (1024, 291)(2368) -29 --> (2368) -29:NI0, pass, PENB
			10'd294 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 17 -> 24
			// srcs: (1031, 302)(2380) -18 --> (2380) -18:PEGB1, pass, PUNB
			10'd295 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 32 -> 16
			// srcs: (1127, 294)(2611) 18 --> (2611) 18:PUGB4, pass, NI0
			10'd296 : rdata = 48'b110001110000100100000000000100000000000000000000;
			// PEs: 56 -> 17
			// srcs: (1158, 295)(2622) 9 --> (2622) 9:PUGB7, pass, PENB
			10'd297 : rdata = 48'b110001110000111100000000000000000000000100000000;
			// PEs: 16 -> 17
			// srcs: (1165, 296)(2611) 18 --> (2611) 18:NI0, pass, PENB
			10'd298 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 8 -> 17
			// srcs: (1166, 298)(2759) -18 --> (2759) -18:PUNB, pass, PENB
			10'd299 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 8 -> 17
			// srcs: (1167, 299)(2904) 27 --> (2904) 27:PUNB, pass, PENB
			10'd300 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 8 -> 17
			// srcs: (1168, 300)(2954) 6 --> (2954) 6:PUNB, pass, PENB
			10'd301 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 8 -> 17
			// srcs: (1169, 301)(3002) -9 --> (3002) -9:PUNB, pass, PENB
			10'd302 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 24 -> 17
			// srcs: (1170, 307)(3037) -9 --> (3037) -9:PUGB3, pass, PENB
			10'd303 : rdata = 48'b110001110000011100000000000000000000000100000000;
			// PEs: 17 -> 40
			// srcs: (1172, 303)(2623) 27 --> (2623) 27:PEGB1, pass, PUGB5
			10'd304 : rdata = 48'b110001110000001000000000000000000000000000001101;
			// PEs: 17 -> 8
			// srcs: (1173, 304)(2771) -20 --> (2771) -20:PEGB1, pass, PUGB1
			10'd305 : rdata = 48'b110001110000001000000000000000000000000000001001;
			// PEs: 17 -> 32
			// srcs: (1174, 305)(2916) 16 --> (2916) 16:PEGB1, pass, PUGB4
			10'd306 : rdata = 48'b110001110000001000000000000000000000000000001100;
			// PEs: 17 -> 56
			// srcs: (1175, 306)(2966) 9 --> (2966) 9:PEGB1, pass, PUGB7
			10'd307 : rdata = 48'b110001110000001000000000000000000000000000001111;
			// PEs: 17 -> 32
			// srcs: (1186, 311)(3038) -37 --> (3038) -37:PEGB1, pass, PUGB4
			10'd308 : rdata = 48'b110001110000001000000000000000000000000000001100;
			// PEs: 8 -> 16
			// srcs: (1423, 308)(2795) -21 --> (2795) -21:PUNB, pass, NI0
			10'd309 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 24 -> 17
			// srcs: (1429, 309)(2843) -10 --> (2843) -10:PUGB3, pass, PENB
			10'd310 : rdata = 48'b110001110000011100000000000000000000000100000000;
			// PEs: 16 -> 17
			// srcs: (1436, 310)(2795) -21 --> (2795) -21:NI0, pass, PENB
			10'd311 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 17 -> 24
			// srcs: (1443, 312)(2844) -31 --> (2844) -31:PEGB1, pass, PUNB
			10'd312 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 8 -> 17
			// srcs: (1525, 313)(3140) 47 --> (3140) 47:PUNB, pass, PENB
			10'd313 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 8 -> 18
			// srcs: (1526, 314)(3140) 47 --> (3140) 47:PUNB, pass, PEGB2
			10'd314 : rdata = 48'b110001101111111100000000000000000000000010100000;
			// PEs: 8 -> 19
			// srcs: (1528, 315)(3140) 47 --> (3140) 47:PUNB, pass, PEGB3
			10'd315 : rdata = 48'b110001101111111100000000000000000000000010110000;
			// PEs: 8 -> 20
			// srcs: (1529, 316)(3140) 47 --> (3140) 47:PUNB, pass, PEGB4
			10'd316 : rdata = 48'b110001101111111100000000000000000000000011000000;
			// PEs: 8 -> 21
			// srcs: (1531, 317)(3140) 47 --> (3140) 47:PUNB, pass, PEGB5
			10'd317 : rdata = 48'b110001101111111100000000000000000000000011010000;
			// PEs: 8 -> 22
			// srcs: (1532, 318)(3140) 47 --> (3140) 47:PUNB, pass, PEGB6
			10'd318 : rdata = 48'b110001101111111100000000000000000000000011100000;
			// PEs: 8 -> 23
			// srcs: (1534, 319)(3140) 47 --> (3140) 47:PUNB, pass, PEGB7
			10'd319 : rdata = 48'b110001101111111100000000000000000000000011110000;
			// PEs: 8 -> 17
			// srcs: (1606, 320)(3140) 47 --> (3140) 47:PUNB, pass, PENB
			10'd320 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 8 -> 18
			// srcs: (1607, 321)(3140) 47 --> (3140) 47:PUNB, pass, PEGB2
			10'd321 : rdata = 48'b110001101111111100000000000000000000000010100000;
			// PEs: 8 -> 19
			// srcs: (1608, 322)(3140) 47 --> (3140) 47:PUNB, pass, PEGB3
			10'd322 : rdata = 48'b110001101111111100000000000000000000000010110000;
			// PEs: 8 -> 20
			// srcs: (1609, 323)(3140) 47 --> (3140) 47:PUNB, pass, PEGB4
			10'd323 : rdata = 48'b110001101111111100000000000000000000000011000000;
			// PEs: 8 -> 17
			// srcs: (1610, 324)(3140) 47 --> (3140) 47:PUNB, pass, PENB
			10'd324 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 8 -> 21
			// srcs: (1611, 325)(3140) 47 --> (3140) 47:PUNB, pass, PEGB5
			10'd325 : rdata = 48'b110001101111111100000000000000000000000011010000;
			// PEs: 8 -> 22
			// srcs: (1612, 326)(3140) 47 --> (3140) 47:PUNB, pass, PEGB6
			10'd326 : rdata = 48'b110001101111111100000000000000000000000011100000;
			// PEs: 8 -> 18
			// srcs: (1613, 327)(3140) 47 --> (3140) 47:PUNB, pass, PEGB2
			10'd327 : rdata = 48'b110001101111111100000000000000000000000010100000;
			// PEs: 8 -> 23
			// srcs: (1614, 328)(3140) 47 --> (3140) 47:PUNB, pass, PEGB7
			10'd328 : rdata = 48'b110001101111111100000000000000000000000011110000;
			// PEs: 8 -> 19
			// srcs: (1616, 329)(3140) 47 --> (3140) 47:PUNB, pass, PEGB3
			10'd329 : rdata = 48'b110001101111111100000000000000000000000010110000;
			// PEs: 8 -> 20
			// srcs: (1619, 330)(3140) 47 --> (3140) 47:PUNB, pass, PEGB4
			10'd330 : rdata = 48'b110001101111111100000000000000000000000011000000;
			// PEs: 8 -> 21
			// srcs: (1622, 331)(3140) 47 --> (3140) 47:PUNB, pass, PEGB5
			10'd331 : rdata = 48'b110001101111111100000000000000000000000011010000;
			// PEs: 8 -> 22
			// srcs: (1625, 332)(3140) 47 --> (3140) 47:PUNB, pass, PEGB6
			10'd332 : rdata = 48'b110001101111111100000000000000000000000011100000;
			// PEs: 8 -> 23
			// srcs: (1628, 333)(3140) 47 --> (3140) 47:PUNB, pass, PEGB7
			10'd333 : rdata = 48'b110001101111111100000000000000000000000011110000;
			// PEs: 8 -> 17
			// srcs: (1687, 334)(3140) 47 --> (3140) 47:PUNB, pass, PENB
			10'd334 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 8 -> 18
			// srcs: (1688, 335)(3140) 47 --> (3140) 47:PUNB, pass, PEGB2
			10'd335 : rdata = 48'b110001101111111100000000000000000000000010100000;
			// PEs: 8 -> 19
			// srcs: (1690, 336)(3140) 47 --> (3140) 47:PUNB, pass, PEGB3
			10'd336 : rdata = 48'b110001101111111100000000000000000000000010110000;
			// PEs: 8 -> 20
			// srcs: (1691, 337)(3140) 47 --> (3140) 47:PUNB, pass, PEGB4
			10'd337 : rdata = 48'b110001101111111100000000000000000000000011000000;
			// PEs: 8 -> 21
			// srcs: (1693, 338)(3140) 47 --> (3140) 47:PUNB, pass, PEGB5
			10'd338 : rdata = 48'b110001101111111100000000000000000000000011010000;
			// PEs: 8 -> 22
			// srcs: (1694, 339)(3140) 47 --> (3140) 47:PUNB, pass, PEGB6
			10'd339 : rdata = 48'b110001101111111100000000000000000000000011100000;
			// PEs: 8 -> 23
			// srcs: (1696, 340)(3140) 47 --> (3140) 47:PUNB, pass, PEGB7
			10'd340 : rdata = 48'b110001101111111100000000000000000000000011110000;
			// PEs: 8 -> 17
			// srcs: (1767, 341)(3140) 47 --> (3140) 47:PUNB, pass, PENB
			10'd341 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 8 -> 18
			// srcs: (1768, 342)(3140) 47 --> (3140) 47:PUNB, pass, PEGB2
			10'd342 : rdata = 48'b110001101111111100000000000000000000000010100000;
			// PEs: 8 -> 19
			// srcs: (1770, 343)(3140) 47 --> (3140) 47:PUNB, pass, PEGB3
			10'd343 : rdata = 48'b110001101111111100000000000000000000000010110000;
			// PEs: 8 -> 20
			// srcs: (1771, 344)(3140) 47 --> (3140) 47:PUNB, pass, PEGB4
			10'd344 : rdata = 48'b110001101111111100000000000000000000000011000000;
			// PEs: 8 -> 21
			// srcs: (1773, 345)(3140) 47 --> (3140) 47:PUNB, pass, PEGB5
			10'd345 : rdata = 48'b110001101111111100000000000000000000000011010000;
			// PEs: 8 -> 22
			// srcs: (1774, 346)(3140) 47 --> (3140) 47:PUNB, pass, PEGB6
			10'd346 : rdata = 48'b110001101111111100000000000000000000000011100000;
			// PEs: 8 -> 23
			// srcs: (1776, 347)(3140) 47 --> (3140) 47:PUNB, pass, PEGB7
			10'd347 : rdata = 48'b110001101111111100000000000000000000000011110000;
			// PEs: 8 -> 17
			// srcs: (1790, 348)(3140) 47 --> (3140) 47:PUNB, pass, PENB
			10'd348 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 8 -> 18
			// srcs: (1793, 349)(3140) 47 --> (3140) 47:PUNB, pass, PEGB2
			10'd349 : rdata = 48'b110001101111111100000000000000000000000010100000;
			// PEs: 8 -> 19
			// srcs: (1796, 350)(3140) 47 --> (3140) 47:PUNB, pass, PEGB3
			10'd350 : rdata = 48'b110001101111111100000000000000000000000010110000;
			// PEs: 8 -> 20
			// srcs: (1799, 351)(3140) 47 --> (3140) 47:PUNB, pass, PEGB4
			10'd351 : rdata = 48'b110001101111111100000000000000000000000011000000;
			// PEs: 8 -> 21
			// srcs: (1806, 352)(3140) 47 --> (3140) 47:PUNB, pass, PEGB5
			10'd352 : rdata = 48'b110001101111111100000000000000000000000011010000;
			// PEs: 8 -> 22
			// srcs: (1809, 353)(3140) 47 --> (3140) 47:PUNB, pass, PEGB6
			10'd353 : rdata = 48'b110001101111111100000000000000000000000011100000;
			// PEs: 8 -> 23
			// srcs: (1812, 354)(3140) 47 --> (3140) 47:PUNB, pass, PEGB7
			10'd354 : rdata = 48'b110001101111111100000000000000000000000011110000;
			// PEs: 8 -> 17
			// srcs: (1849, 355)(3140) 47 --> (3140) 47:PUNB, pass, PENB
			10'd355 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 8 -> 18
			// srcs: (1850, 356)(3140) 47 --> (3140) 47:PUNB, pass, PEGB2
			10'd356 : rdata = 48'b110001101111111100000000000000000000000010100000;
			// PEs: 8 -> 19
			// srcs: (1851, 357)(3140) 47 --> (3140) 47:PUNB, pass, PEGB3
			10'd357 : rdata = 48'b110001101111111100000000000000000000000010110000;
			// PEs: 8 -> 20
			// srcs: (1852, 358)(3140) 47 --> (3140) 47:PUNB, pass, PEGB4
			10'd358 : rdata = 48'b110001101111111100000000000000000000000011000000;
			// PEs: 8 -> 21
			// srcs: (1853, 359)(3140) 47 --> (3140) 47:PUNB, pass, PEGB5
			10'd359 : rdata = 48'b110001101111111100000000000000000000000011010000;
			// PEs: 8 -> 22
			// srcs: (1854, 360)(3140) 47 --> (3140) 47:PUNB, pass, PEGB6
			10'd360 : rdata = 48'b110001101111111100000000000000000000000011100000;
			// PEs: 8 -> 23
			// srcs: (1856, 361)(3140) 47 --> (3140) 47:PUNB, pass, PEGB7
			10'd361 : rdata = 48'b110001101111111100000000000000000000000011110000;
			// PEs: 8 -> 17
			// srcs: (1929, 362)(3140) 47 --> (3140) 47:PUNB, pass, PENB
			10'd362 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 8 -> 18
			// srcs: (1930, 363)(3140) 47 --> (3140) 47:PUNB, pass, PEGB2
			10'd363 : rdata = 48'b110001101111111100000000000000000000000010100000;
			// PEs: 8 -> 19
			// srcs: (1932, 364)(3140) 47 --> (3140) 47:PUNB, pass, PEGB3
			10'd364 : rdata = 48'b110001101111111100000000000000000000000010110000;
			// PEs: 8 -> 20
			// srcs: (1933, 365)(3140) 47 --> (3140) 47:PUNB, pass, PEGB4
			10'd365 : rdata = 48'b110001101111111100000000000000000000000011000000;
			// PEs: 8 -> 21
			// srcs: (1935, 366)(3140) 47 --> (3140) 47:PUNB, pass, PEGB5
			10'd366 : rdata = 48'b110001101111111100000000000000000000000011010000;
			// PEs: 8 -> 22
			// srcs: (1936, 367)(3140) 47 --> (3140) 47:PUNB, pass, PEGB6
			10'd367 : rdata = 48'b110001101111111100000000000000000000000011100000;
			// PEs: 8 -> 23
			// srcs: (1938, 368)(3140) 47 --> (3140) 47:PUNB, pass, PEGB7
			10'd368 : rdata = 48'b110001101111111100000000000000000000000011110000;
			// PEs: 8 -> 17
			// srcs: (1974, 369)(3140) 47 --> (3140) 47:PUNB, pass, PENB
			10'd369 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 8 -> 18
			// srcs: (1977, 370)(3140) 47 --> (3140) 47:PUNB, pass, PEGB2
			10'd370 : rdata = 48'b110001101111111100000000000000000000000010100000;
			// PEs: 8 -> 19
			// srcs: (1980, 371)(3140) 47 --> (3140) 47:PUNB, pass, PEGB3
			10'd371 : rdata = 48'b110001101111111100000000000000000000000010110000;
			// PEs: 8 -> 20
			// srcs: (1983, 372)(3140) 47 --> (3140) 47:PUNB, pass, PEGB4
			10'd372 : rdata = 48'b110001101111111100000000000000000000000011000000;
			// PEs: 8 -> 21
			// srcs: (1986, 373)(3140) 47 --> (3140) 47:PUNB, pass, PEGB5
			10'd373 : rdata = 48'b110001101111111100000000000000000000000011010000;
			// PEs: 8 -> 22
			// srcs: (1989, 374)(3140) 47 --> (3140) 47:PUNB, pass, PEGB6
			10'd374 : rdata = 48'b110001101111111100000000000000000000000011100000;
			// PEs: 8 -> 23
			// srcs: (1992, 375)(3140) 47 --> (3140) 47:PUNB, pass, PEGB7
			10'd375 : rdata = 48'b110001101111111100000000000000000000000011110000;
			// PEs: 8 -> 17
			// srcs: (2009, 376)(3140) 47 --> (3140) 47:PUNB, pass, PENB
			10'd376 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 8 -> 18
			// srcs: (2010, 377)(3140) 47 --> (3140) 47:PUNB, pass, PEGB2
			10'd377 : rdata = 48'b110001101111111100000000000000000000000010100000;
			// PEs: 8 -> 19
			// srcs: (2012, 378)(3140) 47 --> (3140) 47:PUNB, pass, PEGB3
			10'd378 : rdata = 48'b110001101111111100000000000000000000000010110000;
			// PEs: 8 -> 20
			// srcs: (2013, 379)(3140) 47 --> (3140) 47:PUNB, pass, PEGB4
			10'd379 : rdata = 48'b110001101111111100000000000000000000000011000000;
			// PEs: 8 -> 21
			// srcs: (2015, 380)(3140) 47 --> (3140) 47:PUNB, pass, PEGB5
			10'd380 : rdata = 48'b110001101111111100000000000000000000000011010000;
			// PEs: 8 -> 22
			// srcs: (2016, 381)(3140) 47 --> (3140) 47:PUNB, pass, PEGB6
			10'd381 : rdata = 48'b110001101111111100000000000000000000000011100000;
			// PEs: 8 -> 23
			// srcs: (2018, 382)(3140) 47 --> (3140) 47:PUNB, pass, PEGB7
			10'd382 : rdata = 48'b110001101111111100000000000000000000000011110000;
			// PEs: 8 -> 17
			// srcs: (2091, 383)(3140) 47 --> (3140) 47:PUNB, pass, PENB
			10'd383 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 8 -> 18
			// srcs: (2092, 384)(3140) 47 --> (3140) 47:PUNB, pass, PEGB2
			10'd384 : rdata = 48'b110001101111111100000000000000000000000010100000;
			// PEs: 8 -> 19
			// srcs: (2094, 385)(3140) 47 --> (3140) 47:PUNB, pass, PEGB3
			10'd385 : rdata = 48'b110001101111111100000000000000000000000010110000;
			// PEs: 8 -> 20
			// srcs: (2095, 386)(3140) 47 --> (3140) 47:PUNB, pass, PEGB4
			10'd386 : rdata = 48'b110001101111111100000000000000000000000011000000;
			// PEs: 8 -> 21
			// srcs: (2096, 387)(3140) 47 --> (3140) 47:PUNB, pass, PEGB5
			10'd387 : rdata = 48'b110001101111111100000000000000000000000011010000;
			// PEs: 8 -> 22
			// srcs: (2097, 388)(3140) 47 --> (3140) 47:PUNB, pass, PEGB6
			10'd388 : rdata = 48'b110001101111111100000000000000000000000011100000;
			// PEs: 8 -> 23
			// srcs: (2098, 389)(3140) 47 --> (3140) 47:PUNB, pass, PEGB7
			10'd389 : rdata = 48'b110001101111111100000000000000000000000011110000;
			// PEs: 8 -> 17
			// srcs: (2158, 390)(3140) 47 --> (3140) 47:PUNB, pass, PENB
			10'd390 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 8 -> 18
			// srcs: (2161, 391)(3140) 47 --> (3140) 47:PUNB, pass, PEGB2
			10'd391 : rdata = 48'b110001101111111100000000000000000000000010100000;
			// PEs: 8 -> 19
			// srcs: (2164, 392)(3140) 47 --> (3140) 47:PUNB, pass, PEGB3
			10'd392 : rdata = 48'b110001101111111100000000000000000000000010110000;
			// PEs: 8 -> 20
			// srcs: (2167, 393)(3140) 47 --> (3140) 47:PUNB, pass, PEGB4
			10'd393 : rdata = 48'b110001101111111100000000000000000000000011000000;
			// PEs: 8 -> 21
			// srcs: (2170, 394)(3140) 47 --> (3140) 47:PUNB, pass, PEGB5
			10'd394 : rdata = 48'b110001101111111100000000000000000000000011010000;
			// PEs: 8 -> 17
			// srcs: (2171, 395)(3140) 47 --> (3140) 47:PUNB, pass, PENB
			10'd395 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 8 -> 18
			// srcs: (2172, 396)(3140) 47 --> (3140) 47:PUNB, pass, PEGB2
			10'd396 : rdata = 48'b110001101111111100000000000000000000000010100000;
			// PEs: 8 -> 22
			// srcs: (2173, 397)(3140) 47 --> (3140) 47:PUNB, pass, PEGB6
			10'd397 : rdata = 48'b110001101111111100000000000000000000000011100000;
			// PEs: 8 -> 19
			// srcs: (2174, 398)(3140) 47 --> (3140) 47:PUNB, pass, PEGB3
			10'd398 : rdata = 48'b110001101111111100000000000000000000000010110000;
			// PEs: 8 -> 20
			// srcs: (2175, 399)(3140) 47 --> (3140) 47:PUNB, pass, PEGB4
			10'd399 : rdata = 48'b110001101111111100000000000000000000000011000000;
			// PEs: 8 -> 23
			// srcs: (2176, 400)(3140) 47 --> (3140) 47:PUNB, pass, PEGB7
			10'd400 : rdata = 48'b110001101111111100000000000000000000000011110000;
			// PEs: 8 -> 21
			// srcs: (2177, 401)(3140) 47 --> (3140) 47:PUNB, pass, PEGB5
			10'd401 : rdata = 48'b110001101111111100000000000000000000000011010000;
			// PEs: 8 -> 22
			// srcs: (2178, 402)(3140) 47 --> (3140) 47:PUNB, pass, PEGB6
			10'd402 : rdata = 48'b110001101111111100000000000000000000000011100000;
			// PEs: 8 -> 23
			// srcs: (2180, 403)(3140) 47 --> (3140) 47:PUNB, pass, PEGB7
			10'd403 : rdata = 48'b110001101111111100000000000000000000000011110000;
			// PEs: 8 -> 17
			// srcs: (2251, 404)(3140) 47 --> (3140) 47:PUNB, pass, PENB
			10'd404 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 8 -> 18
			// srcs: (2252, 405)(3140) 47 --> (3140) 47:PUNB, pass, PEGB2
			10'd405 : rdata = 48'b110001101111111100000000000000000000000010100000;
			// PEs: 8 -> 19
			// srcs: (2254, 406)(3140) 47 --> (3140) 47:PUNB, pass, PEGB3
			10'd406 : rdata = 48'b110001101111111100000000000000000000000010110000;
			// PEs: 8 -> 20
			// srcs: (2255, 407)(3140) 47 --> (3140) 47:PUNB, pass, PEGB4
			10'd407 : rdata = 48'b110001101111111100000000000000000000000011000000;
			// PEs: 8 -> 21
			// srcs: (2257, 408)(3140) 47 --> (3140) 47:PUNB, pass, PEGB5
			10'd408 : rdata = 48'b110001101111111100000000000000000000000011010000;
			// PEs: 8 -> 22
			// srcs: (2258, 409)(3140) 47 --> (3140) 47:PUNB, pass, PEGB6
			10'd409 : rdata = 48'b110001101111111100000000000000000000000011100000;
			// PEs: 8 -> 23
			// srcs: (2260, 410)(3140) 47 --> (3140) 47:PUNB, pass, PEGB7
			10'd410 : rdata = 48'b110001101111111100000000000000000000000011110000;
			default : rdata = 48'b000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 17) begin
	always @(*) begin
		case(address)
			// PEs: 17, 17 -> 16
			// srcs: (1, 0)(23) -3, (808) -3 --> (1592) 9:ND0, NW0, *, PEGB0
			10'd0 : rdata = 48'b000110110000000001000000000000000000000010000000;
			// PEs: 17, 17 -> 17
			// srcs: (2, 1)(104) 0, (889) -1 --> (1673) 0:ND1, NW1, *, NI0
			10'd1 : rdata = 48'b000110110000000101000000001100000000000000000000;
			// PEs: 17, 17 -> 16
			// srcs: (3, 2)(185) 0, (970) 2 --> (1754) 0:ND2, NW2, *, PEGB0
			10'd2 : rdata = 48'b000110110000001001000000010000000000000010000000;
			// PEs: 17, 17 -> 16
			// srcs: (4, 3)(265) 0, (1050) -3 --> (1834) 0:ND3, NW3, *, PEGB0
			10'd3 : rdata = 48'b000110110000001101000000011000000000000010000000;
			// PEs: 17, 17 -> 17
			// srcs: (5, 4)(347) 1, (1132) 2 --> (1916) 2:ND4, NW4, *, NI1
			10'd4 : rdata = 48'b000110110000010001000000100100001000000000000000;
			// PEs: 17, 17 -> 16
			// srcs: (6, 5)(427) -3, (1212) -1 --> (1996) 3:ND5, NW5, *, PEGB0
			10'd5 : rdata = 48'b000110110000010101000000101000000000000010000000;
			// PEs: 17, 17 -> 16
			// srcs: (7, 6)(507) -3, (1292) 0 --> (2076) 0:ND6, NW6, *, PEGB0
			10'd6 : rdata = 48'b000110110000011001000000110000000000000010000000;
			// PEs: 17, 17 -> 16
			// srcs: (8, 7)(589) 1, (1374) 0 --> (2158) 0:ND7, NW7, *, PEGB0
			10'd7 : rdata = 48'b000110110000011101000000111000000000000010000000;
			// PEs: 17, 17 -> 19
			// srcs: (9, 8)(669) 1, (1454) -1 --> (2238) -1:ND8, NW8, *, PEGB3
			10'd8 : rdata = 48'b000110110000100001000001000000000000000010110000;
			// PEs: 17, 17 -> 21
			// srcs: (10, 9)(749) 1, (1534) 2 --> (2318) 2:ND9, NW9, *, PEGB5
			10'd9 : rdata = 48'b000110110000100101000001001000000000000011010000;
			// PEs: 17, 17 -> 17
			// srcs: (11, 10)(108) 2, (893) 0 --> (1677) 0:ND10, NW10, *, NI2
			10'd10 : rdata = 48'b000110110000101001000001010100010000000000000000;
			// PEs: 17, 17 -> 17
			// srcs: (12, 11)(288) 1, (1073) -2 --> (1857) -2:ND11, NW11, *, NI3
			10'd11 : rdata = 48'b000110110000101101000001011100011000000000000000;
			// PEs: 17, 17 -> 17
			// srcs: (13, 12)(472) -1, (1257) -2 --> (2041) 2:ND12, NW12, *, NI4
			10'd12 : rdata = 48'b000110110000110001000001100100100000000000000000;
			// PEs: 17, 17 -> 17
			// srcs: (14, 13)(656) -1, (1441) 2 --> (2225) -2:ND13, NW13, *, NI5
			10'd13 : rdata = 48'b000110110000110101000001101100101000000000000000;
			// PEs: 16 -> 
			// srcs: (32, 14)(1654) -4 --> (1654) -4:PENB, pass, 
			10'd14 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 16, 17 -> 17
			// srcs: (38, 15)(1653) 0, (1654) -4 --> (2434) -4:PENB, ALU, +, NI6
			10'd15 : rdata = 48'b000011101111111000111111111100110000000000000000;
			// PEs: 16 -> 
			// srcs: (49, 16)(1789) 4 --> (1789) 4:PENB, pass, 
			10'd16 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 16, 17 -> 17
			// srcs: (55, 17)(1788) 3, (1789) 4 --> (2569) 7:PENB, ALU, +, NI7
			10'd17 : rdata = 48'b000011101111111000111111111100111000000000000000;
			// PEs: 16 -> 
			// srcs: (76, 18)(1908) -3 --> (1908) -3:PENB, pass, 
			10'd18 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 16, 17 -> 17
			// srcs: (82, 19)(1907) 0, (1908) -3 --> (2686) -3:PENB, ALU, +, NI8
			10'd19 : rdata = 48'b000011101111111000111111111101000000000000000000;
			// PEs: 16 -> 
			// srcs: (84, 20)(1911) 0 --> (1911) 0:PENB, pass, 
			10'd20 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 16, 17 -> 17
			// srcs: (90, 21)(1910) -2, (1911) 0 --> (2689) -2:PENB, ALU, +, NI9
			10'd21 : rdata = 48'b000011101111111000111111111101001000000000000000;
			// PEs: 16 -> 
			// srcs: (92, 22)(1914) -4 --> (1914) -4:PENB, pass, 
			10'd22 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 16, 17 -> 17
			// srcs: (98, 23)(1913) 2, (1914) -4 --> (2691) -2:PENB, ALU, +, NI10
			10'd23 : rdata = 48'b000011101111111000111111111101010000000000000000;
			// PEs: 16 -> 
			// srcs: (100, 24)(1988) -2 --> (1988) -2:PENB, pass, 
			10'd24 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 16, 17 -> 17
			// srcs: (106, 25)(1987) 4, (1988) -2 --> (2767) 2:PENB, ALU, +, NI11
			10'd25 : rdata = 48'b000011101111111000111111111101011000000000000000;
			// PEs: 16 -> 17
			// srcs: (108, 26)(1991) 1 --> (1991) 1:PENB, pass, NI12
			10'd26 : rdata = 48'b110001101111111000000000000101100000000000000000;
			// PEs: 17 -> 16
			// srcs: (112, 42)(1673) 0 --> (1673) 0:NI0, pass, PEGB0
			10'd27 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 16, 17 -> 17
			// srcs: (114, 27)(1990) -2, (1991) 1 --> (2772) -1:PENB, NI12, +, NI0
			10'd28 : rdata = 48'b000011101111111010100001100100000000000000000000;
			// PEs: 16 -> 
			// srcs: (116, 28)(1994) 0 --> (1994) 0:PENB, pass, 
			10'd29 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 16, 17 -> 17
			// srcs: (122, 29)(1993) 0, (1994) 0 --> (2774) 0:PENB, ALU, +, NI12
			10'd30 : rdata = 48'b000011101111111000111111111101100000000000000000;
			// PEs: 16 -> 17
			// srcs: (124, 30)(2068) 0 --> (2068) 0:PENB, pass, NI13
			10'd31 : rdata = 48'b110001101111111000000000000101101000000000000000;
			// PEs: 17 -> 16
			// srcs: (128, 43)(1916) 2 --> (1916) 2:NI1, pass, PEGB0
			10'd32 : rdata = 48'b110001010000000100000000000000000000000010000000;
			// PEs: 16, 17 -> 17
			// srcs: (130, 31)(2067) -1, (2068) 0 --> (2848) -1:PENB, NI13, +, NI1
			10'd33 : rdata = 48'b000011101111111010100001101100001000000000000000;
			// PEs: 16 -> 
			// srcs: (132, 32)(2071) 2 --> (2071) 2:PENB, pass, 
			10'd34 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 16, 17 -> 17
			// srcs: (138, 33)(2070) 4, (2071) 2 --> (2851) 6:PENB, ALU, +, NI13
			10'd35 : rdata = 48'b000011101111111000111111111101101000000000000000;
			// PEs: 16 -> 
			// srcs: (140, 34)(2074) 4 --> (2074) 4:PENB, pass, 
			10'd36 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 16, 17 -> 17
			// srcs: (146, 35)(2073) 2, (2074) 4 --> (2853) 6:PENB, ALU, +, NI14
			10'd37 : rdata = 48'b000011101111111000111111111101110000000000000000;
			// PEs: 16 -> 17
			// srcs: (148, 36)(2150) 1 --> (2150) 1:PENB, pass, NI15
			10'd38 : rdata = 48'b110001101111111000000000000101111000000000000000;
			// PEs: 17 -> 16
			// srcs: (149, 68)(2691) -2 --> (2691) -2:NI10, pass, PEGB0
			10'd39 : rdata = 48'b110001010000101000000000000000000000000010000000;
			// PEs: 16, 17 -> 17
			// srcs: (154, 37)(2149) 4, (2150) 1 --> (2928) 5:PENB, NI15, +, NI10
			10'd40 : rdata = 48'b000011101111111010100001111101010000000000000000;
			// PEs: 16 -> 17
			// srcs: (156, 38)(2153) 4 --> (2153) 4:PENB, pass, NI15
			10'd41 : rdata = 48'b110001101111111000000000000101111000000000000000;
			// PEs: 17 -> 16
			// srcs: (158, 69)(2767) 2 --> (2767) 2:NI11, pass, PEGB0
			10'd42 : rdata = 48'b110001010000101100000000000000000000000010000000;
			// PEs: 16, 17 -> 17
			// srcs: (162, 39)(2152) 0, (2153) 4 --> (2930) 4:PENB, NI15, +, NI11
			10'd43 : rdata = 48'b000011101111111010100001111101011000000000000000;
			// PEs: 16 -> 
			// srcs: (164, 40)(2156) 2 --> (2156) 2:PENB, pass, 
			10'd44 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 16, 17 -> 17
			// srcs: (170, 41)(2155) 2, (2156) 2 --> (2933) 4:PENB, ALU, +, NI15
			10'd45 : rdata = 48'b000011101111111000111111111101111000000000000000;
			// PEs: 16 -> 
			// srcs: (172, 44)(1585) -3 --> (1585) -3:PENB, pass, 
			10'd46 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 16, 17 -> 16
			// srcs: (178, 45)(2365) -8, (1585) -3 --> (2366) -11:PENB, ALU, +, PEGB0
			10'd47 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 19, 16 -> 17
			// srcs: (179, 46)(2397) -4, (1618) -6 --> (2398) -10:PEGB3, PENB, +, NI16
			10'd48 : rdata = 48'b000011110000011011011111110110000000000000000000;
			// PEs: 21, 16 -> 17
			// srcs: (180, 47)(2408) 6, (1628) 2 --> (2409) 8:PEGB5, PENB, +, NI17
			10'd49 : rdata = 48'b000011110000101011011111110110001000000000000000;
			// PEs: 16 -> 17
			// srcs: (183, 48)(1646) 0 --> (1646) 0:PENB, pass, NI18
			10'd50 : rdata = 48'b110001101111111000000000000110010000000000000000;
			// PEs: 17 -> 16
			// srcs: (185, 58)(2569) 7 --> (2569) 7:NI7, pass, PEGB0
			10'd51 : rdata = 48'b110001010000011100000000000000000000000010000000;
			// PEs: 17 -> 16
			// srcs: (186, 62)(1857) -2 --> (1857) -2:NI3, pass, PEGB0
			10'd52 : rdata = 48'b110001010000001100000000000000000000000010000000;
			// PEs: 17 -> 16
			// srcs: (187, 66)(2686) -3 --> (2686) -3:NI8, pass, PEGB0
			10'd53 : rdata = 48'b110001010000100000000000000000000000000010000000;
			// PEs: 16, 17 -> 17
			// srcs: (189, 49)(2424) -5, (1646) 0 --> (2425) -5:PENB, NI18, +, NI3
			10'd54 : rdata = 48'b000011101111111010100010010100011000000000000000;
			// PEs: 17 -> 16
			// srcs: (196, 67)(2689) -2 --> (2689) -2:NI9, pass, PEGB0
			10'd55 : rdata = 48'b110001010000100100000000000000000000000010000000;
			// PEs: 17 -> 16
			// srcs: (197, 71)(2774) 0 --> (2774) 0:NI12, pass, PEGB0
			10'd56 : rdata = 48'b110001010000110000000000000000000000000010000000;
			// PEs: 17 -> 16
			// srcs: (205, 83)(2933) 4 --> (2933) 4:NI15, pass, PEGB0
			10'd57 : rdata = 48'b110001010000111100000000000000000000000010000000;
			// PEs: 17 -> 16
			// srcs: (215, 95)(2398) -10 --> (2398) -10:NI16, pass, PEGB0
			10'd58 : rdata = 48'b110001010001000000000000000000000000000010000000;
			// PEs: 17 -> 16
			// srcs: (216, 97)(2425) -5 --> (2425) -5:NI3, pass, PEGB0
			10'd59 : rdata = 48'b110001010000001100000000000000000000000010000000;
			// PEs: 17 -> 16
			// srcs: (234, 82)(2930) 4 --> (2930) 4:NI11, pass, PEGB0
			10'd60 : rdata = 48'b110001010000101100000000000000000000000010000000;
			// PEs: 17, 16 -> 16
			// srcs: (248, 50)(2434) -4, (1655) 6 --> (2435) 2:NI6, PENB, +, PEGB0
			10'd61 : rdata = 48'b000011010000011011011111110000000000000010000000;
			// PEs: 16, 17 -> 17
			// srcs: (249, 51)(2457) -2, (1677) 0 --> (2458) -2:PENB, NI2, +, NI3
			10'd62 : rdata = 48'b000011101111111010100000010100011000000000000000;
			// PEs: 16 -> 
			// srcs: (251, 52)(1707) 9 --> (1707) 9:PENB, pass, 
			10'd63 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 16, 17 -> 16
			// srcs: (257, 53)(2485) 8, (1707) 9 --> (2486) 17:PENB, ALU, +, PEGB0
			10'd64 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 16 -> 
			// srcs: (259, 54)(1732) 0 --> (1732) 0:PENB, pass, 
			10'd65 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 16, 17 -> 16
			// srcs: (265, 55)(2510) -2, (1732) 0 --> (2511) -2:PENB, ALU, +, PEGB0
			10'd66 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 16 -> 
			// srcs: (267, 56)(1759) 2 --> (1759) 2:PENB, pass, 
			10'd67 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 16, 17 -> 17
			// srcs: (273, 57)(2537) -4, (1759) 2 --> (2538) -2:PENB, ALU, +, NI2
			10'd68 : rdata = 48'b000011101111111000111111111100010000000000000000;
			// PEs: 17 -> 16
			// srcs: (285, 70)(2772) -1 --> (2772) -1:NI0, pass, PEGB0
			10'd69 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 21, 16 -> 16
			// srcs: (292, 59)(2606) -1, (1827) 3 --> (2607) 2:PEGB5, PENB, +, PEGB0
			10'd70 : rdata = 48'b000011110000101011011111110000000000000010000000;
			// PEs: 16 -> 17
			// srcs: (294, 60)(1839) -6 --> (1839) -6:PENB, pass, NI0
			10'd71 : rdata = 48'b110001101111111000000000000100000000000000000000;
			// PEs: 17 -> 16
			// srcs: (296, 76)(2041) 2 --> (2041) 2:NI4, pass, PEGB0
			10'd72 : rdata = 48'b110001010000010000000000000000000000000010000000;
			// PEs: 16, 17 -> 16
			// srcs: (300, 61)(2617) 4, (1839) -6 --> (2618) -2:PENB, NI0, +, PEGB0
			10'd73 : rdata = 48'b000011101111111010100000000000000000000010000000;
			// PEs: 16, 22 -> 16
			// srcs: (301, 63)(2655) -2, (1876) -2 --> (2656) -4:PENB, PEGB6, +, PEGB0
			10'd74 : rdata = 48'b000011101111111011100001100000000000000010000000;
			// PEs: 16 -> 17
			// srcs: (303, 64)(1900) 0 --> (1900) 0:PENB, pass, NI0
			10'd75 : rdata = 48'b110001101111111000000000000100000000000000000000;
			// PEs: 17 -> 16
			// srcs: (306, 78)(2848) -1 --> (2848) -1:NI1, pass, PEGB0
			10'd76 : rdata = 48'b110001010000000100000000000000000000000010000000;
			// PEs: 16, 17 -> 16
			// srcs: (309, 65)(2678) 4, (1900) 0 --> (2679) 4:PENB, NI0, +, PEGB0
			10'd77 : rdata = 48'b000011101111111010100000000000000000000010000000;
			// PEs: 16 -> 17
			// srcs: (311, 72)(2023) 1 --> (2023) 1:PENB, pass, NI0
			10'd78 : rdata = 48'b110001101111111000000000000100000000000000000000;
			// PEs: 17 -> 16
			// srcs: (314, 79)(2851) 6 --> (2851) 6:NI13, pass, PEGB0
			10'd79 : rdata = 48'b110001010000110100000000000000000000000010000000;
			// PEs: 16, 17 -> 16
			// srcs: (317, 73)(2802) 2, (2023) 1 --> (2803) 3:PENB, NI0, +, PEGB0
			10'd80 : rdata = 48'b000011101111111010100000000000000000000010000000;
			// PEs: 16 -> 17
			// srcs: (319, 74)(2032) 0 --> (2032) 0:PENB, pass, NI0
			10'd81 : rdata = 48'b110001101111111000000000000100000000000000000000;
			// PEs: 17 -> 16
			// srcs: (322, 80)(2853) 6 --> (2853) 6:NI14, pass, PEGB0
			10'd82 : rdata = 48'b110001010000111000000000000000000000000010000000;
			// PEs: 16, 17 -> 16
			// srcs: (325, 75)(2810) -3, (2032) 0 --> (2811) -3:PENB, NI0, +, PEGB0
			10'd83 : rdata = 48'b000011101111111010100000000000000000000010000000;
			// PEs: 17 -> 16
			// srcs: (330, 81)(2928) 5 --> (2928) 5:NI10, pass, PEGB0
			10'd84 : rdata = 48'b110001010000101000000000000000000000000010000000;
			// PEs: 17 -> 16
			// srcs: (346, 96)(2409) 8 --> (2409) 8:NI17, pass, PEGB0
			10'd85 : rdata = 48'b110001010001000100000000000000000000000010000000;
			// PEs: 17 -> 16
			// srcs: (354, 98)(2458) -2 --> (2458) -2:NI3, pass, PEGB0
			10'd86 : rdata = 48'b110001010000001100000000000000000000000010000000;
			// PEs: 17 -> 16
			// srcs: (362, 101)(2538) -2 --> (2538) -2:NI2, pass, PEGB0
			10'd87 : rdata = 48'b110001010000001000000000000000000000000010000000;
			// PEs: 16, 23 -> 16
			// srcs: (387, 77)(2836) 0, (2059) 0 --> (2837) 0:PENB, PEGB7, +, PEGB0
			10'd88 : rdata = 48'b000011101111111011100001110000000000000010000000;
			// PEs: 16 -> 
			// srcs: (389, 84)(2194) -1 --> (2194) -1:PENB, pass, 
			10'd89 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 16, 17 -> 16
			// srcs: (395, 85)(2972) -9, (2194) -1 --> (2973) -10:PENB, ALU, +, PEGB0
			10'd90 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 16, 17 -> 17
			// srcs: (396, 86)(3003) 0, (2225) -2 --> (3004) -2:PENB, NI5, +, NI0
			10'd91 : rdata = 48'b000011101111111010100000101100000000000000000000;
			// PEs: 16, 18 -> 18
			// srcs: (397, 87)(3005) 1, (2228) 0 --> (3006) 1:PENB, PEGB2, +, PENB
			10'd92 : rdata = 48'b000011101111111011100000100000000000000100000000;
			// PEs: 17 -> 18
			// srcs: (404, 112)(3004) -2 --> (3004) -2:NI0, pass, PENB
			10'd93 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 16, 19 -> 17
			// srcs: (558, 88)(3008) -12, (2231) -2 --> (3009) -14:PENB, PEGB3, +, NI0
			10'd94 : rdata = 48'b000011101111111011100000110100000000000000000000;
			// PEs: 16, 20 -> 18
			// srcs: (566, 89)(3010) -4, (2234) 0 --> (3011) -4:PENB, PEGB4, +, PENB
			10'd95 : rdata = 48'b000011101111111011100001000000000000000100000000;
			// PEs: 17 -> 18
			// srcs: (573, 113)(3009) -14 --> (3009) -14:NI0, pass, PENB
			10'd96 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 16, 21 -> 21
			// srcs: (589, 90)(3015) -3, (2237) -3 --> (3016) -6:PENB, PEGB5, +, PEGB5
			10'd97 : rdata = 48'b000011101111111011100001010000000000000011010000;
			// PEs: 16 -> 
			// srcs: (590, 91)(2329) -4 --> (2329) -4:PENB, pass, 
			10'd98 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 16, 17 -> 16
			// srcs: (595, 92)(3105) -1, (2329) -4 --> (3106) -5:PENB, ALU, +, PEGB0
			10'd99 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 16 -> 
			// srcs: (597, 93)(2361) -16 --> (2361) -16:PENB, pass, 
			10'd100 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 16, 17 -> 16
			// srcs: (603, 94)(2359) 9, (2361) -16 --> (2362) -7:PENB, ALU, +, PEGB0
			10'd101 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 16 -> 
			// srcs: (605, 99)(2534) -6 --> (2534) -6:PENB, pass, 
			10'd102 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 16, 17 -> 16
			// srcs: (611, 100)(2532) -2, (2534) -6 --> (2535) -8:PENB, ALU, +, PEGB0
			10'd103 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 16 -> 
			// srcs: (613, 102)(2653) 5 --> (2653) 5:PENB, pass, 
			10'd104 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 16, 17 -> 16
			// srcs: (619, 103)(2651) 5, (2653) 5 --> (2654) 10:PENB, ALU, +, PEGB0
			10'd105 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 16 -> 
			// srcs: (621, 104)(2768) 6 --> (2768) 6:PENB, pass, 
			10'd106 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 16, 17 -> 21
			// srcs: (627, 105)(2766) -4, (2768) 6 --> (2769) 2:PENB, ALU, +, PEGB5
			10'd107 : rdata = 48'b000011101111111000111111111000000000000011010000;
			// PEs: 16 -> 
			// srcs: (629, 106)(2800) -1 --> (2800) -1:PENB, pass, 
			10'd108 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 16, 17 -> 16
			// srcs: (635, 107)(2798) 5, (2800) -1 --> (2801) 4:PENB, ALU, +, PEGB0
			10'd109 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 16 -> 
			// srcs: (637, 108)(2908) -2 --> (2908) -2:PENB, pass, 
			10'd110 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 16, 17 -> 17
			// srcs: (643, 109)(2906) 0, (2908) -2 --> (2909) -2:PENB, ALU, +, NI0
			10'd111 : rdata = 48'b000011101111111000111111111100000000000000000000;
			// PEs: 16 -> 
			// srcs: (653, 110)(2986) -2 --> (2986) -2:PENB, pass, 
			10'd112 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 16, 17 -> 16
			// srcs: (659, 111)(2984) -3, (2986) -2 --> (2987) -5:PENB, ALU, +, PEGB0
			10'd113 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 16 -> 
			// srcs: (728, 114)(2401) -8 --> (2401) -8:PENB, pass, 
			10'd114 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 16, 17 -> 16
			// srcs: (735, 115)(2396) -2, (2401) -8 --> (2402) -10:PENB, ALU, +, PEGB0
			10'd115 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 16 -> 
			// srcs: (737, 116)(2512) 1 --> (2512) 1:PENB, pass, 
			10'd116 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 16, 17 -> 16
			// srcs: (743, 117)(2507) 15, (2512) 1 --> (2513) 16:PENB, ALU, +, PEGB0
			10'd117 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 16 -> 
			// srcs: (981, 118)(2693) -1 --> (2693) -1:PENB, pass, 
			10'd118 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 16, 17 -> 16
			// srcs: (987, 119)(2688) -3, (2693) -1 --> (2694) -4:PENB, ALU, +, PEGB0
			10'd119 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 17, 16 -> 17
			// srcs: (988, 120)(2909) -2, (2914) -9 --> (2915) -11:NI0, PENB, +, NI1
			10'd120 : rdata = 48'b000011010000000011011111110100001000000000000000;
			// PEs: 16 -> 
			// srcs: (990, 121)(2964) -8 --> (2964) -8:PENB, pass, 
			10'd121 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 16, 17 -> 17
			// srcs: (996, 122)(2959) 11, (2964) -8 --> (2965) 3:PENB, ALU, +, NI0
			10'd122 : rdata = 48'b000011101111111000111111111100000000000000000000;
			// PEs: 16 -> 
			// srcs: (1019, 123)(2379) 11 --> (2379) 11:PENB, pass, 
			10'd123 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 16, 17 -> 16
			// srcs: (1026, 124)(2368) -29, (2379) 11 --> (2380) -18:PENB, ALU, +, PEGB0
			10'd124 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 16 -> 
			// srcs: (1160, 125)(2622) 9 --> (2622) 9:PENB, pass, 
			10'd125 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 16, 17 -> 16
			// srcs: (1167, 126)(2611) 18, (2622) 9 --> (2623) 27:PENB, ALU, +, PEGB0
			10'd126 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 16, 21 -> 16
			// srcs: (1168, 127)(2759) -18, (2770) -2 --> (2771) -20:PENB, PEGB5, +, PEGB0
			10'd127 : rdata = 48'b000011101111111011100001010000000000000010000000;
			// PEs: 16, 17 -> 16
			// srcs: (1169, 128)(2904) 27, (2915) -11 --> (2916) 16:PENB, NI1, +, PEGB0
			10'd128 : rdata = 48'b000011101111111010100000001000000000000010000000;
			// PEs: 16, 17 -> 16
			// srcs: (1170, 129)(2954) 6, (2965) 3 --> (2966) 9:PENB, NI0, +, PEGB0
			10'd129 : rdata = 48'b000011101111111010100000000000000000000010000000;
			// PEs: 16, 19 -> 
			// srcs: (1171, 130)(3002) -9, (3013) -19 --> (3014) -28:PENB, PEGB3, +, 
			10'd130 : rdata = 48'b000011101111111011100000110000000000000000000000;
			// PEs: 17, 16 -> 16
			// srcs: (1181, 131)(3014) -28, (3037) -9 --> (3038) -37:ALU, PENB, +, PEGB0
			10'd131 : rdata = 48'b000010011111111111011111110000000000000010000000;
			// PEs: 16 -> 
			// srcs: (1431, 132)(2843) -10 --> (2843) -10:PENB, pass, 
			10'd132 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 16, 17 -> 16
			// srcs: (1438, 133)(2795) -21, (2843) -10 --> (2844) -31:PENB, ALU, +, PEGB0
			10'd133 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 16, 17 -> 18
			// srcs: (1527, 134)(3140) 47, (23) -3 --> (3160) -141:PENB, ND0, *, PENB
			10'd134 : rdata = 48'b000111101111111001100000000000000000000100000000;
			// PEs: 17, 18 -> 17
			// srcs: (1536, 148)(808) -3, (3944) -141 --> (4728) 138:NW0, PEGB2, -, NW0
			10'd135 : rdata = 48'b000100100000000011100000100000000100000000000000;
			// PEs: 16, 17 -> 18
			// srcs: (1608, 135)(3140) 47, (104) 0 --> (3241) 0:PENB, ND1, *, PENB
			10'd136 : rdata = 48'b000111101111111001100000001000000000000100000000;
			// PEs: 16, 17 -> 18
			// srcs: (1612, 136)(3140) 47, (108) 2 --> (3245) 94:PENB, ND10, *, PENB
			10'd137 : rdata = 48'b000111101111111001100001010000000000000100000000;
			// PEs: 17, 18 -> 17
			// srcs: (1617, 149)(889) -1, (4025) 0 --> (4809) -1:NW1, PEGB2, -, NW1
			10'd138 : rdata = 48'b000100100000000111100000100000000100010000000000;
			// PEs: 17, 18 -> 17
			// srcs: (1621, 150)(893) 0, (4029) 94 --> (4813) -94:NW10, PEGB2, -, NW10
			10'd139 : rdata = 48'b000100100000101011100000100000000110100000000000;
			// PEs: 16, 17 -> 18
			// srcs: (1689, 137)(3140) 47, (185) 0 --> (3322) 0:PENB, ND2, *, PENB
			10'd140 : rdata = 48'b000111101111111001100000010000000000000100000000;
			// PEs: 17, 18 -> 17
			// srcs: (1698, 151)(970) 2, (4106) 0 --> (4890) 2:NW2, PEGB2, -, NW2
			10'd141 : rdata = 48'b000100100000001011100000100000000100100000000000;
			// PEs: 16, 17 -> 18
			// srcs: (1769, 138)(3140) 47, (265) 0 --> (3402) 0:PENB, ND3, *, PENB
			10'd142 : rdata = 48'b000111101111111001100000011000000000000100000000;
			// PEs: 17, 18 -> 17
			// srcs: (1778, 152)(1050) -3, (4186) 0 --> (4970) -3:NW3, PEGB2, -, NW3
			10'd143 : rdata = 48'b000100100000001111100000100000000100110000000000;
			// PEs: 16, 17 -> 18
			// srcs: (1792, 139)(3140) 47, (288) 1 --> (3425) 47:PENB, ND11, *, PENB
			10'd144 : rdata = 48'b000111101111111001100001011000000000000100000000;
			// PEs: 17, 18 -> 17
			// srcs: (1801, 153)(1073) -2, (4209) 47 --> (4993) -49:NW11, PEGB2, -, NW11
			10'd145 : rdata = 48'b000100100000101111100000100000000110110000000000;
			// PEs: 16, 17 -> 18
			// srcs: (1851, 140)(3140) 47, (347) 1 --> (3484) 47:PENB, ND4, *, PENB
			10'd146 : rdata = 48'b000111101111111001100000100000000000000100000000;
			// PEs: 17, 18 -> 17
			// srcs: (1860, 154)(1132) 2, (4268) 47 --> (5052) -45:NW4, PEGB2, -, NW4
			10'd147 : rdata = 48'b000100100000010011100000100000000101000000000000;
			// PEs: 16, 17 -> 18
			// srcs: (1931, 141)(3140) 47, (427) -3 --> (3564) -141:PENB, ND5, *, PENB
			10'd148 : rdata = 48'b000111101111111001100000101000000000000100000000;
			// PEs: 17, 18 -> 17
			// srcs: (1940, 155)(1212) -1, (4348) -141 --> (5132) 140:NW5, PEGB2, -, NW5
			10'd149 : rdata = 48'b000100100000010111100000100000000101010000000000;
			// PEs: 16, 17 -> 18
			// srcs: (1976, 142)(3140) 47, (472) -1 --> (3609) -47:PENB, ND12, *, PENB
			10'd150 : rdata = 48'b000111101111111001100001100000000000000100000000;
			// PEs: 17, 18 -> 17
			// srcs: (1985, 156)(1257) -2, (4393) -47 --> (5177) 45:NW12, PEGB2, -, NW12
			10'd151 : rdata = 48'b000100100000110011100000100000000111000000000000;
			// PEs: 16, 17 -> 18
			// srcs: (2011, 143)(3140) 47, (507) -3 --> (3644) -141:PENB, ND6, *, PENB
			10'd152 : rdata = 48'b000111101111111001100000110000000000000100000000;
			// PEs: 17, 18 -> 17
			// srcs: (2020, 157)(1292) 0, (4428) -141 --> (5212) 141:NW6, PEGB2, -, NW6
			10'd153 : rdata = 48'b000100100000011011100000100000000101100000000000;
			// PEs: 16, 17 -> 18
			// srcs: (2093, 144)(3140) 47, (589) 1 --> (3726) 47:PENB, ND7, *, PENB
			10'd154 : rdata = 48'b000111101111111001100000111000000000000100000000;
			// PEs: 17, 18 -> 17
			// srcs: (2102, 158)(1374) 0, (4510) 47 --> (5294) -47:NW7, PEGB2, -, NW7
			10'd155 : rdata = 48'b000100100000011111100000100000000101110000000000;
			// PEs: 16, 17 -> 18
			// srcs: (2160, 145)(3140) 47, (656) -1 --> (3793) -47:PENB, ND13, *, PENB
			10'd156 : rdata = 48'b000111101111111001100001101000000000000100000000;
			// PEs: 17, 18 -> 17
			// srcs: (2169, 159)(1441) 2, (4577) -47 --> (5361) 49:NW13, PEGB2, -, NW13
			10'd157 : rdata = 48'b000100100000110111100000100000000111010000000000;
			// PEs: 16, 17 -> 18
			// srcs: (2173, 146)(3140) 47, (669) 1 --> (3806) 47:PENB, ND8, *, PENB
			10'd158 : rdata = 48'b000111101111111001100001000000000000000100000000;
			// PEs: 17, 18 -> 17
			// srcs: (2182, 160)(1454) -1, (4590) 47 --> (5374) -48:NW8, PEGB2, -, NW8
			10'd159 : rdata = 48'b000100100000100011100000100000000110000000000000;
			// PEs: 16, 17 -> 18
			// srcs: (2253, 147)(3140) 47, (749) 1 --> (3886) 47:PENB, ND9, *, PENB
			10'd160 : rdata = 48'b000111101111111001100001001000000000000100000000;
			// PEs: 17, 18 -> 17
			// srcs: (2262, 161)(1534) 2, (4670) 47 --> (5454) -45:NW9, PEGB2, -, NW9
			10'd161 : rdata = 48'b000100100000100111100000100000000110010000000000;
			default : rdata = 48'b000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 18) begin
	always @(*) begin
		case(address)
			// PEs: 18, 18 -> 16
			// srcs: (1, 0)(24) -3, (809) 1 --> (1593) -3:ND0, NW0, *, PEGB0
			10'd0 : rdata = 48'b000110110000000001000000000000000000000010000000;
			// PEs: 18, 18 -> 18
			// srcs: (2, 1)(105) 0, (890) -2 --> (1674) 0:ND1, NW1, *, NI0
			10'd1 : rdata = 48'b000110110000000101000000001100000000000000000000;
			// PEs: 18, 18 -> 16
			// srcs: (3, 2)(186) -2, (971) 2 --> (1755) -4:ND2, NW2, *, PEGB0
			10'd2 : rdata = 48'b000110110000001001000000010000000000000010000000;
			// PEs: 18, 18 -> 16
			// srcs: (4, 3)(266) 1, (1051) -2 --> (1835) -2:ND3, NW3, *, PEGB0
			10'd3 : rdata = 48'b000110110000001101000000011000000000000010000000;
			// PEs: 18, 18 -> 18
			// srcs: (5, 4)(348) 0, (1133) -2 --> (1917) 0:ND4, NW4, *, NI1
			10'd4 : rdata = 48'b000110110000010001000000100100001000000000000000;
			// PEs: 18, 18 -> 16
			// srcs: (6, 5)(428) -3, (1213) 2 --> (1997) -6:ND5, NW5, *, PEGB0
			10'd5 : rdata = 48'b000110110000010101000000101000000000000010000000;
			// PEs: 18, 18 -> 16
			// srcs: (7, 6)(508) -1, (1293) -1 --> (2077) 1:ND6, NW6, *, PEGB0
			10'd6 : rdata = 48'b000110110000011001000000110000000000000010000000;
			// PEs: 18, 18 -> 16
			// srcs: (8, 7)(590) 1, (1375) -3 --> (2159) -3:ND7, NW7, *, PEGB0
			10'd7 : rdata = 48'b000110110000011101000000111000000000000010000000;
			// PEs: 18, 18 -> 19
			// srcs: (9, 8)(670) 2, (1455) -2 --> (2239) -4:ND8, NW8, *, PENB
			10'd8 : rdata = 48'b000110110000100001000001000000000000000100000000;
			// PEs: 18, 18 -> 21
			// srcs: (10, 9)(750) 0, (1535) 0 --> (2319) 0:ND9, NW9, *, PEGB5
			10'd9 : rdata = 48'b000110110000100101000001001000000000000011010000;
			// PEs: 18, 18 -> 18
			// srcs: (11, 10)(111) -1, (896) -3 --> (1680) 3:ND10, NW10, *, NI2
			10'd10 : rdata = 48'b000110110000101001000001010100010000000000000000;
			// PEs: 18, 18 -> 18
			// srcs: (12, 11)(291) -1, (1076) 0 --> (1860) 0:ND11, NW11, *, NI3
			10'd11 : rdata = 48'b000110110000101101000001011100011000000000000000;
			// PEs: 18, 18 -> 18
			// srcs: (13, 12)(475) 0, (1260) 2 --> (2044) 0:ND12, NW12, *, NI4
			10'd12 : rdata = 48'b000110110000110001000001100100100000000000000000;
			// PEs: 18, 18 -> 17
			// srcs: (14, 13)(659) 0, (1444) 2 --> (2228) 0:ND13, NW13, *, PEGB1
			10'd13 : rdata = 48'b000110110000110101000001101000000000000010010000;
			// PEs: 20 -> 18
			// srcs: (15, 18)(2242) 1 --> (2242) 1:PEGB4, pass, NI5
			10'd14 : rdata = 48'b110001110000100000000000000100101000000000000000;
			// PEs: 16 -> 18
			// srcs: (17, 14)(1578) -6 --> (1578) -6:PEGB0, pass, NI6
			10'd15 : rdata = 48'b110001110000000000000000000100110000000000000000;
			// PEs: 19, 18 -> 22
			// srcs: (18, 19)(2241) 0, (2242) 1 --> (3020) 1:PEGB3, NI5, +, PEGB6
			10'd16 : rdata = 48'b000011110000011010100000101000000000000011100000;
			// PEs: 16, 18 -> 16
			// srcs: (26, 15)(1577) -4, (1578) -6 --> (2360) -10:PEGB0, NI6, +, PEGB0
			10'd17 : rdata = 48'b000011110000000010100000110000000000000010000000;
			// PEs: 16 -> 
			// srcs: (57, 16)(1749) 2 --> (1749) 2:PEGB0, pass, 
			10'd18 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 16, 18 -> 18
			// srcs: (66, 17)(1748) -3, (1749) 2 --> (2528) -1:PEGB0, ALU, +, NI5
			10'd19 : rdata = 48'b000011110000000000111111111100101000000000000000;
			// PEs: 18 -> 16
			// srcs: (118, 22)(1680) 3 --> (1680) 3:NI2, pass, PEGB0
			10'd20 : rdata = 48'b110001010000001000000000000000000000000010000000;
			// PEs: 18 -> 16
			// srcs: (120, 20)(1674) 0 --> (1674) 0:NI0, pass, PEGB0
			10'd21 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 18 -> 16
			// srcs: (128, 23)(2528) -1 --> (2528) -1:NI5, pass, PEGB0
			10'd22 : rdata = 48'b110001010000010100000000000000000000000010000000;
			// PEs: 18 -> 16
			// srcs: (129, 24)(1860) 0 --> (1860) 0:NI3, pass, PEGB0
			10'd23 : rdata = 48'b110001010000001100000000000000000000000010000000;
			// PEs: 18 -> 16
			// srcs: (136, 21)(1917) 0 --> (1917) 0:NI1, pass, PEGB0
			10'd24 : rdata = 48'b110001010000000100000000000000000000000010000000;
			// PEs: 18 -> 16
			// srcs: (210, 25)(2044) 0 --> (2044) 0:NI4, pass, PEGB0
			10'd25 : rdata = 48'b110001010000010000000000000000000000000010000000;
			// PEs: 17 -> 
			// srcs: (399, 26)(3006) 1 --> (3006) 1:PENB, pass, 
			10'd26 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 17, 18 -> 18
			// srcs: (406, 27)(3004) -2, (3006) 1 --> (3007) -1:PENB, ALU, +, NI0
			10'd27 : rdata = 48'b000011101111111000111111111100000000000000000000;
			// PEs: 17 -> 
			// srcs: (568, 28)(3011) -4 --> (3011) -4:PENB, pass, 
			10'd28 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 17, 18 -> 19
			// srcs: (575, 29)(3009) -14, (3011) -4 --> (3012) -18:PENB, ALU, +, PENB
			10'd29 : rdata = 48'b000011101111111000111111111000000000000100000000;
			// PEs: 18 -> 19
			// srcs: (582, 30)(3007) -1 --> (3007) -1:NI0, pass, PENB
			10'd30 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 18, 17 -> 17
			// srcs: (1530, 45)(3) 1, (3160) -141 --> (3944) -141:NM0, PENB, *, PEGB1
			10'd31 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 16, 18 -> 19
			// srcs: (1531, 31)(3140) 47, (24) -3 --> (3161) -141:PEGB0, ND0, *, PENB
			10'd32 : rdata = 48'b000111110000000001100000000000000000000100000000;
			// PEs: 18, 19 -> 18
			// srcs: (1540, 63)(809) 1, (3945) -141 --> (4729) 142:NW0, PEGB3, -, NW0
			10'd33 : rdata = 48'b000100100000000011100000110000000100000000000000;
			// PEs: 18, 17 -> 17
			// srcs: (1611, 46)(3) 1, (3241) 0 --> (4025) 0:NM0, PENB, *, PEGB1
			10'd34 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 16, 18 -> 19
			// srcs: (1612, 32)(3140) 47, (105) 0 --> (3242) 0:PEGB0, ND1, *, PENB
			10'd35 : rdata = 48'b000111110000000001100000001000000000000100000000;
			// PEs: 18, 17 -> 17
			// srcs: (1615, 47)(3) 1, (3245) 94 --> (4029) 94:NM0, PENB, *, PEGB1
			10'd36 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 16, 18 -> 
			// srcs: (1618, 33)(3140) 47, (111) -1 --> (3248) -47:PEGB0, ND10, *, 
			10'd37 : rdata = 48'b000111110000000001100001010000000000000000000000;
			// PEs: 18, 18 -> 18
			// srcs: (1621, 48)(3) 1, (3248) -47 --> (4032) -47:NM0, ALU, *, NI0
			10'd38 : rdata = 48'b000111000000000000111111111100000000000000000000;
			// PEs: 18, 19 -> 18
			// srcs: (1622, 64)(890) -2, (4026) 0 --> (4810) -2:NW1, PEGB3, -, NW1
			10'd39 : rdata = 48'b000100100000000111100000110000000100010000000000;
			// PEs: 18, 18 -> 18
			// srcs: (1624, 65)(896) -3, (4032) -47 --> (4816) 44:NW10, NI0, -, NW10
			10'd40 : rdata = 48'b000100100000101010100000000000000110100000000000;
			// PEs: 18, 17 -> 17
			// srcs: (1692, 49)(3) 1, (3322) 0 --> (4106) 0:NM0, PENB, *, PEGB1
			10'd41 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 16, 18 -> 19
			// srcs: (1693, 34)(3140) 47, (186) -2 --> (3323) -94:PEGB0, ND2, *, PENB
			10'd42 : rdata = 48'b000111110000000001100000010000000000000100000000;
			// PEs: 18, 19 -> 18
			// srcs: (1702, 66)(971) 2, (4107) -94 --> (4891) 96:NW2, PEGB3, -, NW2
			10'd43 : rdata = 48'b000100100000001011100000110000000100100000000000;
			// PEs: 18, 17 -> 17
			// srcs: (1772, 50)(3) 1, (3402) 0 --> (4186) 0:NM0, PENB, *, PEGB1
			10'd44 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 16, 18 -> 19
			// srcs: (1773, 35)(3140) 47, (266) 1 --> (3403) 47:PEGB0, ND3, *, PENB
			10'd45 : rdata = 48'b000111110000000001100000011000000000000100000000;
			// PEs: 18, 19 -> 18
			// srcs: (1782, 67)(1051) -2, (4187) 47 --> (4971) -49:NW3, PEGB3, -, NW3
			10'd46 : rdata = 48'b000100100000001111100000110000000100110000000000;
			// PEs: 18, 17 -> 17
			// srcs: (1795, 51)(3) 1, (3425) 47 --> (4209) 47:NM0, PENB, *, PEGB1
			10'd47 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 16, 18 -> 
			// srcs: (1798, 36)(3140) 47, (291) -1 --> (3428) -47:PEGB0, ND11, *, 
			10'd48 : rdata = 48'b000111110000000001100001011000000000000000000000;
			// PEs: 18, 18 -> 
			// srcs: (1801, 52)(3) 1, (3428) -47 --> (4212) -47:NM0, ALU, *, 
			10'd49 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 18, 18 -> 18
			// srcs: (1804, 68)(1076) 0, (4212) -47 --> (4996) 47:NW11, ALU, -, NW11
			10'd50 : rdata = 48'b000100100000101100111111111000000110110000000000;
			// PEs: 18, 17 -> 17
			// srcs: (1854, 53)(3) 1, (3484) 47 --> (4268) 47:NM0, PENB, *, PEGB1
			10'd51 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 16, 18 -> 19
			// srcs: (1855, 37)(3140) 47, (348) 0 --> (3485) 0:PEGB0, ND4, *, PENB
			10'd52 : rdata = 48'b000111110000000001100000100000000000000100000000;
			// PEs: 18, 19 -> 18
			// srcs: (1864, 69)(1133) -2, (4269) 0 --> (5053) -2:NW4, PEGB3, -, NW4
			10'd53 : rdata = 48'b000100100000010011100000110000000101000000000000;
			// PEs: 18, 17 -> 17
			// srcs: (1934, 54)(3) 1, (3564) -141 --> (4348) -141:NM0, PENB, *, PEGB1
			10'd54 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 16, 18 -> 19
			// srcs: (1935, 38)(3140) 47, (428) -3 --> (3565) -141:PEGB0, ND5, *, PENB
			10'd55 : rdata = 48'b000111110000000001100000101000000000000100000000;
			// PEs: 18, 19 -> 18
			// srcs: (1944, 70)(1213) 2, (4349) -141 --> (5133) 143:NW5, PEGB3, -, NW5
			10'd56 : rdata = 48'b000100100000010111100000110000000101010000000000;
			// PEs: 18, 17 -> 17
			// srcs: (1979, 55)(3) 1, (3609) -47 --> (4393) -47:NM0, PENB, *, PEGB1
			10'd57 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 16, 18 -> 
			// srcs: (1982, 39)(3140) 47, (475) 0 --> (3612) 0:PEGB0, ND12, *, 
			10'd58 : rdata = 48'b000111110000000001100001100000000000000000000000;
			// PEs: 18, 18 -> 
			// srcs: (1985, 56)(3) 1, (3612) 0 --> (4396) 0:NM0, ALU, *, 
			10'd59 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 18, 18 -> 18
			// srcs: (1988, 71)(1260) 2, (4396) 0 --> (5180) 2:NW12, ALU, -, NW12
			10'd60 : rdata = 48'b000100100000110000111111111000000111000000000000;
			// PEs: 18, 17 -> 17
			// srcs: (2014, 57)(3) 1, (3644) -141 --> (4428) -141:NM0, PENB, *, PEGB1
			10'd61 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 16, 18 -> 19
			// srcs: (2015, 40)(3140) 47, (508) -1 --> (3645) -47:PEGB0, ND6, *, PENB
			10'd62 : rdata = 48'b000111110000000001100000110000000000000100000000;
			// PEs: 18, 19 -> 18
			// srcs: (2024, 72)(1293) -1, (4429) -47 --> (5213) 46:NW6, PEGB3, -, NW6
			10'd63 : rdata = 48'b000100100000011011100000110000000101100000000000;
			// PEs: 18, 17 -> 17
			// srcs: (2096, 58)(3) 1, (3726) 47 --> (4510) 47:NM0, PENB, *, PEGB1
			10'd64 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 16, 18 -> 19
			// srcs: (2097, 41)(3140) 47, (590) 1 --> (3727) 47:PEGB0, ND7, *, PENB
			10'd65 : rdata = 48'b000111110000000001100000111000000000000100000000;
			// PEs: 18, 19 -> 18
			// srcs: (2106, 73)(1375) -3, (4511) 47 --> (5295) -50:NW7, PEGB3, -, NW7
			10'd66 : rdata = 48'b000100100000011111100000110000000101110000000000;
			// PEs: 18, 17 -> 17
			// srcs: (2163, 59)(3) 1, (3793) -47 --> (4577) -47:NM0, PENB, *, PEGB1
			10'd67 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 16, 18 -> 
			// srcs: (2166, 42)(3140) 47, (659) 0 --> (3796) 0:PEGB0, ND13, *, 
			10'd68 : rdata = 48'b000111110000000001100001101000000000000000000000;
			// PEs: 18, 18 -> 
			// srcs: (2169, 60)(3) 1, (3796) 0 --> (4580) 0:NM0, ALU, *, 
			10'd69 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 18, 18 -> 18
			// srcs: (2172, 74)(1444) 2, (4580) 0 --> (5364) 2:NW13, ALU, -, NW13
			10'd70 : rdata = 48'b000100100000110100111111111000000111010000000000;
			// PEs: 18, 17 -> 17
			// srcs: (2176, 61)(3) 1, (3806) 47 --> (4590) 47:NM0, PENB, *, PEGB1
			10'd71 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 16, 18 -> 19
			// srcs: (2177, 43)(3140) 47, (670) 2 --> (3807) 94:PEGB0, ND8, *, PENB
			10'd72 : rdata = 48'b000111110000000001100001000000000000000100000000;
			// PEs: 18, 19 -> 18
			// srcs: (2186, 75)(1455) -2, (4591) 94 --> (5375) -96:NW8, PEGB3, -, NW8
			10'd73 : rdata = 48'b000100100000100011100000110000000110000000000000;
			// PEs: 18, 17 -> 17
			// srcs: (2256, 62)(3) 1, (3886) 47 --> (4670) 47:NM0, PENB, *, PEGB1
			10'd74 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 16, 18 -> 19
			// srcs: (2257, 44)(3140) 47, (750) 0 --> (3887) 0:PEGB0, ND9, *, PENB
			10'd75 : rdata = 48'b000111110000000001100001001000000000000100000000;
			// PEs: 18, 19 -> 18
			// srcs: (2266, 76)(1535) 0, (4671) 0 --> (5455) 0:NW9, PEGB3, -, NW9
			10'd76 : rdata = 48'b000100100000100111100000110000000110010000000000;
			default : rdata = 48'b000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 19) begin
	always @(*) begin
		case(address)
			// PEs: 19, 19 -> 16
			// srcs: (1, 0)(26) 0, (811) -2 --> (1595) 0:ND0, NW0, *, PEGB0
			10'd0 : rdata = 48'b000110110000000001000000000000000000000010000000;
			// PEs: 19, 19 -> 16
			// srcs: (2, 1)(106) -2, (891) -2 --> (1675) 4:ND1, NW1, *, PEGB0
			10'd1 : rdata = 48'b000110110000000101000000001000000000000010000000;
			// PEs: 19, 19 -> 16
			// srcs: (3, 2)(188) 2, (973) -2 --> (1757) -4:ND2, NW2, *, PEGB0
			10'd2 : rdata = 48'b000110110000001001000000010000000000000010000000;
			// PEs: 19, 19 -> 16
			// srcs: (4, 3)(268) -1, (1053) -1 --> (1837) 1:ND3, NW3, *, PEGB0
			10'd3 : rdata = 48'b000110110000001101000000011000000000000010000000;
			// PEs: 19, 19 -> 19
			// srcs: (5, 4)(349) -1, (1134) -1 --> (1918) 1:ND4, NW4, *, NI0
			10'd4 : rdata = 48'b000110110000010001000000100100000000000000000000;
			// PEs: 19, 19 -> 16
			// srcs: (6, 5)(430) -2, (1215) -1 --> (1999) 2:ND5, NW5, *, PEGB0
			10'd5 : rdata = 48'b000110110000010101000000101000000000000010000000;
			// PEs: 19, 19 -> 16
			// srcs: (7, 6)(510) 1, (1295) 0 --> (2079) 0:ND6, NW6, *, PEGB0
			10'd6 : rdata = 48'b000110110000011001000000110000000000000010000000;
			// PEs: 19, 19 -> 19
			// srcs: (8, 7)(592) 0, (1377) 2 --> (2161) 0:ND7, NW7, *, NI1
			10'd7 : rdata = 48'b000110110000011101000000111100001000000000000000;
			// PEs: 19, 19 -> 18
			// srcs: (9, 8)(672) 2, (1457) 0 --> (2241) 0:ND8, NW8, *, PEGB2
			10'd8 : rdata = 48'b000110110000100001000001000000000000000010100000;
			// PEs: 19, 19 -> 22
			// srcs: (10, 9)(752) 2, (1537) -1 --> (2321) -2:ND9, NW9, *, PEGB6
			10'd9 : rdata = 48'b000110110000100101000001001000000000000011100000;
			// PEs: 19, 19 -> 16
			// srcs: (11, 10)(114) 1, (899) 1 --> (1683) 1:ND10, NW10, *, PEGB0
			10'd10 : rdata = 48'b000110110000101001000001010000000000000010000000;
			// PEs: 19, 19 -> 19
			// srcs: (12, 11)(294) -2, (1079) -3 --> (1863) 6:ND11, NW11, *, NI2
			10'd11 : rdata = 48'b000110110000101101000001011100010000000000000000;
			// PEs: 19, 19 -> 19
			// srcs: (13, 12)(478) 2, (1263) -2 --> (2047) -4:ND12, NW12, *, NI3
			10'd12 : rdata = 48'b000110110000110001000001100100011000000000000000;
			// PEs: 19, 19 -> 19
			// srcs: (14, 13)(662) 1, (1447) -2 --> (2231) -2:ND13, NW13, *, NI4
			10'd13 : rdata = 48'b000110110000110101000001101100100000000000000000;
			// PEs: 17, 18 -> 21
			// srcs: (15, 18)(2238) -1, (2239) -4 --> (3017) -5:PEGB1, PENB, +, PEGB5
			10'd14 : rdata = 48'b000011110000001011011111110000000000000011010000;
			// PEs: 16 -> 
			// srcs: (21, 14)(1617) -4 --> (1617) -4:PEGB0, pass, 
			10'd15 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 16, 19 -> 17
			// srcs: (30, 15)(1616) 0, (1617) -4 --> (2397) -4:PEGB0, ALU, +, PEGB1
			10'd16 : rdata = 48'b000011110000000000111111111000000000000010010000;
			// PEs: 16 -> 
			// srcs: (60, 16)(1752) 2 --> (1752) 2:PEGB0, pass, 
			10'd17 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 16, 19 -> 19
			// srcs: (69, 17)(1751) 0, (1752) 2 --> (2531) 2:PEGB0, ALU, +, NI5
			10'd18 : rdata = 48'b000011110000000000111111111100101000000000000000;
			// PEs: 19 -> 16
			// srcs: (144, 19)(1918) 1 --> (1918) 1:NI0, pass, PEGB0
			10'd19 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 19 -> 16
			// srcs: (160, 20)(2161) 0 --> (2161) 0:NI1, pass, PEGB0
			10'd20 : rdata = 48'b110001010000000100000000000000000000000010000000;
			// PEs: 19 -> 16
			// srcs: (193, 21)(2531) 2 --> (2531) 2:NI5, pass, PEGB0
			10'd21 : rdata = 48'b110001010000010100000000000000000000000010000000;
			// PEs: 19 -> 16
			// srcs: (218, 23)(2047) -4 --> (2047) -4:NI3, pass, PEGB0
			10'd22 : rdata = 48'b110001010000001100000000000000000000000010000000;
			// PEs: 19 -> 16
			// srcs: (277, 22)(1863) 6 --> (1863) 6:NI2, pass, PEGB0
			10'd23 : rdata = 48'b110001010000001000000000000000000000000010000000;
			// PEs: 19 -> 17
			// srcs: (553, 24)(2231) -2 --> (2231) -2:NI4, pass, PEGB1
			10'd24 : rdata = 48'b110001010000010000000000000000000000000010010000;
			// PEs: 18 -> 
			// srcs: (577, 25)(3012) -18 --> (3012) -18:PENB, pass, 
			10'd25 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 18, 19 -> 17
			// srcs: (584, 26)(3007) -1, (3012) -18 --> (3013) -19:PENB, ALU, +, PEGB1
			10'd26 : rdata = 48'b000011101111111000111111111000000000000010010000;
			// PEs: 16, 19 -> 20
			// srcs: (1533, 27)(3140) 47, (26) 0 --> (3163) 0:PEGB0, ND0, *, PENB
			10'd27 : rdata = 48'b000111110000000001100000000000000000000100000000;
			// PEs: 19, 18 -> 18
			// srcs: (1534, 41)(3) 1, (3161) -141 --> (3945) -141:NM0, PENB, *, PEGB2
			10'd28 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 19, 20 -> 19
			// srcs: (1542, 56)(811) -2, (3947) 0 --> (4731) -2:NW0, PEGB4, -, NW0
			10'd29 : rdata = 48'b000100100000000011100001000000000100000000000000;
			// PEs: 16, 19 -> 20
			// srcs: (1613, 28)(3140) 47, (106) -2 --> (3243) -94:PEGB0, ND1, *, PENB
			10'd30 : rdata = 48'b000111110000000001100000001000000000000100000000;
			// PEs: 19, 18 -> 18
			// srcs: (1615, 42)(3) 1, (3242) 0 --> (4026) 0:NM0, PENB, *, PEGB2
			10'd31 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 16, 19 -> 19
			// srcs: (1621, 29)(3140) 47, (114) 1 --> (3251) 47:PEGB0, ND10, *, NI0
			10'd32 : rdata = 48'b000111110000000001100001010100000000000000000000;
			// PEs: 19, 20 -> 19
			// srcs: (1622, 57)(891) -2, (4027) -94 --> (4811) 92:NW1, PEGB4, -, NW1
			10'd33 : rdata = 48'b000100100000000111100001000000000100010000000000;
			// PEs: 19, 19 -> 
			// srcs: (1624, 43)(3) 1, (3251) 47 --> (4035) 47:NM0, NI0, *, 
			10'd34 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 19, 19 -> 19
			// srcs: (1627, 58)(899) 1, (4035) 47 --> (4819) -46:NW10, ALU, -, NW10
			10'd35 : rdata = 48'b000100100000101000111111111000000110100000000000;
			// PEs: 16, 19 -> 20
			// srcs: (1695, 30)(3140) 47, (188) 2 --> (3325) 94:PEGB0, ND2, *, PENB
			10'd36 : rdata = 48'b000111110000000001100000010000000000000100000000;
			// PEs: 19, 18 -> 18
			// srcs: (1696, 44)(3) 1, (3323) -94 --> (4107) -94:NM0, PENB, *, PEGB2
			10'd37 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 19, 20 -> 19
			// srcs: (1704, 59)(973) -2, (4109) 94 --> (4893) -96:NW2, PEGB4, -, NW2
			10'd38 : rdata = 48'b000100100000001011100001000000000100100000000000;
			// PEs: 16, 19 -> 20
			// srcs: (1775, 31)(3140) 47, (268) -1 --> (3405) -47:PEGB0, ND3, *, PENB
			10'd39 : rdata = 48'b000111110000000001100000011000000000000100000000;
			// PEs: 19, 18 -> 18
			// srcs: (1776, 45)(3) 1, (3403) 47 --> (4187) 47:NM0, PENB, *, PEGB2
			10'd40 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 19, 20 -> 19
			// srcs: (1784, 60)(1053) -1, (4189) -47 --> (4973) 46:NW3, PEGB4, -, NW3
			10'd41 : rdata = 48'b000100100000001111100001000000000100110000000000;
			// PEs: 16, 19 -> 
			// srcs: (1801, 32)(3140) 47, (294) -2 --> (3431) -94:PEGB0, ND11, *, 
			10'd42 : rdata = 48'b000111110000000001100001011000000000000000000000;
			// PEs: 19, 19 -> 
			// srcs: (1804, 46)(3) 1, (3431) -94 --> (4215) -94:NM0, ALU, *, 
			10'd43 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 19, 19 -> 19
			// srcs: (1807, 61)(1079) -3, (4215) -94 --> (4999) 91:NW11, ALU, -, NW11
			10'd44 : rdata = 48'b000100100000101100111111111000000110110000000000;
			// PEs: 16, 19 -> 20
			// srcs: (1856, 33)(3140) 47, (349) -1 --> (3486) -47:PEGB0, ND4, *, PENB
			10'd45 : rdata = 48'b000111110000000001100000100000000000000100000000;
			// PEs: 19, 18 -> 18
			// srcs: (1858, 47)(3) 1, (3485) 0 --> (4269) 0:NM0, PENB, *, PEGB2
			10'd46 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 19, 20 -> 19
			// srcs: (1865, 62)(1134) -1, (4270) -47 --> (5054) 46:NW4, PEGB4, -, NW4
			10'd47 : rdata = 48'b000100100000010011100001000000000101000000000000;
			// PEs: 16, 19 -> 20
			// srcs: (1937, 34)(3140) 47, (430) -2 --> (3567) -94:PEGB0, ND5, *, PENB
			10'd48 : rdata = 48'b000111110000000001100000101000000000000100000000;
			// PEs: 19, 18 -> 18
			// srcs: (1938, 48)(3) 1, (3565) -141 --> (4349) -141:NM0, PENB, *, PEGB2
			10'd49 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 19, 20 -> 19
			// srcs: (1946, 63)(1215) -1, (4351) -94 --> (5135) 93:NW5, PEGB4, -, NW5
			10'd50 : rdata = 48'b000100100000010111100001000000000101010000000000;
			// PEs: 16, 19 -> 
			// srcs: (1985, 35)(3140) 47, (478) 2 --> (3615) 94:PEGB0, ND12, *, 
			10'd51 : rdata = 48'b000111110000000001100001100000000000000000000000;
			// PEs: 19, 19 -> 
			// srcs: (1988, 49)(3) 1, (3615) 94 --> (4399) 94:NM0, ALU, *, 
			10'd52 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 19, 19 -> 19
			// srcs: (1991, 64)(1263) -2, (4399) 94 --> (5183) -96:NW12, ALU, -, NW12
			10'd53 : rdata = 48'b000100100000110000111111111000000111000000000000;
			// PEs: 16, 19 -> 20
			// srcs: (2017, 36)(3140) 47, (510) 1 --> (3647) 47:PEGB0, ND6, *, PENB
			10'd54 : rdata = 48'b000111110000000001100000110000000000000100000000;
			// PEs: 19, 18 -> 18
			// srcs: (2018, 50)(3) 1, (3645) -47 --> (4429) -47:NM0, PENB, *, PEGB2
			10'd55 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 19, 20 -> 19
			// srcs: (2026, 65)(1295) 0, (4431) 47 --> (5215) -47:NW6, PEGB4, -, NW6
			10'd56 : rdata = 48'b000100100000011011100001000000000101100000000000;
			// PEs: 16, 19 -> 20
			// srcs: (2099, 37)(3140) 47, (592) 0 --> (3729) 0:PEGB0, ND7, *, PENB
			10'd57 : rdata = 48'b000111110000000001100000111000000000000100000000;
			// PEs: 19, 18 -> 18
			// srcs: (2100, 51)(3) 1, (3727) 47 --> (4511) 47:NM0, PENB, *, PEGB2
			10'd58 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 19, 20 -> 19
			// srcs: (2108, 66)(1377) 2, (4513) 0 --> (5297) 2:NW7, PEGB4, -, NW7
			10'd59 : rdata = 48'b000100100000011111100001000000000101110000000000;
			// PEs: 16, 19 -> 
			// srcs: (2169, 38)(3140) 47, (662) 1 --> (3799) 47:PEGB0, ND13, *, 
			10'd60 : rdata = 48'b000111110000000001100001101000000000000000000000;
			// PEs: 19, 19 -> 
			// srcs: (2172, 52)(3) 1, (3799) 47 --> (4583) 47:NM0, ALU, *, 
			10'd61 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 19, 19 -> 19
			// srcs: (2175, 67)(1447) -2, (4583) 47 --> (5367) -49:NW13, ALU, -, NW13
			10'd62 : rdata = 48'b000100100000110100111111111000000111010000000000;
			// PEs: 16, 19 -> 19
			// srcs: (2179, 39)(3140) 47, (672) 2 --> (3809) 94:PEGB0, ND8, *, NI0
			10'd63 : rdata = 48'b000111110000000001100001000100000000000000000000;
			// PEs: 19, 18 -> 18
			// srcs: (2180, 53)(3) 1, (3807) 94 --> (4591) 94:NM0, PENB, *, PEGB2
			10'd64 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 19, 19 -> 
			// srcs: (2182, 54)(3) 1, (3809) 94 --> (4593) 94:NM0, NI0, *, 
			10'd65 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 19, 19 -> 19
			// srcs: (2185, 68)(1457) 0, (4593) 94 --> (5377) -94:NW8, ALU, -, NW8
			10'd66 : rdata = 48'b000100100000100000111111111000000110000000000000;
			// PEs: 16, 19 -> 20
			// srcs: (2259, 40)(3140) 47, (752) 2 --> (3889) 94:PEGB0, ND9, *, PENB
			10'd67 : rdata = 48'b000111110000000001100001001000000000000100000000;
			// PEs: 19, 18 -> 18
			// srcs: (2260, 55)(3) 1, (3887) 0 --> (4671) 0:NM0, PENB, *, PEGB2
			10'd68 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 19, 20 -> 19
			// srcs: (2268, 69)(1537) -1, (4673) 94 --> (5457) -95:NW9, PEGB4, -, NW9
			10'd69 : rdata = 48'b000100100000100111100001000000000110010000000000;
			default : rdata = 48'b000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 20) begin
	always @(*) begin
		case(address)
			// PEs: 20, 20 -> 16
			// srcs: (1, 0)(27) -3, (812) 2 --> (1596) -6:ND0, NW0, *, PEGB0
			10'd0 : rdata = 48'b000110110000000001000000000000000000000010000000;
			// PEs: 20, 20 -> 16
			// srcs: (2, 1)(107) 2, (892) -3 --> (1676) -6:ND1, NW1, *, PEGB0
			10'd1 : rdata = 48'b000110110000000101000000001000000000000010000000;
			// PEs: 20, 20 -> 16
			// srcs: (3, 2)(189) 0, (974) -2 --> (1758) 0:ND2, NW2, *, PEGB0
			10'd2 : rdata = 48'b000110110000001001000000010000000000000010000000;
			// PEs: 20, 20 -> 16
			// srcs: (4, 3)(269) -1, (1054) -3 --> (1838) 3:ND3, NW3, *, PEGB0
			10'd3 : rdata = 48'b000110110000001101000000011000000000000010000000;
			// PEs: 20, 20 -> 20
			// srcs: (5, 4)(350) 2, (1135) 2 --> (1919) 4:ND4, NW4, *, NI0
			10'd4 : rdata = 48'b000110110000010001000000100100000000000000000000;
			// PEs: 20, 20 -> 16
			// srcs: (6, 5)(431) -3, (1216) -2 --> (2000) 6:ND5, NW5, *, PEGB0
			10'd5 : rdata = 48'b000110110000010101000000101000000000000010000000;
			// PEs: 20, 20 -> 16
			// srcs: (7, 6)(511) 0, (1296) 1 --> (2080) 0:ND6, NW6, *, PEGB0
			10'd6 : rdata = 48'b000110110000011001000000110000000000000010000000;
			// PEs: 20, 20 -> 20
			// srcs: (8, 7)(593) 2, (1378) 2 --> (2162) 4:ND7, NW7, *, NI1
			10'd7 : rdata = 48'b000110110000011101000000111100001000000000000000;
			// PEs: 20, 20 -> 18
			// srcs: (9, 8)(673) 1, (1458) 1 --> (2242) 1:ND8, NW8, *, PEGB2
			10'd8 : rdata = 48'b000110110000100001000001000000000000000010100000;
			// PEs: 20, 20 -> 22
			// srcs: (10, 9)(753) -2, (1538) -2 --> (2322) 4:ND9, NW9, *, PEGB6
			10'd9 : rdata = 48'b000110110000100101000001001000000000000011100000;
			// PEs: 20, 20 -> 20
			// srcs: (11, 10)(117) 1, (902) -1 --> (1686) -1:ND10, NW10, *, NI2
			10'd10 : rdata = 48'b000110110000101001000001010100010000000000000000;
			// PEs: 20, 20 -> 20
			// srcs: (12, 11)(297) 1, (1082) -3 --> (1866) -3:ND11, NW11, *, NI3
			10'd11 : rdata = 48'b000110110000101101000001011100011000000000000000;
			// PEs: 20, 20 -> 20
			// srcs: (13, 12)(481) -1, (1266) 0 --> (2050) 0:ND12, NW12, *, NI4
			10'd12 : rdata = 48'b000110110000110001000001100100100000000000000000;
			// PEs: 20, 20 -> 17
			// srcs: (14, 13)(665) 0, (1450) 2 --> (2234) 0:ND13, NW13, *, PEGB1
			10'd13 : rdata = 48'b000110110000110101000001101000000000000010010000;
			// PEs: 22 -> 
			// srcs: (15, 18)(2245) -6 --> (2245) -6:PEGB6, pass, 
			10'd14 : rdata = 48'b110001110000110000000000000000000000000000000000;
			// PEs: 21, 20 -> 20
			// srcs: (17, 19)(2244) 4, (2245) -6 --> (3022) -2:PEGB5, ALU, +, NI5
			10'd15 : rdata = 48'b000011110000101000111111111100101000000000000000;
			// PEs: 16 -> 
			// srcs: (23, 14)(1620) 0 --> (1620) 0:PEGB0, pass, 
			10'd16 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 16, 20 -> 16
			// srcs: (32, 15)(1619) 0, (1620) 0 --> (2399) 0:PEGB0, ALU, +, PEGB0
			10'd17 : rdata = 48'b000011110000000000111111111000000000000010000000;
			// PEs: 16 -> 
			// srcs: (68, 16)(1823) 0 --> (1823) 0:PEGB0, pass, 
			10'd18 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 16, 20 -> 20
			// srcs: (77, 17)(1822) 0, (1823) 0 --> (2603) 0:PEGB0, ALU, +, NI6
			10'd19 : rdata = 48'b000011110000000000111111111100110000000000000000;
			// PEs: 20 -> 16
			// srcs: (152, 20)(1919) 4 --> (1919) 4:NI0, pass, PEGB0
			10'd20 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 20 -> 16
			// srcs: (168, 21)(2162) 4 --> (2162) 4:NI1, pass, PEGB0
			10'd21 : rdata = 48'b110001010000000100000000000000000000000010000000;
			// PEs: 20 -> 16
			// srcs: (194, 23)(2603) 0 --> (2603) 0:NI6, pass, PEGB0
			10'd22 : rdata = 48'b110001010000011000000000000000000000000010000000;
			// PEs: 20 -> 16
			// srcs: (202, 24)(1866) -3 --> (1866) -3:NI3, pass, PEGB0
			10'd23 : rdata = 48'b110001010000001100000000000000000000000010000000;
			// PEs: 20 -> 16
			// srcs: (205, 25)(2050) 0 --> (2050) 0:NI4, pass, PEGB0
			10'd24 : rdata = 48'b110001010000010000000000000000000000000010000000;
			// PEs: 20 -> 16
			// srcs: (264, 22)(1686) -1 --> (1686) -1:NI2, pass, PEGB0
			10'd25 : rdata = 48'b110001010000001000000000000000000000000010000000;
			// PEs: 20 -> 16
			// srcs: (338, 26)(3022) -2 --> (3022) -2:NI5, pass, PEGB0
			10'd26 : rdata = 48'b110001010000010100000000000000000000000010000000;
			// PEs: 16, 20 -> 21
			// srcs: (1534, 27)(3140) 47, (27) -3 --> (3164) -141:PEGB0, ND0, *, PENB
			10'd27 : rdata = 48'b000111110000000001100000000000000000000100000000;
			// PEs: 20, 19 -> 19
			// srcs: (1536, 41)(3) 1, (3163) 0 --> (3947) 0:NM0, PENB, *, PEGB3
			10'd28 : rdata = 48'b000111000000000011011111110000000000000010110000;
			// PEs: 20, 21 -> 20
			// srcs: (1543, 56)(812) 2, (3948) -141 --> (4732) 143:NW0, PEGB5, -, NW0
			10'd29 : rdata = 48'b000100100000000011100001010000000100000000000000;
			// PEs: 16, 20 -> 21
			// srcs: (1614, 28)(3140) 47, (107) 2 --> (3244) 94:PEGB0, ND1, *, PENB
			10'd30 : rdata = 48'b000111110000000001100000001000000000000100000000;
			// PEs: 20, 19 -> 19
			// srcs: (1616, 42)(3) 1, (3243) -94 --> (4027) -94:NM0, PENB, *, PEGB3
			10'd31 : rdata = 48'b000111000000000011011111110000000000000010110000;
			// PEs: 20, 21 -> 20
			// srcs: (1623, 57)(892) -3, (4028) 94 --> (4812) -97:NW1, PEGB5, -, NW1
			10'd32 : rdata = 48'b000100100000000111100001010000000100010000000000;
			// PEs: 16, 20 -> 
			// srcs: (1624, 29)(3140) 47, (117) 1 --> (3254) 47:PEGB0, ND10, *, 
			10'd33 : rdata = 48'b000111110000000001100001010000000000000000000000;
			// PEs: 20, 20 -> 
			// srcs: (1627, 43)(3) 1, (3254) 47 --> (4038) 47:NM0, ALU, *, 
			10'd34 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 20, 20 -> 20
			// srcs: (1630, 58)(902) -1, (4038) 47 --> (4822) -48:NW10, ALU, -, NW10
			10'd35 : rdata = 48'b000100100000101000111111111000000110100000000000;
			// PEs: 16, 20 -> 21
			// srcs: (1696, 30)(3140) 47, (189) 0 --> (3326) 0:PEGB0, ND2, *, PENB
			10'd36 : rdata = 48'b000111110000000001100000010000000000000100000000;
			// PEs: 20, 19 -> 19
			// srcs: (1698, 44)(3) 1, (3325) 94 --> (4109) 94:NM0, PENB, *, PEGB3
			10'd37 : rdata = 48'b000111000000000011011111110000000000000010110000;
			// PEs: 20, 21 -> 20
			// srcs: (1705, 59)(974) -2, (4110) 0 --> (4894) -2:NW2, PEGB5, -, NW2
			10'd38 : rdata = 48'b000100100000001011100001010000000100100000000000;
			// PEs: 16, 20 -> 21
			// srcs: (1776, 31)(3140) 47, (269) -1 --> (3406) -47:PEGB0, ND3, *, PENB
			10'd39 : rdata = 48'b000111110000000001100000011000000000000100000000;
			// PEs: 20, 19 -> 19
			// srcs: (1778, 45)(3) 1, (3405) -47 --> (4189) -47:NM0, PENB, *, PEGB3
			10'd40 : rdata = 48'b000111000000000011011111110000000000000010110000;
			// PEs: 20, 21 -> 20
			// srcs: (1785, 60)(1054) -3, (4190) -47 --> (4974) 44:NW3, PEGB5, -, NW3
			10'd41 : rdata = 48'b000100100000001111100001010000000100110000000000;
			// PEs: 16, 20 -> 
			// srcs: (1804, 32)(3140) 47, (297) 1 --> (3434) 47:PEGB0, ND11, *, 
			10'd42 : rdata = 48'b000111110000000001100001011000000000000000000000;
			// PEs: 20, 20 -> 
			// srcs: (1807, 46)(3) 1, (3434) 47 --> (4218) 47:NM0, ALU, *, 
			10'd43 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 20, 20 -> 20
			// srcs: (1810, 61)(1082) -3, (4218) 47 --> (5002) -50:NW11, ALU, -, NW11
			10'd44 : rdata = 48'b000100100000101100111111111000000110110000000000;
			// PEs: 16, 20 -> 21
			// srcs: (1857, 33)(3140) 47, (350) 2 --> (3487) 94:PEGB0, ND4, *, PENB
			10'd45 : rdata = 48'b000111110000000001100000100000000000000100000000;
			// PEs: 20, 19 -> 19
			// srcs: (1859, 47)(3) 1, (3486) -47 --> (4270) -47:NM0, PENB, *, PEGB3
			10'd46 : rdata = 48'b000111000000000011011111110000000000000010110000;
			// PEs: 20, 21 -> 20
			// srcs: (1866, 62)(1135) 2, (4271) 94 --> (5055) -92:NW4, PEGB5, -, NW4
			10'd47 : rdata = 48'b000100100000010011100001010000000101000000000000;
			// PEs: 16, 20 -> 21
			// srcs: (1938, 34)(3140) 47, (431) -3 --> (3568) -141:PEGB0, ND5, *, PENB
			10'd48 : rdata = 48'b000111110000000001100000101000000000000100000000;
			// PEs: 20, 19 -> 19
			// srcs: (1940, 48)(3) 1, (3567) -94 --> (4351) -94:NM0, PENB, *, PEGB3
			10'd49 : rdata = 48'b000111000000000011011111110000000000000010110000;
			// PEs: 20, 21 -> 20
			// srcs: (1947, 63)(1216) -2, (4352) -141 --> (5136) 139:NW5, PEGB5, -, NW5
			10'd50 : rdata = 48'b000100100000010111100001010000000101010000000000;
			// PEs: 16, 20 -> 
			// srcs: (1988, 35)(3140) 47, (481) -1 --> (3618) -47:PEGB0, ND12, *, 
			10'd51 : rdata = 48'b000111110000000001100001100000000000000000000000;
			// PEs: 20, 20 -> 
			// srcs: (1991, 49)(3) 1, (3618) -47 --> (4402) -47:NM0, ALU, *, 
			10'd52 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 20, 20 -> 20
			// srcs: (1994, 64)(1266) 0, (4402) -47 --> (5186) 47:NW12, ALU, -, NW12
			10'd53 : rdata = 48'b000100100000110000111111111000000111000000000000;
			// PEs: 16, 20 -> 21
			// srcs: (2018, 36)(3140) 47, (511) 0 --> (3648) 0:PEGB0, ND6, *, PENB
			10'd54 : rdata = 48'b000111110000000001100000110000000000000100000000;
			// PEs: 20, 19 -> 19
			// srcs: (2020, 50)(3) 1, (3647) 47 --> (4431) 47:NM0, PENB, *, PEGB3
			10'd55 : rdata = 48'b000111000000000011011111110000000000000010110000;
			// PEs: 20, 21 -> 20
			// srcs: (2027, 65)(1296) 1, (4432) 0 --> (5216) 1:NW6, PEGB5, -, NW6
			10'd56 : rdata = 48'b000100100000011011100001010000000101100000000000;
			// PEs: 16, 20 -> 20
			// srcs: (2100, 37)(3140) 47, (593) 2 --> (3730) 94:PEGB0, ND7, *, NI0
			10'd57 : rdata = 48'b000111110000000001100000111100000000000000000000;
			// PEs: 20, 19 -> 19
			// srcs: (2102, 51)(3) 1, (3729) 0 --> (4513) 0:NM0, PENB, *, PEGB3
			10'd58 : rdata = 48'b000111000000000011011111110000000000000010110000;
			// PEs: 20, 20 -> 
			// srcs: (2103, 52)(3) 1, (3730) 94 --> (4514) 94:NM0, NI0, *, 
			10'd59 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 20, 20 -> 20
			// srcs: (2106, 66)(1378) 2, (4514) 94 --> (5298) -92:NW7, ALU, -, NW7
			10'd60 : rdata = 48'b000100100000011100111111111000000101110000000000;
			// PEs: 16, 20 -> 
			// srcs: (2172, 38)(3140) 47, (665) 0 --> (3802) 0:PEGB0, ND13, *, 
			10'd61 : rdata = 48'b000111110000000001100001101000000000000000000000;
			// PEs: 20, 20 -> 
			// srcs: (2175, 53)(3) 1, (3802) 0 --> (4586) 0:NM0, ALU, *, 
			10'd62 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 20, 20 -> 20
			// srcs: (2178, 67)(1450) 2, (4586) 0 --> (5370) 2:NW13, ALU, -, NW13
			10'd63 : rdata = 48'b000100100000110100111111111000000111010000000000;
			// PEs: 16, 20 -> 
			// srcs: (2180, 39)(3140) 47, (673) 1 --> (3810) 47:PEGB0, ND8, *, 
			10'd64 : rdata = 48'b000111110000000001100001000000000000000000000000;
			// PEs: 20, 20 -> 
			// srcs: (2183, 54)(3) 1, (3810) 47 --> (4594) 47:NM0, ALU, *, 
			10'd65 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 20, 20 -> 20
			// srcs: (2186, 68)(1458) 1, (4594) 47 --> (5378) -46:NW8, ALU, -, NW8
			10'd66 : rdata = 48'b000100100000100000111111111000000110000000000000;
			// PEs: 16, 20 -> 21
			// srcs: (2260, 40)(3140) 47, (753) -2 --> (3890) -94:PEGB0, ND9, *, PENB
			10'd67 : rdata = 48'b000111110000000001100001001000000000000100000000;
			// PEs: 20, 19 -> 19
			// srcs: (2262, 55)(3) 1, (3889) 94 --> (4673) 94:NM0, PENB, *, PEGB3
			10'd68 : rdata = 48'b000111000000000011011111110000000000000010110000;
			// PEs: 20, 21 -> 20
			// srcs: (2269, 69)(1538) -2, (4674) -94 --> (5458) 92:NW9, PEGB5, -, NW9
			10'd69 : rdata = 48'b000100100000100111100001010000000110010000000000;
			default : rdata = 48'b000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 21) begin
	always @(*) begin
		case(address)
			// PEs: 21, 21 -> 16
			// srcs: (1, 0)(29) 2, (814) 2 --> (1598) 4:ND0, NW0, *, PEGB0
			10'd0 : rdata = 48'b000110110000000001000000000000000000000010000000;
			// PEs: 21, 21 -> 16
			// srcs: (2, 1)(109) -1, (894) 1 --> (1678) -1:ND1, NW1, *, PEGB0
			10'd1 : rdata = 48'b000110110000000101000000001000000000000010000000;
			// PEs: 21, 21 -> 16
			// srcs: (3, 2)(191) -2, (976) 2 --> (1760) -4:ND2, NW2, *, PEGB0
			10'd2 : rdata = 48'b000110110000001001000000010000000000000010000000;
			// PEs: 21, 21 -> 16
			// srcs: (4, 3)(271) -1, (1056) 1 --> (1840) -1:ND3, NW3, *, PEGB0
			10'd3 : rdata = 48'b000110110000001101000000011000000000000010000000;
			// PEs: 21, 21 -> 16
			// srcs: (5, 4)(351) -3, (1136) -2 --> (1920) 6:ND4, NW4, *, PEGB0
			10'd4 : rdata = 48'b000110110000010001000000100000000000000010000000;
			// PEs: 21, 21 -> 16
			// srcs: (6, 5)(433) -2, (1218) 2 --> (2002) -4:ND5, NW5, *, PEGB0
			10'd5 : rdata = 48'b000110110000010101000000101000000000000010000000;
			// PEs: 21, 21 -> 16
			// srcs: (7, 6)(513) 2, (1298) 1 --> (2082) 2:ND6, NW6, *, PEGB0
			10'd6 : rdata = 48'b000110110000011001000000110000000000000010000000;
			// PEs: 21, 21 -> 16
			// srcs: (8, 7)(594) -3, (1379) -1 --> (2163) 3:ND7, NW7, *, PEGB0
			10'd7 : rdata = 48'b000110110000011101000000111000000000000010000000;
			// PEs: 21, 21 -> 20
			// srcs: (9, 8)(675) 2, (1460) 2 --> (2244) 4:ND8, NW8, *, PEGB4
			10'd8 : rdata = 48'b000110110000100001000001000000000000000011000000;
			// PEs: 21, 21 -> 23
			// srcs: (10, 9)(755) 2, (1540) 2 --> (2324) 4:ND9, NW9, *, PEGB7
			10'd9 : rdata = 48'b000110110000100101000001001000000000000011110000;
			// PEs: 21, 21 -> 16
			// srcs: (11, 10)(120) -2, (905) 0 --> (1689) 0:ND10, NW10, *, PEGB0
			10'd10 : rdata = 48'b000110110000101001000001010000000000000010000000;
			// PEs: 21, 21 -> 16
			// srcs: (12, 11)(304) 1, (1089) 2 --> (1873) 2:ND11, NW11, *, PEGB0
			10'd11 : rdata = 48'b000110110000101101000001011000000000000010000000;
			// PEs: 21, 21 -> 16
			// srcs: (13, 12)(484) -2, (1269) -2 --> (2053) 4:ND12, NW12, *, PEGB0
			10'd12 : rdata = 48'b000110110000110001000001100000000000000010000000;
			// PEs: 21, 21 -> 21
			// srcs: (14, 13)(668) 1, (1453) -3 --> (2237) -3:ND13, NW13, *, NI0
			10'd13 : rdata = 48'b000110110000110101000001101100000000000000000000;
			// PEs: 18 -> 
			// srcs: (15, 18)(2319) 0 --> (2319) 0:PEGB2, pass, 
			10'd14 : rdata = 48'b110001110000010000000000000000000000000000000000;
			// PEs: 17, 21 -> 16
			// srcs: (18, 19)(2318) 2, (2319) 0 --> (3096) 2:PEGB1, ALU, +, PEGB0
			10'd15 : rdata = 48'b000011110000001000111111111000000000000010000000;
			// PEs: 19 -> 
			// srcs: (20, 21)(3017) -5 --> (3017) -5:PEGB3, pass, 
			10'd16 : rdata = 48'b110001110000011000000000000000000000000000000000;
			// PEs: 21, 22 -> 21
			// srcs: (23, 22)(3017) -5, (2240) 0 --> (3018) -5:ALU, PEGB6, +, NI1
			10'd17 : rdata = 48'b000010011111111111100001100100001000000000000000;
			// PEs: 16 -> 
			// srcs: (25, 14)(1627) 6 --> (1627) 6:PEGB0, pass, 
			10'd18 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 16, 21 -> 17
			// srcs: (34, 15)(1626) 0, (1627) 6 --> (2408) 6:PEGB0, ALU, +, PEGB1
			10'd19 : rdata = 48'b000011110000000000111111111000000000000010010000;
			// PEs: 16 -> 
			// srcs: (71, 16)(1826) -2 --> (1826) -2:PEGB0, pass, 
			10'd20 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 16, 21 -> 17
			// srcs: (80, 17)(1825) 1, (1826) -2 --> (2606) -1:PEGB0, ALU, +, PEGB1
			10'd21 : rdata = 48'b000011110000000000111111111000000000000010010000;
			// PEs: 21 -> 17
			// srcs: (584, 20)(2237) -3 --> (2237) -3:NI0, pass, PEGB1
			10'd22 : rdata = 48'b110001010000000000000000000000000000000010010000;
			// PEs: 17, 21 -> 16
			// srcs: (595, 23)(3016) -6, (3018) -5 --> (3019) -11:PEGB1, NI1, +, PEGB0
			10'd23 : rdata = 48'b000011110000001010100000001000000000000010000000;
			// PEs: 16 -> 
			// srcs: (641, 24)(2764) -4 --> (2764) -4:PEGB0, pass, 
			10'd24 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 21, 17 -> 17
			// srcs: (643, 25)(2764) -4, (2769) 2 --> (2770) -2:ALU, PEGB1, +, PEGB1
			10'd25 : rdata = 48'b000010011111111111100000010000000000000010010000;
			// PEs: 16, 21 -> 22
			// srcs: (1536, 26)(3140) 47, (29) 2 --> (3166) 94:PEGB0, ND0, *, PENB
			10'd26 : rdata = 48'b000111110000000001100000000000000000000100000000;
			// PEs: 21, 20 -> 20
			// srcs: (1537, 40)(3) 1, (3164) -141 --> (3948) -141:NM0, PENB, *, PEGB4
			10'd27 : rdata = 48'b000111000000000011011111110000000000000011000000;
			// PEs: 21, 22 -> 21
			// srcs: (1545, 56)(814) 2, (3950) 94 --> (4734) -92:NW0, PEGB6, -, NW0
			10'd28 : rdata = 48'b000100100000000011100001100000000100000000000000;
			// PEs: 16, 21 -> 22
			// srcs: (1616, 27)(3140) 47, (109) -1 --> (3246) -47:PEGB0, ND1, *, PENB
			10'd29 : rdata = 48'b000111110000000001100000001000000000000100000000;
			// PEs: 21, 20 -> 20
			// srcs: (1617, 41)(3) 1, (3244) 94 --> (4028) 94:NM0, PENB, *, PEGB4
			10'd30 : rdata = 48'b000111000000000011011111110000000000000011000000;
			// PEs: 21, 22 -> 21
			// srcs: (1625, 57)(894) 1, (4030) -47 --> (4814) 48:NW1, PEGB6, -, NW1
			10'd31 : rdata = 48'b000100100000000111100001100000000100010000000000;
			// PEs: 16, 21 -> 
			// srcs: (1627, 28)(3140) 47, (120) -2 --> (3257) -94:PEGB0, ND10, *, 
			10'd32 : rdata = 48'b000111110000000001100001010000000000000000000000;
			// PEs: 21, 21 -> 
			// srcs: (1630, 42)(3) 1, (3257) -94 --> (4041) -94:NM0, ALU, *, 
			10'd33 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 21, 21 -> 21
			// srcs: (1633, 58)(905) 0, (4041) -94 --> (4825) 94:NW10, ALU, -, NW10
			10'd34 : rdata = 48'b000100100000101000111111111000000110100000000000;
			// PEs: 16, 21 -> 22
			// srcs: (1698, 29)(3140) 47, (191) -2 --> (3328) -94:PEGB0, ND2, *, PENB
			10'd35 : rdata = 48'b000111110000000001100000010000000000000100000000;
			// PEs: 21, 20 -> 20
			// srcs: (1699, 43)(3) 1, (3326) 0 --> (4110) 0:NM0, PENB, *, PEGB4
			10'd36 : rdata = 48'b000111000000000011011111110000000000000011000000;
			// PEs: 21, 22 -> 21
			// srcs: (1707, 59)(976) 2, (4112) -94 --> (4896) 96:NW2, PEGB6, -, NW2
			10'd37 : rdata = 48'b000100100000001011100001100000000100100000000000;
			// PEs: 16, 21 -> 21
			// srcs: (1778, 30)(3140) 47, (271) -1 --> (3408) -47:PEGB0, ND3, *, NI0
			10'd38 : rdata = 48'b000111110000000001100000011100000000000000000000;
			// PEs: 21, 20 -> 20
			// srcs: (1779, 44)(3) 1, (3406) -47 --> (4190) -47:NM0, PENB, *, PEGB4
			10'd39 : rdata = 48'b000111000000000011011111110000000000000011000000;
			// PEs: 21, 21 -> 
			// srcs: (1781, 45)(3) 1, (3408) -47 --> (4192) -47:NM0, NI0, *, 
			10'd40 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 21, 21 -> 21
			// srcs: (1784, 60)(1056) 1, (4192) -47 --> (4976) 48:NW3, ALU, -, NW3
			10'd41 : rdata = 48'b000100100000001100111111111000000100110000000000;
			// PEs: 16, 21 -> 
			// srcs: (1811, 31)(3140) 47, (304) 1 --> (3441) 47:PEGB0, ND11, *, 
			10'd42 : rdata = 48'b000111110000000001100001011000000000000000000000;
			// PEs: 21, 21 -> 
			// srcs: (1814, 46)(3) 1, (3441) 47 --> (4225) 47:NM0, ALU, *, 
			10'd43 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 21, 21 -> 21
			// srcs: (1817, 61)(1089) 2, (4225) 47 --> (5009) -45:NW11, ALU, -, NW11
			10'd44 : rdata = 48'b000100100000101100111111111000000110110000000000;
			// PEs: 16, 21 -> 22
			// srcs: (1858, 32)(3140) 47, (351) -3 --> (3488) -141:PEGB0, ND4, *, PENB
			10'd45 : rdata = 48'b000111110000000001100000100000000000000100000000;
			// PEs: 21, 20 -> 20
			// srcs: (1860, 47)(3) 1, (3487) 94 --> (4271) 94:NM0, PENB, *, PEGB4
			10'd46 : rdata = 48'b000111000000000011011111110000000000000011000000;
			// PEs: 21, 22 -> 21
			// srcs: (1867, 62)(1136) -2, (4272) -141 --> (5056) 139:NW4, PEGB6, -, NW4
			10'd47 : rdata = 48'b000100100000010011100001100000000101000000000000;
			// PEs: 16, 21 -> 22
			// srcs: (1940, 33)(3140) 47, (433) -2 --> (3570) -94:PEGB0, ND5, *, PENB
			10'd48 : rdata = 48'b000111110000000001100000101000000000000100000000;
			// PEs: 21, 20 -> 20
			// srcs: (1941, 48)(3) 1, (3568) -141 --> (4352) -141:NM0, PENB, *, PEGB4
			10'd49 : rdata = 48'b000111000000000011011111110000000000000011000000;
			// PEs: 21, 22 -> 21
			// srcs: (1949, 63)(1218) 2, (4354) -94 --> (5138) 96:NW5, PEGB6, -, NW5
			10'd50 : rdata = 48'b000100100000010111100001100000000101010000000000;
			// PEs: 16, 21 -> 
			// srcs: (1991, 34)(3140) 47, (484) -2 --> (3621) -94:PEGB0, ND12, *, 
			10'd51 : rdata = 48'b000111110000000001100001100000000000000000000000;
			// PEs: 21, 21 -> 
			// srcs: (1994, 49)(3) 1, (3621) -94 --> (4405) -94:NM0, ALU, *, 
			10'd52 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 21, 21 -> 21
			// srcs: (1997, 64)(1269) -2, (4405) -94 --> (5189) 92:NW12, ALU, -, NW12
			10'd53 : rdata = 48'b000100100000110000111111111000000111000000000000;
			// PEs: 16, 21 -> 21
			// srcs: (2020, 35)(3140) 47, (513) 2 --> (3650) 94:PEGB0, ND6, *, NI0
			10'd54 : rdata = 48'b000111110000000001100000110100000000000000000000;
			// PEs: 21, 20 -> 20
			// srcs: (2021, 50)(3) 1, (3648) 0 --> (4432) 0:NM0, PENB, *, PEGB4
			10'd55 : rdata = 48'b000111000000000011011111110000000000000011000000;
			// PEs: 21, 21 -> 
			// srcs: (2023, 51)(3) 1, (3650) 94 --> (4434) 94:NM0, NI0, *, 
			10'd56 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 21, 21 -> 21
			// srcs: (2026, 65)(1298) 1, (4434) 94 --> (5218) -93:NW6, ALU, -, NW6
			10'd57 : rdata = 48'b000100100000011000111111111000000101100000000000;
			// PEs: 16, 21 -> 
			// srcs: (2101, 36)(3140) 47, (594) -3 --> (3731) -141:PEGB0, ND7, *, 
			10'd58 : rdata = 48'b000111110000000001100000111000000000000000000000;
			// PEs: 21, 21 -> 
			// srcs: (2104, 52)(3) 1, (3731) -141 --> (4515) -141:NM0, ALU, *, 
			10'd59 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 21, 21 -> 21
			// srcs: (2107, 66)(1379) -1, (4515) -141 --> (5299) 140:NW7, ALU, -, NW7
			10'd60 : rdata = 48'b000100100000011100111111111000000101110000000000;
			// PEs: 16, 21 -> 
			// srcs: (2175, 37)(3140) 47, (668) 1 --> (3805) 47:PEGB0, ND13, *, 
			10'd61 : rdata = 48'b000111110000000001100001101000000000000000000000;
			// PEs: 21, 21 -> 
			// srcs: (2178, 53)(3) 1, (3805) 47 --> (4589) 47:NM0, ALU, *, 
			10'd62 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 21, 21 -> 21
			// srcs: (2181, 67)(1453) -3, (4589) 47 --> (5373) -50:NW13, ALU, -, NW13
			10'd63 : rdata = 48'b000100100000110100111111111000000111010000000000;
			// PEs: 16, 21 -> 
			// srcs: (2182, 38)(3140) 47, (675) 2 --> (3812) 94:PEGB0, ND8, *, 
			10'd64 : rdata = 48'b000111110000000001100001000000000000000000000000;
			// PEs: 21, 21 -> 
			// srcs: (2185, 54)(3) 1, (3812) 94 --> (4596) 94:NM0, ALU, *, 
			10'd65 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 21, 21 -> 21
			// srcs: (2188, 68)(1460) 2, (4596) 94 --> (5380) -92:NW8, ALU, -, NW8
			10'd66 : rdata = 48'b000100100000100000111111111000000110000000000000;
			// PEs: 16, 21 -> 22
			// srcs: (2262, 39)(3140) 47, (755) 2 --> (3892) 94:PEGB0, ND9, *, PENB
			10'd67 : rdata = 48'b000111110000000001100001001000000000000100000000;
			// PEs: 21, 20 -> 20
			// srcs: (2263, 55)(3) 1, (3890) -94 --> (4674) -94:NM0, PENB, *, PEGB4
			10'd68 : rdata = 48'b000111000000000011011111110000000000000011000000;
			// PEs: 21, 22 -> 21
			// srcs: (2271, 69)(1540) 2, (4676) 94 --> (5460) -92:NW9, PEGB6, -, NW9
			10'd69 : rdata = 48'b000100100000100111100001100000000110010000000000;
			default : rdata = 48'b000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 22) begin
	always @(*) begin
		case(address)
			// PEs: 22, 22 -> 16
			// srcs: (1, 0)(30) 1, (815) -2 --> (1599) -2:ND0, NW0, *, PEGB0
			10'd0 : rdata = 48'b000110110000000001000000000000000000000010000000;
			// PEs: 22, 22 -> 16
			// srcs: (2, 1)(110) 2, (895) -2 --> (1679) -4:ND1, NW1, *, PEGB0
			10'd1 : rdata = 48'b000110110000000101000000001000000000000010000000;
			// PEs: 22, 22 -> 16
			// srcs: (3, 2)(192) 1, (977) -1 --> (1761) -1:ND2, NW2, *, PEGB0
			10'd2 : rdata = 48'b000110110000001001000000010000000000000010000000;
			// PEs: 22, 22 -> 16
			// srcs: (4, 3)(272) 1, (1057) -1 --> (1841) -1:ND3, NW3, *, PEGB0
			10'd3 : rdata = 48'b000110110000001101000000011000000000000010000000;
			// PEs: 22, 22 -> 16
			// srcs: (5, 4)(352) -3, (1137) 2 --> (1921) -6:ND4, NW4, *, PEGB0
			10'd4 : rdata = 48'b000110110000010001000000100000000000000010000000;
			// PEs: 22, 22 -> 16
			// srcs: (6, 5)(434) 2, (1219) 1 --> (2003) 2:ND5, NW5, *, PEGB0
			10'd5 : rdata = 48'b000110110000010101000000101000000000000010000000;
			// PEs: 22, 22 -> 16
			// srcs: (7, 6)(514) 2, (1299) 0 --> (2083) 0:ND6, NW6, *, PEGB0
			10'd6 : rdata = 48'b000110110000011001000000110000000000000010000000;
			// PEs: 22, 22 -> 16
			// srcs: (8, 7)(595) 2, (1380) 2 --> (2164) 4:ND7, NW7, *, PEGB0
			10'd7 : rdata = 48'b000110110000011101000000111000000000000010000000;
			// PEs: 22, 22 -> 20
			// srcs: (9, 8)(676) -3, (1461) 2 --> (2245) -6:ND8, NW8, *, PEGB4
			10'd8 : rdata = 48'b000110110000100001000001000000000000000011000000;
			// PEs: 22, 22 -> 23
			// srcs: (10, 9)(756) 2, (1541) -2 --> (2325) -4:ND9, NW9, *, PENB
			10'd9 : rdata = 48'b000110110000100101000001001000000000000100000000;
			// PEs: 22, 22 -> 22
			// srcs: (11, 10)(123) 0, (908) 2 --> (1692) 0:ND10, NW10, *, NI0
			10'd10 : rdata = 48'b000110110000101001000001010100000000000000000000;
			// PEs: 22, 22 -> 17
			// srcs: (12, 11)(307) 2, (1092) -1 --> (1876) -2:ND11, NW11, *, PEGB1
			10'd11 : rdata = 48'b000110110000101101000001011000000000000010010000;
			// PEs: 22, 22 -> 22
			// srcs: (13, 12)(487) 0, (1272) 2 --> (2056) 0:ND12, NW12, *, NI1
			10'd12 : rdata = 48'b000110110000110001000001100100001000000000000000;
			// PEs: 22, 22 -> 21
			// srcs: (14, 13)(671) 0, (1456) -2 --> (2240) 0:ND13, NW13, *, PEGB5
			10'd13 : rdata = 48'b000110110000110101000001101000000000000011010000;
			// PEs: 20 -> 
			// srcs: (15, 18)(2322) 4 --> (2322) 4:PEGB4, pass, 
			10'd14 : rdata = 48'b110001110000100000000000000000000000000000000000;
			// PEs: 19, 22 -> 22
			// srcs: (18, 19)(2321) -2, (2322) 4 --> (3100) 2:PEGB3, ALU, +, NI2
			10'd15 : rdata = 48'b000011110000011000111111111100010000000000000000;
			// PEs: 18 -> 
			// srcs: (23, 22)(3020) 1 --> (3020) 1:PEGB2, pass, 
			10'd16 : rdata = 48'b110001110000010000000000000000000000000000000000;
			// PEs: 22, 23 -> 22
			// srcs: (26, 23)(3020) 1, (2243) -2 --> (3021) -1:ALU, PEGB7, +, NI3
			10'd17 : rdata = 48'b000010011111111111100001110100011000000000000000;
			// PEs: 16 -> 
			// srcs: (28, 14)(1630) -2 --> (1630) -2:PEGB0, pass, 
			10'd18 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 16, 22 -> 16
			// srcs: (37, 15)(1629) 2, (1630) -2 --> (2411) 0:PEGB0, ALU, +, PEGB0
			10'd19 : rdata = 48'b000011110000000000111111111000000000000010000000;
			// PEs: 16 -> 
			// srcs: (73, 16)(1829) 0 --> (1829) 0:PEGB0, pass, 
			10'd20 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 16, 22 -> 16
			// srcs: (82, 17)(1828) 0, (1829) 0 --> (2608) 0:PEGB0, ALU, +, PEGB0
			10'd21 : rdata = 48'b000011110000000000111111111000000000000010000000;
			// PEs: 22 -> 16
			// srcs: (185, 20)(1692) 0 --> (1692) 0:NI0, pass, PEGB0
			10'd22 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 22 -> 16
			// srcs: (205, 24)(3100) 2 --> (3100) 2:NI2, pass, PEGB0
			10'd23 : rdata = 48'b110001010000001000000000000000000000000010000000;
			// PEs: 22 -> 16
			// srcs: (226, 21)(2056) 0 --> (2056) 0:NI1, pass, PEGB0
			10'd24 : rdata = 48'b110001010000000100000000000000000000000010000000;
			// PEs: 22 -> 16
			// srcs: (398, 25)(3021) -1 --> (3021) -1:NI3, pass, PEGB0
			10'd25 : rdata = 48'b110001010000001100000000000000000000000010000000;
			// PEs: 16, 22 -> 23
			// srcs: (1537, 26)(3140) 47, (30) 1 --> (3167) 47:PEGB0, ND0, *, PENB
			10'd26 : rdata = 48'b000111110000000001100000000000000000000100000000;
			// PEs: 22, 21 -> 21
			// srcs: (1539, 40)(3) 1, (3166) 94 --> (3950) 94:NM0, PENB, *, PEGB5
			10'd27 : rdata = 48'b000111000000000011011111110000000000000011010000;
			// PEs: 22, 23 -> 22
			// srcs: (1546, 56)(815) -2, (3951) 47 --> (4735) -49:NW0, PEGB7, -, NW0
			10'd28 : rdata = 48'b000100100000000011100001110000000100000000000000;
			// PEs: 16, 22 -> 23
			// srcs: (1617, 27)(3140) 47, (110) 2 --> (3247) 94:PEGB0, ND1, *, PENB
			10'd29 : rdata = 48'b000111110000000001100000001000000000000100000000;
			// PEs: 22, 21 -> 21
			// srcs: (1619, 41)(3) 1, (3246) -47 --> (4030) -47:NM0, PENB, *, PEGB5
			10'd30 : rdata = 48'b000111000000000011011111110000000000000011010000;
			// PEs: 22, 23 -> 22
			// srcs: (1626, 57)(895) -2, (4031) 94 --> (4815) -96:NW1, PEGB7, -, NW1
			10'd31 : rdata = 48'b000100100000000111100001110000000100010000000000;
			// PEs: 16, 22 -> 
			// srcs: (1630, 28)(3140) 47, (123) 0 --> (3260) 0:PEGB0, ND10, *, 
			10'd32 : rdata = 48'b000111110000000001100001010000000000000000000000;
			// PEs: 22, 22 -> 
			// srcs: (1633, 42)(3) 1, (3260) 0 --> (4044) 0:NM0, ALU, *, 
			10'd33 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 22, 22 -> 22
			// srcs: (1636, 58)(908) 2, (4044) 0 --> (4828) 2:NW10, ALU, -, NW10
			10'd34 : rdata = 48'b000100100000101000111111111000000110100000000000;
			// PEs: 16, 22 -> 22
			// srcs: (1699, 29)(3140) 47, (192) 1 --> (3329) 47:PEGB0, ND2, *, NI0
			10'd35 : rdata = 48'b000111110000000001100000010100000000000000000000;
			// PEs: 22, 21 -> 21
			// srcs: (1701, 43)(3) 1, (3328) -94 --> (4112) -94:NM0, PENB, *, PEGB5
			10'd36 : rdata = 48'b000111000000000011011111110000000000000011010000;
			// PEs: 22, 22 -> 
			// srcs: (1702, 44)(3) 1, (3329) 47 --> (4113) 47:NM0, NI0, *, 
			10'd37 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 22, 22 -> 22
			// srcs: (1705, 59)(977) -1, (4113) 47 --> (4897) -48:NW2, ALU, -, NW2
			10'd38 : rdata = 48'b000100100000001000111111111000000100100000000000;
			// PEs: 16, 22 -> 
			// srcs: (1779, 30)(3140) 47, (272) 1 --> (3409) 47:PEGB0, ND3, *, 
			10'd39 : rdata = 48'b000111110000000001100000011000000000000000000000;
			// PEs: 22, 22 -> 
			// srcs: (1782, 45)(3) 1, (3409) 47 --> (4193) 47:NM0, ALU, *, 
			10'd40 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 22, 22 -> 22
			// srcs: (1785, 60)(1057) -1, (4193) 47 --> (4977) -48:NW3, ALU, -, NW3
			10'd41 : rdata = 48'b000100100000001100111111111000000100110000000000;
			// PEs: 16, 22 -> 
			// srcs: (1814, 31)(3140) 47, (307) 2 --> (3444) 94:PEGB0, ND11, *, 
			10'd42 : rdata = 48'b000111110000000001100001011000000000000000000000;
			// PEs: 22, 22 -> 
			// srcs: (1817, 46)(3) 1, (3444) 94 --> (4228) 94:NM0, ALU, *, 
			10'd43 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 22, 22 -> 22
			// srcs: (1820, 61)(1092) -1, (4228) 94 --> (5012) -95:NW11, ALU, -, NW11
			10'd44 : rdata = 48'b000100100000101100111111111000000110110000000000;
			// PEs: 16, 22 -> 23
			// srcs: (1859, 32)(3140) 47, (352) -3 --> (3489) -141:PEGB0, ND4, *, PENB
			10'd45 : rdata = 48'b000111110000000001100000100000000000000100000000;
			// PEs: 22, 21 -> 21
			// srcs: (1861, 47)(3) 1, (3488) -141 --> (4272) -141:NM0, PENB, *, PEGB5
			10'd46 : rdata = 48'b000111000000000011011111110000000000000011010000;
			// PEs: 22, 23 -> 22
			// srcs: (1868, 62)(1137) 2, (4273) -141 --> (5057) 143:NW4, PEGB7, -, NW4
			10'd47 : rdata = 48'b000100100000010011100001110000000101000000000000;
			// PEs: 16, 22 -> 22
			// srcs: (1941, 33)(3140) 47, (434) 2 --> (3571) 94:PEGB0, ND5, *, NI0
			10'd48 : rdata = 48'b000111110000000001100000101100000000000000000000;
			// PEs: 22, 21 -> 21
			// srcs: (1943, 48)(3) 1, (3570) -94 --> (4354) -94:NM0, PENB, *, PEGB5
			10'd49 : rdata = 48'b000111000000000011011111110000000000000011010000;
			// PEs: 22, 22 -> 
			// srcs: (1944, 49)(3) 1, (3571) 94 --> (4355) 94:NM0, NI0, *, 
			10'd50 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 22, 22 -> 22
			// srcs: (1947, 63)(1219) 1, (4355) 94 --> (5139) -93:NW5, ALU, -, NW5
			10'd51 : rdata = 48'b000100100000010100111111111000000101010000000000;
			// PEs: 16, 22 -> 
			// srcs: (1994, 34)(3140) 47, (487) 0 --> (3624) 0:PEGB0, ND12, *, 
			10'd52 : rdata = 48'b000111110000000001100001100000000000000000000000;
			// PEs: 22, 22 -> 
			// srcs: (1997, 50)(3) 1, (3624) 0 --> (4408) 0:NM0, ALU, *, 
			10'd53 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 22, 22 -> 22
			// srcs: (2000, 64)(1272) 2, (4408) 0 --> (5192) 2:NW12, ALU, -, NW12
			10'd54 : rdata = 48'b000100100000110000111111111000000111000000000000;
			// PEs: 16, 22 -> 
			// srcs: (2021, 35)(3140) 47, (514) 2 --> (3651) 94:PEGB0, ND6, *, 
			10'd55 : rdata = 48'b000111110000000001100000110000000000000000000000;
			// PEs: 22, 22 -> 
			// srcs: (2024, 51)(3) 1, (3651) 94 --> (4435) 94:NM0, ALU, *, 
			10'd56 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 22, 22 -> 22
			// srcs: (2027, 65)(1299) 0, (4435) 94 --> (5219) -94:NW6, ALU, -, NW6
			10'd57 : rdata = 48'b000100100000011000111111111000000101100000000000;
			// PEs: 16, 22 -> 
			// srcs: (2102, 36)(3140) 47, (595) 2 --> (3732) 94:PEGB0, ND7, *, 
			10'd58 : rdata = 48'b000111110000000001100000111000000000000000000000;
			// PEs: 22, 22 -> 
			// srcs: (2105, 52)(3) 1, (3732) 94 --> (4516) 94:NM0, ALU, *, 
			10'd59 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 22, 22 -> 22
			// srcs: (2108, 66)(1380) 2, (4516) 94 --> (5300) -92:NW7, ALU, -, NW7
			10'd60 : rdata = 48'b000100100000011100111111111000000101110000000000;
			// PEs: 16, 22 -> 
			// srcs: (2178, 37)(3140) 47, (671) 0 --> (3808) 0:PEGB0, ND13, *, 
			10'd61 : rdata = 48'b000111110000000001100001101000000000000000000000;
			// PEs: 22, 22 -> 22
			// srcs: (2181, 53)(3) 1, (3808) 0 --> (4592) 0:NM0, ALU, *, NI0
			10'd62 : rdata = 48'b000111000000000000111111111100000000000000000000;
			// PEs: 16, 22 -> 22
			// srcs: (2183, 38)(3140) 47, (676) -3 --> (3813) -141:PEGB0, ND8, *, NI1
			10'd63 : rdata = 48'b000111110000000001100001000100001000000000000000;
			// PEs: 22, 22 -> 22
			// srcs: (2184, 67)(1456) -2, (4592) 0 --> (5376) -2:NW13, NI0, -, NW13
			10'd64 : rdata = 48'b000100100000110110100000000000000111010000000000;
			// PEs: 22, 22 -> 
			// srcs: (2186, 54)(3) 1, (3813) -141 --> (4597) -141:NM0, NI1, *, 
			10'd65 : rdata = 48'b000111000000000010100000001000000000000000000000;
			// PEs: 22, 22 -> 22
			// srcs: (2189, 68)(1461) 2, (4597) -141 --> (5381) 143:NW8, ALU, -, NW8
			10'd66 : rdata = 48'b000100100000100000111111111000000110000000000000;
			// PEs: 16, 22 -> 23
			// srcs: (2263, 39)(3140) 47, (756) 2 --> (3893) 94:PEGB0, ND9, *, PENB
			10'd67 : rdata = 48'b000111110000000001100001001000000000000100000000;
			// PEs: 22, 21 -> 21
			// srcs: (2265, 55)(3) 1, (3892) 94 --> (4676) 94:NM0, PENB, *, PEGB5
			10'd68 : rdata = 48'b000111000000000011011111110000000000000011010000;
			// PEs: 22, 23 -> 22
			// srcs: (2272, 69)(1541) -2, (4677) 94 --> (5461) -96:NW9, PEGB7, -, NW9
			10'd69 : rdata = 48'b000100100000100111100001110000000110010000000000;
			default : rdata = 48'b000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 23) begin
	always @(*) begin
		case(address)
			// PEs: 23, 23 -> 16
			// srcs: (1, 0)(32) -2, (817) -2 --> (1601) 4:ND0, NW0, *, PENB
			10'd0 : rdata = 48'b000110110000000001000000000000000000000100000000;
			// PEs: 23, 23 -> 16
			// srcs: (2, 1)(112) -1, (897) -3 --> (1681) 3:ND1, NW1, *, PENB
			10'd1 : rdata = 48'b000110110000000101000000001000000000000100000000;
			// PEs: 23, 23 -> 16
			// srcs: (3, 2)(194) 0, (979) -2 --> (1763) 0:ND2, NW2, *, PENB
			10'd2 : rdata = 48'b000110110000001001000000010000000000000100000000;
			// PEs: 23, 23 -> 16
			// srcs: (4, 3)(274) 1, (1059) 1 --> (1843) 1:ND3, NW3, *, PENB
			10'd3 : rdata = 48'b000110110000001101000000011000000000000100000000;
			// PEs: 23, 23 -> 16
			// srcs: (5, 4)(354) -3, (1139) 2 --> (1923) -6:ND4, NW4, *, PENB
			10'd4 : rdata = 48'b000110110000010001000000100000000000000100000000;
			// PEs: 23, 23 -> 16
			// srcs: (6, 5)(436) -1, (1221) -1 --> (2005) 1:ND5, NW5, *, PENB
			10'd5 : rdata = 48'b000110110000010101000000101000000000000100000000;
			// PEs: 23, 23 -> 16
			// srcs: (7, 6)(516) 0, (1301) -3 --> (2085) 0:ND6, NW6, *, PENB
			10'd6 : rdata = 48'b000110110000011001000000110000000000000100000000;
			// PEs: 23, 23 -> 16
			// srcs: (8, 7)(596) -1, (1381) 0 --> (2165) 0:ND7, NW7, *, PENB
			10'd7 : rdata = 48'b000110110000011101000000111000000000000100000000;
			// PEs: 23, 23 -> 16
			// srcs: (9, 8)(678) 1, (1463) -2 --> (2247) -2:ND8, NW8, *, PENB
			10'd8 : rdata = 48'b000110110000100001000001000000000000000100000000;
			// PEs: 23, 23 -> 16
			// srcs: (10, 9)(758) -3, (1543) 0 --> (2327) 0:ND9, NW9, *, PENB
			10'd9 : rdata = 48'b000110110000100101000001001000000000000100000000;
			// PEs: 23, 23 -> 23
			// srcs: (11, 10)(126) -1, (911) -3 --> (1695) 3:ND10, NW10, *, NI0
			10'd10 : rdata = 48'b000110110000101001000001010100000000000000000000;
			// PEs: 23, 23 -> 23
			// srcs: (12, 11)(310) 2, (1095) 2 --> (1879) 4:ND11, NW11, *, NI1
			10'd11 : rdata = 48'b000110110000101101000001011100001000000000000000;
			// PEs: 23, 23 -> 17
			// srcs: (13, 12)(490) 0, (1275) -2 --> (2059) 0:ND12, NW12, *, PEGB1
			10'd12 : rdata = 48'b000110110000110001000001100000000000000010010000;
			// PEs: 23, 23 -> 22
			// srcs: (14, 13)(674) -1, (1459) 2 --> (2243) -2:ND13, NW13, *, PEGB6
			10'd13 : rdata = 48'b000110110000110101000001101000000000000011100000;
			// PEs: 21, 22 -> 23
			// srcs: (16, 18)(2324) 4, (2325) -4 --> (3102) 0:PEGB5, PENB, +, NI2
			10'd14 : rdata = 48'b000011110000101011011111110100010000000000000000;
			// PEs: 16 -> 
			// srcs: (31, 14)(1633) -6 --> (1633) -6:PEGB0, pass, 
			10'd15 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 16, 23 -> 16
			// srcs: (40, 15)(1632) 0, (1633) -6 --> (2413) -6:PEGB0, ALU, +, PENB
			10'd16 : rdata = 48'b000011110000000000111111111000000000000100000000;
			// PEs: 16 -> 
			// srcs: (75, 16)(1832) 9 --> (1832) 9:PEGB0, pass, 
			10'd17 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 16, 23 -> 23
			// srcs: (84, 17)(1831) -3, (1832) 9 --> (2612) 6:PEGB0, ALU, +, NI3
			10'd18 : rdata = 48'b000011110000000000111111111100011000000000000000;
			// PEs: 23 -> 16
			// srcs: (120, 21)(1695) 3 --> (1695) 3:NI0, pass, PENB
			10'd19 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 23 -> 16
			// srcs: (141, 23)(1879) 4 --> (1879) 4:NI1, pass, PENB
			10'd20 : rdata = 48'b110001010000000100000000000000000000000100000000;
			// PEs: 23 -> 16
			// srcs: (242, 24)(3102) 0 --> (3102) 0:NI2, pass, PENB
			10'd21 : rdata = 48'b110001010000001000000000000000000000000100000000;
			// PEs: 16 -> 
			// srcs: (250, 19)(1672) 1 --> (1672) 1:PEGB0, pass, 
			10'd22 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 16, 23 -> 16
			// srcs: (259, 20)(1671) 2, (1672) 1 --> (2454) 3:PEGB0, ALU, +, PENB
			10'd23 : rdata = 48'b000011110000000000111111111000000000000100000000;
			// PEs: 23 -> 16
			// srcs: (272, 22)(2612) 6 --> (2612) 6:NI3, pass, PENB
			10'd24 : rdata = 48'b110001010000001100000000000000000000000100000000;
			// PEs: 16, 23 -> 23
			// srcs: (1539, 25)(3140) 47, (32) -2 --> (3169) -94:PEGB0, ND0, *, NI0
			10'd25 : rdata = 48'b000111110000000001100000000100000000000000000000;
			// PEs: 23, 22 -> 22
			// srcs: (1540, 39)(3) 1, (3167) 47 --> (3951) 47:NM0, PENB, *, PEGB6
			10'd26 : rdata = 48'b000111000000000011011111110000000000000011100000;
			// PEs: 23, 23 -> 
			// srcs: (1542, 40)(3) 1, (3169) -94 --> (3953) -94:NM0, NI0, *, 
			10'd27 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 23, 23 -> 23
			// srcs: (1545, 57)(817) -2, (3953) -94 --> (4737) 92:NW0, ALU, -, NW0
			10'd28 : rdata = 48'b000100100000000000111111111000000100000000000000;
			// PEs: 16, 23 -> 23
			// srcs: (1619, 26)(3140) 47, (112) -1 --> (3249) -47:PEGB0, ND1, *, NI0
			10'd29 : rdata = 48'b000111110000000001100000001100000000000000000000;
			// PEs: 23, 22 -> 22
			// srcs: (1620, 41)(3) 1, (3247) 94 --> (4031) 94:NM0, PENB, *, PEGB6
			10'd30 : rdata = 48'b000111000000000011011111110000000000000011100000;
			// PEs: 23, 23 -> 
			// srcs: (1622, 42)(3) 1, (3249) -47 --> (4033) -47:NM0, NI0, *, 
			10'd31 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 23, 23 -> 23
			// srcs: (1625, 58)(897) -3, (4033) -47 --> (4817) 44:NW1, ALU, -, NW1
			10'd32 : rdata = 48'b000100100000000100111111111000000100010000000000;
			// PEs: 16, 23 -> 
			// srcs: (1633, 27)(3140) 47, (126) -1 --> (3263) -47:PEGB0, ND10, *, 
			10'd33 : rdata = 48'b000111110000000001100001010000000000000000000000;
			// PEs: 23, 23 -> 
			// srcs: (1636, 43)(3) 1, (3263) -47 --> (4047) -47:NM0, ALU, *, 
			10'd34 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 23, 23 -> 23
			// srcs: (1639, 59)(911) -3, (4047) -47 --> (4831) 44:NW10, ALU, -, NW10
			10'd35 : rdata = 48'b000100100000101000111111111000000110100000000000;
			// PEs: 16, 23 -> 
			// srcs: (1701, 28)(3140) 47, (194) 0 --> (3331) 0:PEGB0, ND2, *, 
			10'd36 : rdata = 48'b000111110000000001100000010000000000000000000000;
			// PEs: 23, 23 -> 
			// srcs: (1704, 44)(3) 1, (3331) 0 --> (4115) 0:NM0, ALU, *, 
			10'd37 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 23, 23 -> 23
			// srcs: (1707, 60)(979) -2, (4115) 0 --> (4899) -2:NW2, ALU, -, NW2
			10'd38 : rdata = 48'b000100100000001000111111111000000100100000000000;
			// PEs: 16, 23 -> 
			// srcs: (1781, 29)(3140) 47, (274) 1 --> (3411) 47:PEGB0, ND3, *, 
			10'd39 : rdata = 48'b000111110000000001100000011000000000000000000000;
			// PEs: 23, 23 -> 
			// srcs: (1784, 45)(3) 1, (3411) 47 --> (4195) 47:NM0, ALU, *, 
			10'd40 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 23, 23 -> 23
			// srcs: (1787, 61)(1059) 1, (4195) 47 --> (4979) -46:NW3, ALU, -, NW3
			10'd41 : rdata = 48'b000100100000001100111111111000000100110000000000;
			// PEs: 16, 23 -> 
			// srcs: (1817, 30)(3140) 47, (310) 2 --> (3447) 94:PEGB0, ND11, *, 
			10'd42 : rdata = 48'b000111110000000001100001011000000000000000000000;
			// PEs: 23, 23 -> 
			// srcs: (1820, 46)(3) 1, (3447) 94 --> (4231) 94:NM0, ALU, *, 
			10'd43 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 23, 23 -> 23
			// srcs: (1823, 62)(1095) 2, (4231) 94 --> (5015) -92:NW11, ALU, -, NW11
			10'd44 : rdata = 48'b000100100000101100111111111000000110110000000000;
			// PEs: 16, 23 -> 23
			// srcs: (1861, 31)(3140) 47, (354) -3 --> (3491) -141:PEGB0, ND4, *, NI0
			10'd45 : rdata = 48'b000111110000000001100000100100000000000000000000;
			// PEs: 23, 22 -> 22
			// srcs: (1862, 47)(3) 1, (3489) -141 --> (4273) -141:NM0, PENB, *, PEGB6
			10'd46 : rdata = 48'b000111000000000011011111110000000000000011100000;
			// PEs: 23, 23 -> 
			// srcs: (1864, 48)(3) 1, (3491) -141 --> (4275) -141:NM0, NI0, *, 
			10'd47 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 23, 23 -> 23
			// srcs: (1867, 63)(1139) 2, (4275) -141 --> (5059) 143:NW4, ALU, -, NW4
			10'd48 : rdata = 48'b000100100000010000111111111000000101000000000000;
			// PEs: 16, 23 -> 
			// srcs: (1943, 32)(3140) 47, (436) -1 --> (3573) -47:PEGB0, ND5, *, 
			10'd49 : rdata = 48'b000111110000000001100000101000000000000000000000;
			// PEs: 23, 23 -> 
			// srcs: (1946, 49)(3) 1, (3573) -47 --> (4357) -47:NM0, ALU, *, 
			10'd50 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 23, 23 -> 23
			// srcs: (1949, 64)(1221) -1, (4357) -47 --> (5141) 46:NW5, ALU, -, NW5
			10'd51 : rdata = 48'b000100100000010100111111111000000101010000000000;
			// PEs: 16, 23 -> 
			// srcs: (1997, 33)(3140) 47, (490) 0 --> (3627) 0:PEGB0, ND12, *, 
			10'd52 : rdata = 48'b000111110000000001100001100000000000000000000000;
			// PEs: 23, 23 -> 
			// srcs: (2000, 50)(3) 1, (3627) 0 --> (4411) 0:NM0, ALU, *, 
			10'd53 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 23, 23 -> 23
			// srcs: (2003, 65)(1275) -2, (4411) 0 --> (5195) -2:NW12, ALU, -, NW12
			10'd54 : rdata = 48'b000100100000110000111111111000000111000000000000;
			// PEs: 16, 23 -> 
			// srcs: (2023, 34)(3140) 47, (516) 0 --> (3653) 0:PEGB0, ND6, *, 
			10'd55 : rdata = 48'b000111110000000001100000110000000000000000000000;
			// PEs: 23, 23 -> 
			// srcs: (2026, 51)(3) 1, (3653) 0 --> (4437) 0:NM0, ALU, *, 
			10'd56 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 23, 23 -> 23
			// srcs: (2029, 66)(1301) -3, (4437) 0 --> (5221) -3:NW6, ALU, -, NW6
			10'd57 : rdata = 48'b000100100000011000111111111000000101100000000000;
			// PEs: 16, 23 -> 
			// srcs: (2103, 35)(3140) 47, (596) -1 --> (3733) -47:PEGB0, ND7, *, 
			10'd58 : rdata = 48'b000111110000000001100000111000000000000000000000;
			// PEs: 23, 23 -> 
			// srcs: (2106, 52)(3) 1, (3733) -47 --> (4517) -47:NM0, ALU, *, 
			10'd59 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 23, 23 -> 23
			// srcs: (2109, 67)(1381) 0, (4517) -47 --> (5301) 47:NW7, ALU, -, NW7
			10'd60 : rdata = 48'b000100100000011100111111111000000101110000000000;
			// PEs: 16, 23 -> 
			// srcs: (2181, 36)(3140) 47, (674) -1 --> (3811) -47:PEGB0, ND13, *, 
			10'd61 : rdata = 48'b000111110000000001100001101000000000000000000000;
			// PEs: 23, 23 -> 23
			// srcs: (2184, 53)(3) 1, (3811) -47 --> (4595) -47:NM0, ALU, *, NI0
			10'd62 : rdata = 48'b000111000000000000111111111100000000000000000000;
			// PEs: 16, 23 -> 23
			// srcs: (2185, 37)(3140) 47, (678) 1 --> (3815) 47:PEGB0, ND8, *, NI1
			10'd63 : rdata = 48'b000111110000000001100001000100001000000000000000;
			// PEs: 23, 23 -> 23
			// srcs: (2187, 68)(1459) 2, (4595) -47 --> (5379) 49:NW13, NI0, -, NW13
			10'd64 : rdata = 48'b000100100000110110100000000000000111010000000000;
			// PEs: 23, 23 -> 
			// srcs: (2188, 54)(3) 1, (3815) 47 --> (4599) 47:NM0, NI1, *, 
			10'd65 : rdata = 48'b000111000000000010100000001000000000000000000000;
			// PEs: 23, 23 -> 23
			// srcs: (2191, 69)(1463) -2, (4599) 47 --> (5383) -49:NW8, ALU, -, NW8
			10'd66 : rdata = 48'b000100100000100000111111111000000110000000000000;
			// PEs: 16, 23 -> 23
			// srcs: (2265, 38)(3140) 47, (758) -3 --> (3895) -141:PEGB0, ND9, *, NI0
			10'd67 : rdata = 48'b000111110000000001100001001100000000000000000000;
			// PEs: 23, 22 -> 22
			// srcs: (2266, 55)(3) 1, (3893) 94 --> (4677) 94:NM0, PENB, *, PEGB6
			10'd68 : rdata = 48'b000111000000000011011111110000000000000011100000;
			// PEs: 23, 23 -> 
			// srcs: (2268, 56)(3) 1, (3895) -141 --> (4679) -141:NM0, NI0, *, 
			10'd69 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 23, 23 -> 23
			// srcs: (2271, 70)(1543) 0, (4679) -141 --> (5463) 141:NW9, ALU, -, NW9
			10'd70 : rdata = 48'b000100100000100100111111111000000110010000000000;
			default : rdata = 48'b000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 24) begin
	always @(*) begin
		case(address)
			// PEs: 25 -> 8
			// srcs: (6, 0)(1602) -4 --> (1602) -4:PEGB1, pass, PUGB1
			10'd0 : rdata = 48'b110001110000001000000000000000000000000000001001;
			// PEs: 26 -> 8
			// srcs: (7, 1)(1604) -1 --> (1604) -1:PEGB2, pass, PUGB1
			10'd1 : rdata = 48'b110001110000010000000000000000000000000000001001;
			// PEs: 27 -> 8
			// srcs: (8, 2)(1605) -2 --> (1605) -2:PEGB3, pass, PUGB1
			10'd2 : rdata = 48'b110001110000011000000000000000000000000000001001;
			// PEs: 28 -> 8
			// srcs: (9, 3)(1607) -2 --> (1607) -2:PEGB4, pass, PUGB1
			10'd3 : rdata = 48'b110001110000100000000000000000000000000000001001;
			// PEs: 29 -> 8
			// srcs: (10, 4)(1608) 0 --> (1608) 0:PEGB5, pass, PUGB1
			10'd4 : rdata = 48'b110001110000101000000000000000000000000000001001;
			// PEs: 30 -> 8
			// srcs: (11, 5)(1610) -6 --> (1610) -6:PEGB6, pass, PUGB1
			10'd5 : rdata = 48'b110001110000110000000000000000000000000000001001;
			// PEs: 31 -> 8
			// srcs: (12, 6)(1611) -2 --> (1611) -2:PENB, pass, PUGB1
			10'd6 : rdata = 48'b110001101111111000000000000000000000000000001001;
			// PEs: 48 -> 24
			// srcs: (13, 7)(1635) -1 --> (1635) -1:PUGB6, pass, NI0
			10'd7 : rdata = 48'b110001110000110100000000000100000000000000000000;
			// PEs: 48 -> 26
			// srcs: (14, 8)(1636) 0 --> (1636) 0:PUGB6, pass, PEGB2
			10'd8 : rdata = 48'b110001110000110100000000000000000000000010100000;
			// PEs: 48 -> 24
			// srcs: (15, 10)(1638) 0 --> (1638) 0:PUGB6, pass, NI1
			10'd9 : rdata = 48'b110001110000110100000000000100001000000000000000;
			// PEs: 48 -> 27
			// srcs: (16, 11)(1639) 3 --> (1639) 3:PUGB6, pass, PEGB3
			10'd10 : rdata = 48'b110001110000110100000000000000000000000010110000;
			// PEs: 48 -> 24
			// srcs: (17, 13)(1641) -6 --> (1641) -6:PUGB6, pass, NI2
			10'd11 : rdata = 48'b110001110000110100000000000100010000000000000000;
			// PEs: 56 -> 28
			// srcs: (18, 14)(1642) 1 --> (1642) 1:PUGB7, pass, PEGB4
			10'd12 : rdata = 48'b110001110000111100000000000000000000000011000000;
			// PEs: 56 -> 24
			// srcs: (19, 16)(1644) -1 --> (1644) -1:PUGB7, pass, NI3
			10'd13 : rdata = 48'b110001110000111100000000000100011000000000000000;
			// PEs: 56 -> 29
			// srcs: (20, 17)(1645) -4 --> (1645) -4:PUGB7, pass, PEGB5
			10'd14 : rdata = 48'b110001110000111100000000000000000000000011010000;
			// PEs: 56 -> 24
			// srcs: (21, 19)(1647) 2 --> (1647) 2:PUGB7, pass, NI4
			10'd15 : rdata = 48'b110001110000111100000000000100100000000000000000;
			// PEs: 56 -> 30
			// srcs: (22, 20)(1648) -6 --> (1648) -6:PUGB7, pass, PEGB6
			10'd16 : rdata = 48'b110001110000111100000000000000000000000011100000;
			// PEs: 24 -> 26
			// srcs: (23, 9)(1635) -1 --> (1635) -1:NI0, pass, PEGB2
			10'd17 : rdata = 48'b110001010000000000000000000000000000000010100000;
			// PEs: 56 -> 24
			// srcs: (24, 22)(1650) 9 --> (1650) 9:PUGB7, pass, NI0
			10'd18 : rdata = 48'b110001110000111100000000000100000000000000000000;
			// PEs: 24 -> 27
			// srcs: (25, 12)(1638) 0 --> (1638) 0:NI1, pass, PEGB3
			10'd19 : rdata = 48'b110001010000000100000000000000000000000010110000;
			// PEs: 56 -> 31
			// srcs: (26, 23)(1651) -2 --> (1651) -2:PUGB7, pass, PEGB7
			10'd20 : rdata = 48'b110001110000111100000000000000000000000011110000;
			// PEs: 24 -> 28
			// srcs: (27, 15)(1641) -6 --> (1641) -6:NI2, pass, PEGB4
			10'd21 : rdata = 48'b110001010000001000000000000000000000000011000000;
			// PEs: 0 -> 24
			// srcs: (28, 25)(1656) 0 --> (1656) 0:PUGB0, pass, NI1
			10'd22 : rdata = 48'b110001110000000100000000000100001000000000000000;
			// PEs: 24 -> 29
			// srcs: (29, 18)(1644) -1 --> (1644) -1:NI3, pass, PEGB5
			10'd23 : rdata = 48'b110001010000001100000000000000000000000011010000;
			// PEs: 0 -> 25
			// srcs: (30, 26)(1657) 1 --> (1657) 1:PUGB0, pass, PENB
			10'd24 : rdata = 48'b110001110000000100000000000000000000000100000000;
			// PEs: 24 -> 30
			// srcs: (31, 21)(1647) 2 --> (1647) 2:NI4, pass, PEGB6
			10'd25 : rdata = 48'b110001010000010000000000000000000000000011100000;
			// PEs: 25 -> 32
			// srcs: (32, 28)(1682) -2 --> (1682) -2:PEGB1, pass, PUNB
			10'd26 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 26 -> 32
			// srcs: (33, 29)(1684) 1 --> (1684) 1:PEGB2, pass, PUNB
			10'd27 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 27 -> 32
			// srcs: (34, 30)(1685) 0 --> (1685) 0:PEGB3, pass, PUNB
			10'd28 : rdata = 48'b110001110000011000000000000000000000001000000000;
			// PEs: 24 -> 31
			// srcs: (35, 24)(1650) 9 --> (1650) 9:NI0, pass, PEGB7
			10'd29 : rdata = 48'b110001010000000000000000000000000000000011110000;
			// PEs: 24 -> 25
			// srcs: (36, 27)(1656) 0 --> (1656) 0:NI1, pass, PENB
			10'd30 : rdata = 48'b110001010000000100000000000000000000000100000000;
			// PEs: 28 -> 32
			// srcs: (37, 31)(1687) -2 --> (1687) -2:PEGB4, pass, PUNB
			10'd31 : rdata = 48'b110001110000100000000000000000000000001000000000;
			// PEs: 29 -> 32
			// srcs: (38, 32)(1688) -3 --> (1688) -3:PEGB5, pass, PUNB
			10'd32 : rdata = 48'b110001110000101000000000000000000000001000000000;
			// PEs: 30 -> 32
			// srcs: (39, 33)(1690) 9 --> (1690) 9:PEGB6, pass, PUNB
			10'd33 : rdata = 48'b110001110000110000000000000000000000001000000000;
			// PEs: 31 -> 32
			// srcs: (40, 34)(1691) 6 --> (1691) 6:PENB, pass, PUNB
			10'd34 : rdata = 48'b110001101111111000000000000000000000001000000000;
			// PEs: 25 -> 32
			// srcs: (41, 41)(1764) 0 --> (1764) 0:PEGB1, pass, PUNB
			10'd35 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 26 -> 32
			// srcs: (42, 42)(1766) -3 --> (1766) -3:PEGB2, pass, PUNB
			10'd36 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 16 -> 24
			// srcs: (43, 35)(1757) -4 --> (1757) -4:PUNB, pass, NI0
			10'd37 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 16 -> 26
			// srcs: (44, 36)(1758) 0 --> (1758) 0:PUNB, pass, PEGB2
			10'd38 : rdata = 48'b110001101111111100000000000000000000000010100000;
			// PEs: 16 -> 24
			// srcs: (45, 38)(1760) -4 --> (1760) -4:PUNB, pass, NI1
			10'd39 : rdata = 48'b110001101111111100000000000100001000000000000000;
			// PEs: 16 -> 27
			// srcs: (46, 39)(1761) -1 --> (1761) -1:PUNB, pass, PEGB3
			10'd40 : rdata = 48'b110001101111111100000000000000000000000010110000;
			// PEs: 27 -> 32
			// srcs: (47, 43)(1767) 0 --> (1767) 0:PEGB3, pass, PUNB
			10'd41 : rdata = 48'b110001110000011000000000000000000000001000000000;
			// PEs: 40 -> 24
			// srcs: (48, 44)(1791) 0 --> (1791) 0:PUGB5, pass, NI2
			10'd42 : rdata = 48'b110001110000101100000000000100010000000000000000;
			// PEs: 40 -> 25
			// srcs: (49, 45)(1792) 0 --> (1792) 0:PUGB5, pass, PENB
			10'd43 : rdata = 48'b110001110000101100000000000000000000000100000000;
			// PEs: 16 -> 24
			// srcs: (50, 47)(1834) 0 --> (1834) 0:PUNB, pass, NI3
			10'd44 : rdata = 48'b110001101111111100000000000100011000000000000000;
			// PEs: 16 -> 28
			// srcs: (51, 48)(1835) -2 --> (1835) -2:PUNB, pass, PEGB4
			10'd45 : rdata = 48'b110001101111111100000000000000000000000011000000;
			// PEs: 25 -> 32
			// srcs: (52, 56)(1844) 9 --> (1844) 9:PEGB1, pass, PUNB
			10'd46 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 24 -> 26
			// srcs: (53, 37)(1757) -4 --> (1757) -4:NI0, pass, PEGB2
			10'd47 : rdata = 48'b110001010000000000000000000000000000000010100000;
			// PEs: 16 -> 24
			// srcs: (54, 50)(1837) 1 --> (1837) 1:PUNB, pass, NI0
			10'd48 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 24 -> 27
			// srcs: (55, 40)(1760) -4 --> (1760) -4:NI1, pass, PEGB3
			10'd49 : rdata = 48'b110001010000000100000000000000000000000010110000;
			// PEs: 24 -> 25
			// srcs: (56, 46)(1791) 0 --> (1791) 0:NI2, pass, PENB
			10'd50 : rdata = 48'b110001010000001000000000000000000000000100000000;
			// PEs: 26 -> 32
			// srcs: (57, 57)(1846) 0 --> (1846) 0:PEGB2, pass, PUNB
			10'd51 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 16 -> 29
			// srcs: (58, 51)(1838) 3 --> (1838) 3:PUNB, pass, PEGB5
			10'd52 : rdata = 48'b110001101111111100000000000000000000000011010000;
			// PEs: 16 -> 24
			// srcs: (59, 53)(1840) -1 --> (1840) -1:PUNB, pass, NI1
			10'd53 : rdata = 48'b110001101111111100000000000100001000000000000000;
			// PEs: 24 -> 28
			// srcs: (60, 49)(1834) 0 --> (1834) 0:NI3, pass, PEGB4
			10'd54 : rdata = 48'b110001010000001100000000000000000000000011000000;
			// PEs: 16 -> 30
			// srcs: (61, 54)(1841) -1 --> (1841) -1:PUNB, pass, PEGB6
			10'd55 : rdata = 48'b110001101111111100000000000000000000000011100000;
			// PEs: 27 -> 32
			// srcs: (62, 58)(1847) 0 --> (1847) 0:PEGB3, pass, PUNB
			10'd56 : rdata = 48'b110001110000011000000000000000000000001000000000;
			// PEs: 28 -> 32
			// srcs: (63, 59)(1849) 0 --> (1849) 0:PEGB4, pass, PUNB
			10'd57 : rdata = 48'b110001110000100000000000000000000000001000000000;
			// PEs: 29 -> 32
			// srcs: (64, 60)(1850) 3 --> (1850) 3:PEGB5, pass, PUNB
			10'd58 : rdata = 48'b110001110000101000000000000000000000001000000000;
			// PEs: 30 -> 32
			// srcs: (65, 61)(1852) 2 --> (1852) 2:PEGB6, pass, PUNB
			10'd59 : rdata = 48'b110001110000110000000000000000000000001000000000;
			// PEs: 31 -> 32
			// srcs: (66, 62)(1853) -2 --> (1853) -2:PENB, pass, PUNB
			10'd60 : rdata = 48'b110001101111111000000000000000000000001000000000;
			// PEs: 24 -> 29
			// srcs: (67, 52)(1837) 1 --> (1837) 1:NI0, pass, PEGB5
			10'd61 : rdata = 48'b110001010000000000000000000000000000000011010000;
			// PEs: 16 -> 24
			// srcs: (68, 63)(1920) 6 --> (1920) 6:PUNB, pass, NI0
			10'd62 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 26 -> 32
			// srcs: (69, 67)(1926) -2 --> (1926) -2:PEGB2, pass, PUNB
			10'd63 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 24 -> 30
			// srcs: (70, 55)(1840) -1 --> (1840) -1:NI1, pass, PEGB6
			10'd64 : rdata = 48'b110001010000000100000000000000000000000011100000;
			// PEs: 27 -> 32
			// srcs: (71, 68)(1927) -2 --> (1927) -2:PEGB3, pass, PUNB
			10'd65 : rdata = 48'b110001110000011000000000000000000000001000000000;
			// PEs: 28 -> 32
			// srcs: (72, 69)(1929) 2 --> (1929) 2:PEGB4, pass, PUNB
			10'd66 : rdata = 48'b110001110000100000000000000000000000001000000000;
			// PEs: 16 -> 25
			// srcs: (73, 64)(1921) -6 --> (1921) -6:PUNB, pass, PENB
			10'd67 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 29 -> 32
			// srcs: (74, 70)(1930) -3 --> (1930) -3:PEGB5, pass, PUNB
			10'd68 : rdata = 48'b110001110000101000000000000000000000001000000000;
			// PEs: 30 -> 32
			// srcs: (75, 71)(1932) -4 --> (1932) -4:PEGB6, pass, PUNB
			10'd69 : rdata = 48'b110001110000110000000000000000000000001000000000;
			// PEs: 31 -> 32
			// srcs: (76, 72)(1933) 0 --> (1933) 0:PENB, pass, PUNB
			10'd70 : rdata = 48'b110001101111111000000000000000000000001000000000;
			// PEs: 26 -> 32
			// srcs: (77, 83)(2008) 0 --> (2008) 0:PEGB2, pass, PUNB
			10'd71 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 16 -> 31
			// srcs: (78, 66)(1923) -6 --> (1923) -6:PUNB, pass, PEGB7
			10'd72 : rdata = 48'b110001101111111100000000000000000000000011110000;
			// PEs: 24 -> 25
			// srcs: (79, 65)(1920) 6 --> (1920) 6:NI0, pass, PENB
			10'd73 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 16 -> 24
			// srcs: (80, 73)(1996) 3 --> (1996) 3:PUNB, pass, NI0
			10'd74 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 27 -> 32
			// srcs: (81, 84)(2009) -3 --> (2009) -3:PEGB3, pass, PUNB
			10'd75 : rdata = 48'b110001110000011000000000000000000000001000000000;
			// PEs: 28 -> 32
			// srcs: (82, 85)(2011) -6 --> (2011) -6:PEGB4, pass, PUNB
			10'd76 : rdata = 48'b110001110000100000000000000000000000001000000000;
			// PEs: 29 -> 32
			// srcs: (83, 86)(2012) -4 --> (2012) -4:PEGB5, pass, PUNB
			10'd77 : rdata = 48'b110001110000101000000000000000000000001000000000;
			// PEs: 26 -> 32
			// srcs: (84, 97)(2088) -2 --> (2088) -2:PEGB2, pass, PUNB
			10'd78 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 16 -> 25
			// srcs: (85, 74)(1997) -6 --> (1997) -6:PUNB, pass, PENB
			10'd79 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 27 -> 32
			// srcs: (86, 98)(2089) 0 --> (2089) 0:PEGB3, pass, PUNB
			10'd80 : rdata = 48'b110001110000011000000000000000000000001000000000;
			// PEs: 28 -> 32
			// srcs: (87, 99)(2091) 0 --> (2091) 0:PEGB4, pass, PUNB
			10'd81 : rdata = 48'b110001110000100000000000000000000000001000000000;
			// PEs: 29 -> 32
			// srcs: (88, 100)(2092) 0 --> (2092) 0:PEGB5, pass, PUNB
			10'd82 : rdata = 48'b110001110000101000000000000000000000001000000000;
			// PEs: 30 -> 32
			// srcs: (89, 101)(2094) 4 --> (2094) 4:PEGB6, pass, PUNB
			10'd83 : rdata = 48'b110001110000110000000000000000000000001000000000;
			// PEs: 31 -> 32
			// srcs: (90, 102)(2095) 0 --> (2095) 0:PENB, pass, PUNB
			10'd84 : rdata = 48'b110001101111111000000000000000000000001000000000;
			// PEs: 24 -> 25
			// srcs: (91, 75)(1996) 3 --> (1996) 3:NI0, pass, PENB
			10'd85 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 16 -> 24
			// srcs: (92, 76)(1999) 2 --> (1999) 2:PUNB, pass, NI0
			10'd86 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 16 -> 25
			// srcs: (93, 77)(2000) 6 --> (2000) 6:PUNB, pass, PENB
			10'd87 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 26 -> 32
			// srcs: (94, 107)(2168) 0 --> (2168) 0:PEGB2, pass, PUNB
			10'd88 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 27 -> 32
			// srcs: (95, 108)(2169) -2 --> (2169) -2:PEGB3, pass, PUNB
			10'd89 : rdata = 48'b110001110000011000000000000000000000001000000000;
			// PEs: 28 -> 32
			// srcs: (96, 109)(2171) 4 --> (2171) 4:PEGB4, pass, PUNB
			10'd90 : rdata = 48'b110001110000100000000000000000000000001000000000;
			// PEs: 29 -> 32
			// srcs: (97, 110)(2172) 0 --> (2172) 0:PEGB5, pass, PUNB
			10'd91 : rdata = 48'b110001110000101000000000000000000000001000000000;
			// PEs: 30 -> 32
			// srcs: (98, 111)(2174) 3 --> (2174) 3:PEGB6, pass, PUNB
			10'd92 : rdata = 48'b110001110000110000000000000000000000001000000000;
			// PEs: 24 -> 25
			// srcs: (99, 78)(1999) 2 --> (1999) 2:NI0, pass, PENB
			10'd93 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 16 -> 24
			// srcs: (100, 79)(2002) -4 --> (2002) -4:PUNB, pass, NI0
			10'd94 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 16 -> 25
			// srcs: (101, 80)(2003) 2 --> (2003) 2:PUNB, pass, PENB
			10'd95 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 16 -> 26
			// srcs: (102, 82)(2005) 1 --> (2005) 1:PUNB, pass, PEGB2
			10'd96 : rdata = 48'b110001101111111100000000000000000000000010100000;
			// PEs: 31 -> 32
			// srcs: (103, 112)(2175) 6 --> (2175) 6:PENB, pass, PUNB
			10'd97 : rdata = 48'b110001101111111000000000000000000000001000000000;
			// PEs: 28 -> 0
			// srcs: (104, 141)(2422) -5 --> (2422) -5:PEGB4, pass, PUGB0
			10'd98 : rdata = 48'b110001110000100000000000000000000000000000001000;
			// PEs: 29 -> 16
			// srcs: (105, 142)(2424) -5 --> (2424) -5:PEGB5, pass, PUGB2
			10'd99 : rdata = 48'b110001110000101000000000000000000000000000001010;
			// PEs: 31 -> 8
			// srcs: (106, 144)(2431) 7 --> (2431) 7:PENB, pass, PUGB1
			10'd100 : rdata = 48'b110001101111111000000000000000000000000000001001;
			// PEs: 24 -> 25
			// srcs: (107, 81)(2002) -4 --> (2002) -4:NI0, pass, PENB
			10'd101 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 16 -> 24
			// srcs: (108, 87)(2076) 0 --> (2076) 0:PUNB, pass, NI0
			10'd102 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 16 -> 25
			// srcs: (109, 88)(2077) 1 --> (2077) 1:PUNB, pass, PENB
			10'd103 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 25 -> 40
			// srcs: (110, 145)(2436) 1 --> (2436) 1:PEGB1, pass, PUGB5
			10'd104 : rdata = 48'b110001110000001000000000000000000000000000001101;
			// PEs: 28 -> 32
			// srcs: (111, 118)(1769) -2 --> (1769) -2:PEGB4, pass, PUNB
			10'd105 : rdata = 48'b110001110000100000000000000000000000001000000000;
			// PEs: 26 -> 40
			// srcs: (112, 151)(1701) -1 --> (1701) -1:PEGB2, pass, PUGB5
			10'd106 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 27 -> 0
			// srcs: (113, 152)(1704) -2 --> (1704) -2:PEGB3, pass, PUGB0
			10'd107 : rdata = 48'b110001110000011000000000000000000000000000001000;
			// PEs: 30 -> 56
			// srcs: (114, 155)(1713) -2 --> (1713) -2:PEGB6, pass, PUGB7
			10'd108 : rdata = 48'b110001110000110000000000000000000000000000001111;
			// PEs: 24 -> 25
			// srcs: (115, 89)(2076) 0 --> (2076) 0:NI0, pass, PENB
			10'd109 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 16 -> 24
			// srcs: (116, 90)(2079) 0 --> (2079) 0:PUNB, pass, NI0
			10'd110 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 16 -> 25
			// srcs: (117, 91)(2080) 0 --> (2080) 0:PUNB, pass, PENB
			10'd111 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 30 -> 56
			// srcs: (118, 171)(2619) -2 --> (2619) -2:PEGB6, pass, PUGB7
			10'd112 : rdata = 48'b110001110000110000000000000000000000000000001111;
			// PEs: 29 -> 32
			// srcs: (119, 119)(1770) 0 --> (1770) 0:PEGB5, pass, PUNB
			10'd113 : rdata = 48'b110001110000101000000000000000000000001000000000;
			// PEs: 28 -> 16
			// srcs: (121, 153)(1707) 9 --> (1707) 9:PEGB4, pass, PUGB2
			10'd114 : rdata = 48'b110001110000100000000000000000000000000000001010;
			// PEs: 29 -> 40
			// srcs: (122, 154)(1710) 2 --> (1710) 2:PEGB5, pass, PUGB5
			10'd115 : rdata = 48'b110001110000101000000000000000000000000000001101;
			// PEs: 24 -> 25
			// srcs: (123, 92)(2079) 0 --> (2079) 0:NI0, pass, PENB
			10'd116 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 16 -> 24
			// srcs: (124, 93)(2082) 2 --> (2082) 2:PUNB, pass, NI0
			10'd117 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 16 -> 25
			// srcs: (125, 94)(2083) 0 --> (2083) 0:PUNB, pass, PENB
			10'd118 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 16 -> 27
			// srcs: (126, 96)(2085) 0 --> (2085) 0:PUNB, pass, PEGB3
			10'd119 : rdata = 48'b110001101111111100000000000000000000000010110000;
			// PEs: 30 -> 32
			// srcs: (127, 120)(1771) 1 --> (1771) 1:PEGB6, pass, PUNB
			10'd120 : rdata = 48'b110001110000110000000000000000000000001000000000;
			// PEs: 31 -> 0
			// srcs: (128, 156)(1716) -2 --> (1716) -2:PENB, pass, PUGB0
			10'd121 : rdata = 48'b110001101111111000000000000000000000000000001000;
			// PEs: 26 -> 16
			// srcs: (129, 163)(2537) -4 --> (2537) -4:PEGB2, pass, PUGB2
			10'd122 : rdata = 48'b110001110000010000000000000000000000000000001010;
			// PEs: 25 -> 40
			// srcs: (130, 165)(2571) 0 --> (2571) 0:PEGB1, pass, PUGB5
			10'd123 : rdata = 48'b110001110000001000000000000000000000000000001101;
			// PEs: 24 -> 25
			// srcs: (131, 95)(2082) 2 --> (2082) 2:NI0, pass, PENB
			10'd124 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 16 -> 24
			// srcs: (132, 103)(2158) 0 --> (2158) 0:PUNB, pass, NI0
			10'd125 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 16 -> 25
			// srcs: (133, 104)(2159) -3 --> (2159) -3:PUNB, pass, PENB
			10'd126 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 31 -> 32
			// srcs: (134, 121)(1772) 0 --> (1772) 0:PENB, pass, PUNB
			10'd127 : rdata = 48'b110001101111111000000000000000000000001000000000;
			// PEs: 28 -> 48
			// srcs: (135, 181)(1891) 2 --> (1891) 2:PEGB4, pass, PUGB6
			10'd128 : rdata = 48'b110001110000100000000000000000000000000000001110;
			// PEs: 29 -> 56
			// srcs: (136, 182)(1894) 4 --> (1894) 4:PEGB5, pass, PUGB7
			10'd129 : rdata = 48'b110001110000101000000000000000000000000000001111;
			// PEs: 30 -> 8
			// srcs: (137, 183)(1897) -2 --> (1897) -2:PEGB6, pass, PUGB1
			10'd130 : rdata = 48'b110001110000110000000000000000000000000000001001;
			// PEs: 25 -> 8
			// srcs: (138, 193)(2777) -3 --> (2777) -3:PEGB1, pass, PUGB1
			10'd131 : rdata = 48'b110001110000001000000000000000000000000000001001;
			// PEs: 24 -> 25
			// srcs: (139, 105)(2158) 0 --> (2158) 0:NI0, pass, PENB
			10'd132 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 16 -> 25
			// srcs: (140, 106)(2165) 0 --> (2165) 0:PUNB, pass, PENB
			10'd133 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 16 -> 25
			// srcs: (141, 113)(2247) -2 --> (2247) -2:PUNB, pass, PENB
			10'd134 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 16 -> 25
			// srcs: (142, 114)(2327) 0 --> (2327) 0:PUNB, pass, PENB
			10'd135 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 30 -> 32
			// srcs: (143, 128)(2014) 0 --> (2014) 0:PEGB6, pass, PUNB
			10'd136 : rdata = 48'b110001110000110000000000000000000000001000000000;
			// PEs: 28 -> 40
			// srcs: (144, 169)(2614) -2 --> (2614) -2:PEGB4, pass, PUGB5
			10'd137 : rdata = 48'b110001110000100000000000000000000000000000001101;
			// PEs: 29 -> 16
			// srcs: (145, 170)(2617) 4 --> (2617) 4:PEGB5, pass, PUGB2
			10'd138 : rdata = 48'b110001110000101000000000000000000000000000001010;
			// PEs: 26 -> 0
			// srcs: (146, 179)(1885) -2 --> (1885) -2:PEGB2, pass, PUGB0
			10'd139 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 27 -> 40
			// srcs: (147, 180)(1888) -2 --> (1888) -2:PEGB3, pass, PUGB5
			10'd140 : rdata = 48'b110001110000011000000000000000000000000000001101;
			// PEs: 31 -> 32
			// srcs: (148, 129)(2015) 4 --> (2015) 4:PENB, pass, PUNB
			10'd141 : rdata = 48'b110001101111111000000000000000000000001000000000;
			// PEs: 27 -> 32
			// srcs: (149, 140)(2419) 3 --> (2419) 3:PEGB3, pass, PUNB
			10'd142 : rdata = 48'b110001110000011000000000000000000000001000000000;
			// PEs: 25 -> 56
			// srcs: (150, 194)(2779) 8 --> (2779) 8:PEGB1, pass, PUGB7
			10'd143 : rdata = 48'b110001110000001000000000000000000000000000001111;
			// PEs: 25 -> 8
			// srcs: (151, 195)(2783) -2 --> (2783) -2:PEGB1, pass, PUGB1
			10'd144 : rdata = 48'b110001110000001000000000000000000000000000001001;
			// PEs: 31 -> 16
			// srcs: (154, 184)(1900) 0 --> (1900) 0:PENB, pass, PUGB2
			10'd145 : rdata = 48'b110001101111111000000000000000000000000000001010;
			// PEs: 25 -> 16
			// srcs: (155, 225)(3105) -1 --> (3105) -1:PEGB1, pass, PUGB2
			10'd146 : rdata = 48'b110001110000001000000000000000000000000000001010;
			// PEs: 25 -> 32
			// srcs: (157, 150)(1698) -4 --> (1698) -4:PEGB1, pass, PUNB
			10'd147 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 26 -> 48
			// srcs: (159, 196)(2785) 4 --> (2785) 4:PEGB2, pass, PUGB6
			10'd148 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 28 -> 8
			// srcs: (160, 228)(3114) 4 --> (3114) 4:PEGB4, pass, PUGB1
			10'd149 : rdata = 48'b110001110000100000000000000000000000000000001001;
			// PEs: 25 -> 32
			// srcs: (165, 178)(1882) 0 --> (1882) 0:PEGB1, pass, PUNB
			10'd150 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 25 -> 48
			// srcs: (167, 211)(2935) -3 --> (2935) -3:PEGB1, pass, PUGB6
			10'd151 : rdata = 48'b110001110000001000000000000000000000000000001110;
			// PEs: 31 -> 48
			// srcs: (172, 218)(2268) 1 --> (2268) 1:PENB, pass, PUGB6
			10'd152 : rdata = 48'b110001101111111000000000000000000000000000001110;
			// PEs: 25 -> 32
			// srcs: (173, 185)(2700) 0 --> (2700) 0:PEGB1, pass, PUNB
			10'd153 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 31 -> 32
			// srcs: (178, 186)(2703) -8 --> (2703) -8:PENB, pass, PUNB
			10'd154 : rdata = 48'b110001101111111000000000000000000000001000000000;
			// PEs: 27 -> 32
			// srcs: (179, 207)(2864) 3 --> (2864) 3:PEGB3, pass, PUNB
			10'd155 : rdata = 48'b110001110000011000000000000000000000001000000000;
			// PEs: 31 -> 48
			// srcs: (180, 226)(3107) -6 --> (3107) -6:PENB, pass, PUGB6
			10'd156 : rdata = 48'b110001101111111000000000000000000000000000001110;
			// PEs: 25 -> 32
			// srcs: (187, 212)(2946) 0 --> (2946) 0:PEGB1, pass, PUNB
			10'd157 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 30 -> 32
			// srcs: (195, 217)(2265) 2 --> (2265) 2:PEGB6, pass, PUNB
			10'd158 : rdata = 48'b110001110000110000000000000000000000001000000000;
			// PEs: 16 -> 24
			// srcs: (227, 115)(1673) 0 --> (1673) 0:PUNB, pass, NI0
			10'd159 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 16 -> 27
			// srcs: (243, 116)(1674) 0 --> (1674) 0:PUNB, pass, PEGB3
			10'd160 : rdata = 48'b110001101111111100000000000000000000000010110000;
			// PEs: 24 -> 27
			// srcs: (252, 117)(1673) 0 --> (1673) 0:NI0, pass, PEGB3
			10'd161 : rdata = 48'b110001010000000000000000000000000000000010110000;
			// PEs: 16 -> 24
			// srcs: (256, 122)(1916) 2 --> (1916) 2:PUNB, pass, NI0
			10'd162 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 16 -> 25
			// srcs: (272, 123)(1917) 0 --> (1917) 0:PUNB, pass, PENB
			10'd163 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (278, 124)(1916) 2 --> (1916) 2:NI0, pass, PENB
			10'd164 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 16 -> 24
			// srcs: (288, 125)(1918) 1 --> (1918) 1:PUNB, pass, NI0
			10'd165 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 16 -> 25
			// srcs: (304, 126)(1919) 4 --> (1919) 4:PUNB, pass, PENB
			10'd166 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (310, 127)(1918) 1 --> (1918) 1:NI0, pass, PENB
			10'd167 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 16 -> 24
			// srcs: (317, 130)(2161) 0 --> (2161) 0:PUNB, pass, NI0
			10'd168 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 16 -> 25
			// srcs: (333, 131)(2162) 4 --> (2162) 4:PUNB, pass, PENB
			10'd169 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (339, 132)(2161) 0 --> (2161) 0:NI0, pass, PENB
			10'd170 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 16 -> 24
			// srcs: (340, 133)(2163) 3 --> (2163) 3:PUNB, pass, NI0
			10'd171 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 16 -> 25
			// srcs: (341, 134)(2164) 4 --> (2164) 4:PUNB, pass, PENB
			10'd172 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (347, 135)(2163) 3 --> (2163) 3:NI0, pass, PENB
			10'd173 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 8 -> 24
			// srcs: (348, 136)(2386) -3 --> (2386) -3:PUGB1, pass, NI0
			10'd174 : rdata = 48'b110001110000001100000000000100000000000000000000;
			// PEs: 56 -> 25
			// srcs: (349, 137)(1606) 6 --> (1606) 6:PUGB7, pass, PENB
			10'd175 : rdata = 48'b110001110000111100000000000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (355, 138)(2386) -3 --> (2386) -3:NI0, pass, PENB
			10'd176 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 0 -> 25
			// srcs: (356, 139)(1637) 0 --> (1637) 0:PUGB0, pass, PENB
			10'd177 : rdata = 48'b110001110000000100000000000000000000000100000000;
			// PEs: 0 -> 25
			// srcs: (357, 143)(1649) 0 --> (1649) 0:PUGB0, pass, PENB
			10'd178 : rdata = 48'b110001110000000100000000000000000000000100000000;
			// PEs: 16 -> 25
			// srcs: (358, 146)(2454) 3 --> (2454) 3:PUNB, pass, PENB
			10'd179 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 32 -> 24
			// srcs: (359, 147)(2466) 1 --> (2466) 1:PUGB4, pass, NI0
			10'd180 : rdata = 48'b110001110000100100000000000100000000000000000000;
			// PEs: 25 -> 32
			// srcs: (362, 232)(2387) 3 --> (2387) 3:PEGB1, pass, PUNB
			10'd181 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 25 -> 32
			// srcs: (363, 236)(2418) -1 --> (2418) -1:PEGB1, pass, PUNB
			10'd182 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 16 -> 25
			// srcs: (522, 148)(1686) -1 --> (1686) -1:PUNB, pass, PENB
			10'd183 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (528, 149)(2466) 1 --> (2466) 1:NI0, pass, PENB
			10'd184 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 0 -> 24
			// srcs: (529, 157)(2505) 8 --> (2505) 8:PUGB0, pass, NI0
			10'd185 : rdata = 48'b110001110000000100000000000100000000000000000000;
			// PEs: 32 -> 25
			// srcs: (530, 158)(1726) 6 --> (1726) 6:PUGB4, pass, PENB
			10'd186 : rdata = 48'b110001110000100100000000000000000000000100000000;
			// PEs: 25 -> 48
			// srcs: (535, 239)(2467) 0 --> (2467) 0:PEGB1, pass, PUGB6
			10'd187 : rdata = 48'b110001110000001000000000000000000000000000001110;
			// PEs: 24 -> 25
			// srcs: (536, 159)(2505) 8 --> (2505) 8:NI0, pass, PENB
			10'd188 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 0 -> 24
			// srcs: (537, 160)(2526) 0 --> (2526) 0:PUGB0, pass, NI0
			10'd189 : rdata = 48'b110001110000000100000000000100000000000000000000;
			// PEs: 40 -> 25
			// srcs: (538, 161)(1747) 0 --> (1747) 0:PUGB5, pass, PENB
			10'd190 : rdata = 48'b110001110000101100000000000000000000000100000000;
			// PEs: 25 -> 32
			// srcs: (543, 243)(2506) 14 --> (2506) 14:PEGB1, pass, PUNB
			10'd191 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 24 -> 25
			// srcs: (544, 162)(2526) 0 --> (2526) 0:NI0, pass, PENB
			10'd192 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 40 -> 25
			// srcs: (545, 164)(1762) 0 --> (1762) 0:PUGB5, pass, PENB
			10'd193 : rdata = 48'b110001110000101100000000000000000000000100000000;
			// PEs: 16 -> 24
			// srcs: (546, 166)(2612) 6 --> (2612) 6:PUNB, pass, NI0
			10'd194 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 0 -> 25
			// srcs: (547, 167)(1833) 0 --> (1833) 0:PUGB0, pass, PENB
			10'd195 : rdata = 48'b110001110000000100000000000000000000000100000000;
			// PEs: 25 -> 32
			// srcs: (551, 244)(2527) 0 --> (2527) 0:PEGB1, pass, PUNB
			10'd196 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 26 -> 32
			// srcs: (552, 255)(2699) 7 --> (2699) 7:PEGB2, pass, PUNB
			10'd197 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 24 -> 25
			// srcs: (558, 168)(2612) 6 --> (2612) 6:NI0, pass, PENB
			10'd198 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 32 -> 24
			// srcs: (559, 172)(2624) 10 --> (2624) 10:PUGB4, pass, NI0
			10'd199 : rdata = 48'b110001110000100100000000000100000000000000000000;
			// PEs: 8 -> 25
			// srcs: (560, 173)(1845) 0 --> (1845) 0:PUGB1, pass, PENB
			10'd200 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 25 -> 56
			// srcs: (565, 249)(2613) 6 --> (2613) 6:PEGB1, pass, PUGB7
			10'd201 : rdata = 48'b110001110000001000000000000000000000000000001111;
			// PEs: 24 -> 25
			// srcs: (566, 174)(2624) 10 --> (2624) 10:NI0, pass, PENB
			10'd202 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 40 -> 24
			// srcs: (567, 175)(2640) 1 --> (2640) 1:PUGB5, pass, NI0
			10'd203 : rdata = 48'b110001110000101100000000000100000000000000000000;
			// PEs: 16 -> 25
			// srcs: (568, 176)(1863) 6 --> (1863) 6:PUNB, pass, PENB
			10'd204 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 25 -> 0
			// srcs: (573, 250)(2625) 10 --> (2625) 10:PEGB1, pass, PUGB0
			10'd205 : rdata = 48'b110001110000001000000000000000000000000000001000;
			// PEs: 24 -> 25
			// srcs: (574, 177)(2640) 1 --> (2640) 1:NI0, pass, PENB
			10'd206 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 8 -> 24
			// srcs: (575, 187)(2760) 0 --> (2760) 0:PUGB1, pass, NI0
			10'd207 : rdata = 48'b110001110000001100000000000100000000000000000000;
			// PEs: 56 -> 25
			// srcs: (576, 188)(1980) 0 --> (1980) 0:PUGB7, pass, PENB
			10'd208 : rdata = 48'b110001110000111100000000000000000000000100000000;
			// PEs: 25 -> 40
			// srcs: (581, 251)(2641) 7 --> (2641) 7:PEGB1, pass, PUGB5
			10'd209 : rdata = 48'b110001110000001000000000000000000000000000001101;
			// PEs: 24 -> 25
			// srcs: (582, 189)(2760) 0 --> (2760) 0:NI0, pass, PENB
			10'd210 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 16 -> 24
			// srcs: (583, 190)(2772) -1 --> (2772) -1:PUNB, pass, NI0
			10'd211 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 56 -> 25
			// srcs: (584, 191)(1992) 4 --> (1992) 4:PUGB7, pass, PENB
			10'd212 : rdata = 48'b110001110000111100000000000000000000000100000000;
			// PEs: 25 -> 8
			// srcs: (589, 256)(2761) 0 --> (2761) 0:PEGB1, pass, PUGB1
			10'd213 : rdata = 48'b110001110000001000000000000000000000000000001001;
			// PEs: 24 -> 25
			// srcs: (590, 192)(2772) -1 --> (2772) -1:NI0, pass, PENB
			10'd214 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 56 -> 24
			// srcs: (591, 197)(2820) 3 --> (2820) 3:PUGB7, pass, NI0
			10'd215 : rdata = 48'b110001110000111100000000000100000000000000000000;
			// PEs: 16 -> 25
			// srcs: (592, 198)(2041) 2 --> (2041) 2:PUNB, pass, PENB
			10'd216 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 25 -> 32
			// srcs: (597, 257)(2773) 3 --> (2773) 3:PEGB1, pass, PUNB
			10'd217 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 24 -> 25
			// srcs: (598, 199)(2820) 3 --> (2820) 3:NI0, pass, PENB
			10'd218 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 0 -> 24
			// srcs: (599, 200)(2831) -4 --> (2831) -4:PUGB0, pass, NI0
			10'd219 : rdata = 48'b110001110000000100000000000100000000000000000000;
			// PEs: 16 -> 25
			// srcs: (600, 201)(2053) 4 --> (2053) 4:PUNB, pass, PENB
			10'd220 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 25 -> 32
			// srcs: (605, 261)(2821) 5 --> (2821) 5:PEGB1, pass, PUNB
			10'd221 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 24 -> 25
			// srcs: (606, 202)(2831) -4 --> (2831) -4:NI0, pass, PENB
			10'd222 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 8 -> 25
			// srcs: (607, 203)(2838) -8 --> (2838) -8:PUGB1, pass, PENB
			10'd223 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 16 -> 25
			// srcs: (608, 204)(2848) -1 --> (2848) -1:PUNB, pass, PENB
			10'd224 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 16 -> 25
			// srcs: (609, 205)(2851) 6 --> (2851) 6:PUNB, pass, PENB
			10'd225 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 16 -> 25
			// srcs: (610, 206)(2853) 6 --> (2853) 6:PUNB, pass, PENB
			10'd226 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 16 -> 24
			// srcs: (611, 208)(2928) 5 --> (2928) 5:PUNB, pass, NI0
			10'd227 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 48 -> 25
			// srcs: (612, 209)(2151) 0 --> (2151) 0:PUGB6, pass, PENB
			10'd228 : rdata = 48'b110001110000110100000000000000000000000100000000;
			// PEs: 25 -> 0
			// srcs: (613, 262)(2832) 0 --> (2832) 0:PEGB1, pass, PUGB0
			10'd229 : rdata = 48'b110001110000001000000000000000000000000000001000;
			// PEs: 30 -> 32
			// srcs: (621, 265)(2863) 0 --> (2863) 0:PEGB6, pass, PUNB
			10'd230 : rdata = 48'b110001110000110000000000000000000000001000000000;
			// PEs: 25 -> 8
			// srcs: (622, 264)(2849) -1 --> (2849) -1:PEGB1, pass, PUGB1
			10'd231 : rdata = 48'b110001110000001000000000000000000000000000001001;
			// PEs: 26 -> 32
			// srcs: (623, 267)(2945) 11 --> (2945) 11:PEGB2, pass, PUNB
			10'd232 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 24 -> 25
			// srcs: (630, 210)(2928) 5 --> (2928) 5:NI0, pass, PENB
			10'd233 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 56 -> 24
			// srcs: (631, 213)(2983) -1 --> (2983) -1:PUGB7, pass, NI0
			10'd234 : rdata = 48'b110001110000111100000000000100000000000000000000;
			// PEs: 8 -> 25
			// srcs: (632, 214)(2206) -2 --> (2206) -2:PUGB1, pass, PENB
			10'd235 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 25 -> 56
			// srcs: (637, 266)(2929) 5 --> (2929) 5:PEGB1, pass, PUGB7
			10'd236 : rdata = 48'b110001110000001000000000000000000000000000001111;
			// PEs: 24 -> 25
			// srcs: (638, 215)(2983) -1 --> (2983) -1:NI0, pass, PENB
			10'd237 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 25 -> 16
			// srcs: (645, 271)(2984) -3 --> (2984) -3:PEGB1, pass, PUGB2
			10'd238 : rdata = 48'b110001110000001000000000000000000000000000001010;
			// PEs: 16 -> 25
			// srcs: (664, 216)(3022) -2 --> (3022) -2:PUNB, pass, PENB
			10'd239 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 48 -> 24
			// srcs: (665, 219)(3059) -4 --> (3059) -4:PUGB6, pass, NI0
			10'd240 : rdata = 48'b110001110000110100000000000100000000000000000000;
			// PEs: 32 -> 25
			// srcs: (666, 220)(2283) -6 --> (2283) -6:PUGB4, pass, PENB
			10'd241 : rdata = 48'b110001110000100100000000000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (672, 221)(3059) -4 --> (3059) -4:NI0, pass, PENB
			10'd242 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 0 -> 24
			// srcs: (673, 222)(3080) 0 --> (3080) 0:PUGB0, pass, NI0
			10'd243 : rdata = 48'b110001110000000100000000000100000000000000000000;
			// PEs: 40 -> 25
			// srcs: (674, 223)(2304) 1 --> (2304) 1:PUGB5, pass, PENB
			10'd244 : rdata = 48'b110001110000101100000000000000000000000100000000;
			// PEs: 25 -> 56
			// srcs: (679, 273)(3060) -10 --> (3060) -10:PEGB1, pass, PUGB7
			10'd245 : rdata = 48'b110001110000001000000000000000000000000000001111;
			// PEs: 24 -> 25
			// srcs: (680, 224)(3080) 0 --> (3080) 0:NI0, pass, PENB
			10'd246 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 48 -> 25
			// srcs: (681, 227)(2335) -2 --> (2335) -2:PUGB6, pass, PENB
			10'd247 : rdata = 48'b110001110000110100000000000000000000000100000000;
			// PEs: 32 -> 24
			// srcs: (682, 229)(3123) 7 --> (3123) 7:PUGB4, pass, NI0
			10'd248 : rdata = 48'b110001110000100100000000000100000000000000000000;
			// PEs: 56 -> 25
			// srcs: (683, 230)(2347) 2 --> (2347) 2:PUGB7, pass, PENB
			10'd249 : rdata = 48'b110001110000111100000000000000000000000100000000;
			// PEs: 25 -> 40
			// srcs: (687, 277)(3081) 1 --> (3081) 1:PEGB1, pass, PUGB5
			10'd250 : rdata = 48'b110001110000001000000000000000000000000000001101;
			// PEs: 24 -> 25
			// srcs: (694, 231)(3123) 7 --> (3123) 7:NI0, pass, PENB
			10'd251 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 56 -> 24
			// srcs: (695, 233)(2407) -2 --> (2407) -2:PUGB7, pass, NI0
			10'd252 : rdata = 48'b110001110000111100000000000100000000000000000000;
			// PEs: 16 -> 25
			// srcs: (696, 234)(2409) 8 --> (2409) 8:PUNB, pass, PENB
			10'd253 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 25 -> 0
			// srcs: (697, 278)(3113) -6 --> (3113) -6:PEGB1, pass, PUGB0
			10'd254 : rdata = 48'b110001110000001000000000000000000000000000001000;
			// PEs: 25 -> 32
			// srcs: (701, 279)(3124) 9 --> (3124) 9:PEGB1, pass, PUNB
			10'd255 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 24 -> 25
			// srcs: (702, 235)(2407) -2 --> (2407) -2:NI0, pass, PENB
			10'd256 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 8 -> 25
			// srcs: (703, 237)(2432) 7 --> (2432) 7:PUGB1, pass, PENB
			10'd257 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 16 -> 25
			// srcs: (704, 238)(2458) -2 --> (2458) -2:PUNB, pass, PENB
			10'd258 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 40 -> 24
			// srcs: (705, 240)(2490) 2 --> (2490) 2:PUGB5, pass, NI0
			10'd259 : rdata = 48'b110001110000101100000000000100000000000000000000;
			// PEs: 56 -> 25
			// srcs: (706, 241)(2492) -8 --> (2492) -8:PUGB7, pass, PENB
			10'd260 : rdata = 48'b110001110000111100000000000000000000000100000000;
			// PEs: 25 -> 32
			// srcs: (709, 283)(2410) 6 --> (2410) 6:PEGB1, pass, PUNB
			10'd261 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 25 -> 32
			// srcs: (710, 284)(2433) 3 --> (2433) 3:PEGB1, pass, PUNB
			10'd262 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 24 -> 25
			// srcs: (712, 242)(2490) 2 --> (2490) 2:NI0, pass, PENB
			10'd263 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 16 -> 25
			// srcs: (713, 245)(2538) -2 --> (2538) -2:PUNB, pass, PENB
			10'd264 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 8 -> 24
			// srcs: (714, 246)(2602) 13 --> (2602) 13:PUGB1, pass, NI0
			10'd265 : rdata = 48'b110001110000001100000000000100000000000000000000;
			// PEs: 56 -> 25
			// srcs: (715, 247)(2604) 3 --> (2604) 3:PUGB7, pass, PENB
			10'd266 : rdata = 48'b110001110000111100000000000000000000000100000000;
			// PEs: 25 -> 0
			// srcs: (719, 286)(2493) -6 --> (2493) -6:PEGB1, pass, PUGB0
			10'd267 : rdata = 48'b110001110000001000000000000000000000000000001000;
			// PEs: 25 -> 48
			// srcs: (720, 290)(2541) -7 --> (2541) -7:PEGB1, pass, PUGB6
			10'd268 : rdata = 48'b110001110000001000000000000000000000000000001110;
			// PEs: 24 -> 25
			// srcs: (721, 248)(2602) 13 --> (2602) 13:NI0, pass, PENB
			10'd269 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 32 -> 24
			// srcs: (722, 252)(2662) 0 --> (2662) 0:PUGB4, pass, NI0
			10'd270 : rdata = 48'b110001110000100100000000000100000000000000000000;
			// PEs: 0 -> 25
			// srcs: (723, 253)(2664) -4 --> (2664) -4:PUGB0, pass, PENB
			10'd271 : rdata = 48'b110001110000000100000000000000000000000100000000;
			// PEs: 25 -> 32
			// srcs: (728, 291)(2605) 16 --> (2605) 16:PEGB1, pass, PUNB
			10'd272 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 24 -> 25
			// srcs: (729, 254)(2662) 0 --> (2662) 0:NI0, pass, PENB
			10'd273 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 8 -> 24
			// srcs: (730, 258)(2778) -3 --> (2778) -3:PUGB1, pass, NI0
			10'd274 : rdata = 48'b110001110000001100000000000100000000000000000000;
			// PEs: 56 -> 25
			// srcs: (731, 259)(2780) 8 --> (2780) 8:PUGB7, pass, PENB
			10'd275 : rdata = 48'b110001110000111100000000000000000000000100000000;
			// PEs: 25 -> 0
			// srcs: (736, 292)(2665) -4 --> (2665) -4:PEGB1, pass, PUGB0
			10'd276 : rdata = 48'b110001110000001000000000000000000000000000001000;
			// PEs: 24 -> 25
			// srcs: (737, 260)(2778) -3 --> (2778) -3:NI0, pass, PENB
			10'd277 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 16 -> 25
			// srcs: (738, 263)(2837) 0 --> (2837) 0:PUNB, pass, PENB
			10'd278 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 32 -> 24
			// srcs: (739, 268)(2961) -1 --> (2961) -1:PUGB4, pass, NI0
			10'd279 : rdata = 48'b110001110000100100000000000100000000000000000000;
			// PEs: 56 -> 25
			// srcs: (740, 269)(2963) -7 --> (2963) -7:PUGB7, pass, PENB
			10'd280 : rdata = 48'b110001110000111100000000000000000000000100000000;
			// PEs: 26 -> 0
			// srcs: (741, 298)(2855) 13 --> (2855) 13:PEGB2, pass, PUGB0
			10'd281 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 25 -> 32
			// srcs: (744, 293)(2781) 5 --> (2781) 5:PEGB1, pass, PUNB
			10'd282 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 25 -> 56
			// srcs: (745, 297)(2840) -8 --> (2840) -8:PEGB1, pass, PUGB7
			10'd283 : rdata = 48'b110001110000001000000000000000000000000000001111;
			// PEs: 24 -> 25
			// srcs: (746, 270)(2961) -1 --> (2961) -1:NI0, pass, PENB
			10'd284 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 32 -> 24
			// srcs: (747, 274)(3076) 4 --> (3076) 4:PUGB4, pass, NI0
			10'd285 : rdata = 48'b110001110000100100000000000100000000000000000000;
			// PEs: 0 -> 25
			// srcs: (748, 275)(3078) -2 --> (3078) -2:PUGB0, pass, PENB
			10'd286 : rdata = 48'b110001110000000100000000000000000000000100000000;
			// PEs: 27 -> 32
			// srcs: (749, 299)(2861) 3 --> (2861) 3:PEGB3, pass, PUNB
			10'd287 : rdata = 48'b110001110000011000000000000000000000001000000000;
			// PEs: 25 -> 16
			// srcs: (753, 303)(2964) -8 --> (2964) -8:PEGB1, pass, PUGB2
			10'd288 : rdata = 48'b110001110000001000000000000000000000000000001010;
			// PEs: 24 -> 25
			// srcs: (754, 276)(3076) 4 --> (3076) 4:NI0, pass, PENB
			10'd289 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 8 -> 24
			// srcs: (755, 280)(3129) 9 --> (3129) 9:PUGB1, pass, NI0
			10'd290 : rdata = 48'b110001110000001100000000000100000000000000000000;
			// PEs: 40 -> 25
			// srcs: (756, 281)(3131) -2 --> (3131) -2:PUGB5, pass, PENB
			10'd291 : rdata = 48'b110001110000101100000000000000000000000100000000;
			// PEs: 25 -> 40
			// srcs: (761, 308)(3079) 2 --> (3079) 2:PEGB1, pass, PUGB5
			10'd292 : rdata = 48'b110001110000001000000000000000000000000000001101;
			// PEs: 24 -> 25
			// srcs: (762, 282)(3129) 9 --> (3129) 9:NI0, pass, PENB
			10'd293 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 56 -> 25
			// srcs: (763, 285)(2464) 0 --> (2464) 0:PUGB7, pass, PENB
			10'd294 : rdata = 48'b110001110000111100000000000000000000000100000000;
			// PEs: 32 -> 24
			// srcs: (764, 287)(2530) -1 --> (2530) -1:PUGB4, pass, NI0
			10'd295 : rdata = 48'b110001110000100100000000000100000000000000000000;
			// PEs: 25 -> 32
			// srcs: (769, 309)(3132) 7 --> (3132) 7:PEGB1, pass, PUNB
			10'd296 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 25 -> 56
			// srcs: (770, 310)(2465) 1 --> (2465) 1:PEGB1, pass, PUGB7
			10'd297 : rdata = 48'b110001110000001000000000000000000000000000001111;
			// PEs: 16 -> 29
			// srcs: (775, 272)(3021) -1 --> (3021) -1:PUNB, pass, PEGB5
			10'd298 : rdata = 48'b110001101111111100000000000000000000000011010000;
			// PEs: 16 -> 25
			// srcs: (776, 288)(2535) -8 --> (2535) -8:PUNB, pass, PENB
			10'd299 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (782, 289)(2530) -1 --> (2530) -1:NI0, pass, PENB
			10'd300 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 16 -> 24
			// srcs: (783, 294)(2801) 4 --> (2801) 4:PUNB, pass, NI0
			10'd301 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 48 -> 25
			// srcs: (784, 295)(2806) 2 --> (2806) 2:PUGB6, pass, PENB
			10'd302 : rdata = 48'b110001110000110100000000000000000000000100000000;
			// PEs: 16 -> 28
			// srcs: (785, 304)(3019) -11 --> (3019) -11:PUNB, pass, PEGB4
			10'd303 : rdata = 48'b110001101111111100000000000000000000000011000000;
			// PEs: 25 -> 0
			// srcs: (789, 314)(2536) -9 --> (2536) -9:PEGB1, pass, PUGB0
			10'd304 : rdata = 48'b110001110000001000000000000000000000000000001000;
			// PEs: 24 -> 25
			// srcs: (790, 296)(2801) 4 --> (2801) 4:NI0, pass, PENB
			10'd305 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 48 -> 24
			// srcs: (791, 300)(2921) -1 --> (2921) -1:PUGB6, pass, NI0
			10'd306 : rdata = 48'b110001110000110100000000000100000000000000000000;
			// PEs: 32 -> 25
			// srcs: (792, 301)(2926) -2 --> (2926) -2:PUGB4, pass, PENB
			10'd307 : rdata = 48'b110001110000100100000000000000000000000100000000;
			// PEs: 25 -> 8
			// srcs: (797, 315)(2807) 6 --> (2807) 6:PEGB1, pass, PUGB1
			10'd308 : rdata = 48'b110001110000001000000000000000000000000000001001;
			// PEs: 24 -> 25
			// srcs: (798, 302)(2921) -1 --> (2921) -1:NI0, pass, PENB
			10'd309 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 40 -> 24
			// srcs: (799, 305)(3056) -4 --> (3056) -4:PUGB5, pass, NI0
			10'd310 : rdata = 48'b110001110000101100000000000100000000000000000000;
			// PEs: 56 -> 25
			// srcs: (800, 306)(3061) -15 --> (3061) -15:PUGB7, pass, PENB
			10'd311 : rdata = 48'b110001110000111100000000000000000000000100000000;
			// PEs: 25 -> 56
			// srcs: (805, 319)(2927) -3 --> (2927) -3:PEGB1, pass, PUGB7
			10'd312 : rdata = 48'b110001110000001000000000000000000000000000001111;
			// PEs: 24 -> 25
			// srcs: (806, 307)(3056) -4 --> (3056) -4:NI0, pass, PENB
			10'd313 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 16 -> 24
			// srcs: (807, 311)(2513) 16 --> (2513) 16:PUNB, pass, NI0
			10'd314 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 40 -> 25
			// srcs: (808, 312)(2524) 3 --> (2524) 3:PUGB5, pass, PENB
			10'd315 : rdata = 48'b110001110000101100000000000000000000000100000000;
			// PEs: 31 -> 16
			// srcs: (809, 326)(3037) -9 --> (3037) -9:PENB, pass, PUGB2
			10'd316 : rdata = 48'b110001101111111000000000000000000000000000001010;
			// PEs: 25 -> 56
			// srcs: (813, 320)(3062) -19 --> (3062) -19:PEGB1, pass, PUGB7
			10'd317 : rdata = 48'b110001110000001000000000000000000000000000001111;
			// PEs: 24 -> 25
			// srcs: (814, 313)(2513) 16 --> (2513) 16:NI0, pass, PENB
			10'd318 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 40 -> 24
			// srcs: (815, 316)(2830) 1 --> (2830) 1:PUGB5, pass, NI0
			10'd319 : rdata = 48'b110001110000101100000000000100000000000000000000;
			// PEs: 25 -> 32
			// srcs: (821, 324)(2525) 19 --> (2525) 19:PEGB1, pass, PUNB
			10'd320 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 56 -> 25
			// srcs: (1167, 317)(2841) -14 --> (2841) -14:PUGB7, pass, PENB
			10'd321 : rdata = 48'b110001110000111100000000000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (1174, 318)(2830) 1 --> (2830) 1:NI0, pass, PENB
			10'd322 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 16 -> 24
			// srcs: (1175, 321)(2380) -18 --> (2380) -18:PUNB, pass, NI0
			10'd323 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 32 -> 25
			// srcs: (1176, 322)(2403) -6 --> (2403) -6:PUGB4, pass, PENB
			10'd324 : rdata = 48'b110001110000100100000000000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (1182, 323)(2380) -18 --> (2380) -18:NI0, pass, PENB
			10'd325 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 8 -> 25
			// srcs: (1416, 325)(2819) 3 --> (2819) 3:PUGB1, pass, PENB
			10'd326 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 48 -> 25
			// srcs: (1417, 327)(2452) 14 --> (2452) 14:PUGB6, pass, PENB
			10'd327 : rdata = 48'b110001110000110100000000000000000000000100000000;
			// PEs: 25 -> 16
			// srcs: (1424, 328)(2843) -10 --> (2843) -10:PEGB1, pass, PUGB2
			10'd328 : rdata = 48'b110001110000001000000000000000000000000000001010;
			// PEs: 25 -> 0
			// srcs: (1425, 332)(2453) -10 --> (2453) -10:PEGB1, pass, PUGB0
			10'd329 : rdata = 48'b110001110000001000000000000000000000000000001000;
			// PEs: 48 -> 24
			// srcs: (1426, 329)(2892) 28 --> (2892) 28:PUGB6, pass, NI0
			10'd330 : rdata = 48'b110001110000110100000000000100000000000000000000;
			// PEs: 32 -> 25
			// srcs: (1427, 330)(2940) 27 --> (2940) 27:PUGB4, pass, PENB
			10'd331 : rdata = 48'b110001110000100100000000000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (1433, 331)(2892) 28 --> (2892) 28:NI0, pass, PENB
			10'd332 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 16 -> 25
			// srcs: (1445, 333)(2844) -31 --> (2844) -31:PUNB, pass, PENB
			10'd333 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 25 -> 48
			// srcs: (1453, 334)(2942) 24 --> (2942) 24:PEGB1, pass, PUGB6
			10'd334 : rdata = 48'b110001110000001000000000000000000000000000001110;
			// PEs: 8 -> 25
			// srcs: (1538, 335)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd335 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 26
			// srcs: (1540, 336)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd336 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 27
			// srcs: (1541, 337)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd337 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 28
			// srcs: (1543, 338)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd338 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 29
			// srcs: (1544, 339)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd339 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 30
			// srcs: (1546, 340)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd340 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 31
			// srcs: (1547, 341)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd341 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 25
			// srcs: (1618, 342)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd342 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 26
			// srcs: (1620, 343)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd343 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 27
			// srcs: (1621, 344)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd344 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 28
			// srcs: (1623, 345)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd345 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 29
			// srcs: (1624, 346)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd346 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 30
			// srcs: (1626, 347)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd347 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 31
			// srcs: (1627, 348)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd348 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 25
			// srcs: (1634, 349)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd349 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 26
			// srcs: (1637, 350)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd350 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 27
			// srcs: (1640, 351)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd351 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 28
			// srcs: (1643, 352)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd352 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 29
			// srcs: (1646, 353)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd353 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 30
			// srcs: (1649, 354)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd354 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 31
			// srcs: (1652, 355)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd355 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 25
			// srcs: (1700, 356)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd356 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 26
			// srcs: (1702, 357)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd357 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 27
			// srcs: (1703, 358)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd358 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 28
			// srcs: (1705, 359)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd359 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 29
			// srcs: (1706, 360)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd360 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 30
			// srcs: (1707, 361)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd361 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 31
			// srcs: (1708, 362)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd362 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 25
			// srcs: (1780, 363)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd363 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 26
			// srcs: (1782, 364)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd364 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 27
			// srcs: (1783, 365)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd365 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 28
			// srcs: (1785, 366)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd366 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 29
			// srcs: (1786, 367)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd367 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 30
			// srcs: (1788, 368)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd368 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 31
			// srcs: (1789, 369)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd369 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 25
			// srcs: (1818, 370)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd370 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 26
			// srcs: (1821, 371)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd371 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 27
			// srcs: (1824, 372)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd372 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 28
			// srcs: (1827, 373)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd373 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 29
			// srcs: (1830, 374)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd374 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 30
			// srcs: (1833, 375)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd375 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 31
			// srcs: (1836, 376)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd376 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 25
			// srcs: (1860, 377)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd377 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 26
			// srcs: (1862, 378)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd378 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 27
			// srcs: (1863, 379)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd379 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 28
			// srcs: (1865, 380)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd380 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 29
			// srcs: (1866, 381)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd381 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 30
			// srcs: (1868, 382)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd382 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 31
			// srcs: (1869, 383)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd383 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 25
			// srcs: (1942, 384)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd384 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 26
			// srcs: (1944, 385)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd385 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 27
			// srcs: (1945, 386)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd386 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 28
			// srcs: (1947, 387)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd387 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 29
			// srcs: (1948, 388)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd388 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 30
			// srcs: (1950, 389)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd389 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 31
			// srcs: (1951, 390)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd390 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 25
			// srcs: (1998, 391)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd391 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 26
			// srcs: (2005, 392)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd392 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 27
			// srcs: (2008, 393)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd393 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 28
			// srcs: (2011, 394)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd394 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 29
			// srcs: (2014, 395)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd395 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 30
			// srcs: (2017, 396)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd396 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 31
			// srcs: (2020, 397)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd397 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 25
			// srcs: (2022, 398)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd398 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 26
			// srcs: (2024, 399)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd399 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 27
			// srcs: (2025, 400)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd400 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 28
			// srcs: (2027, 401)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd401 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 29
			// srcs: (2028, 402)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd402 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 30
			// srcs: (2030, 403)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd403 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 31
			// srcs: (2031, 404)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd404 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 25
			// srcs: (2102, 405)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd405 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 26
			// srcs: (2104, 406)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd406 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 27
			// srcs: (2105, 407)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd407 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 28
			// srcs: (2107, 408)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd408 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 29
			// srcs: (2108, 409)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd409 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 30
			// srcs: (2110, 410)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd410 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 31
			// srcs: (2111, 411)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd411 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 25
			// srcs: (2182, 412)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd412 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 25
			// srcs: (2184, 413)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd413 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 26
			// srcs: (2185, 414)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd414 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 26
			// srcs: (2186, 415)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd415 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 27
			// srcs: (2187, 416)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd416 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 27
			// srcs: (2188, 417)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd417 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 28
			// srcs: (2189, 418)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd418 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 29
			// srcs: (2190, 419)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd419 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 28
			// srcs: (2191, 420)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd420 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 30
			// srcs: (2192, 421)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd421 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 31
			// srcs: (2193, 422)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd422 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 29
			// srcs: (2194, 423)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd423 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 30
			// srcs: (2201, 424)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd424 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 31
			// srcs: (2204, 425)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd425 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 25
			// srcs: (2264, 426)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd426 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 26
			// srcs: (2266, 427)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd427 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 27
			// srcs: (2267, 428)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd428 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 28
			// srcs: (2269, 429)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd429 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 29
			// srcs: (2270, 430)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd430 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 30
			// srcs: (2272, 431)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd431 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 31
			// srcs: (2273, 432)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd432 : rdata = 48'b110001110000001100000000000000000000000011110000;
			default : rdata = 48'b000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 25) begin
	always @(*) begin
		case(address)
			// PEs: 25, 25 -> 24
			// srcs: (1, 0)(33) 2, (818) -2 --> (1602) -4:ND0, NW0, *, PEGB0
			10'd0 : rdata = 48'b000110110000000001000000000000000000000010000000;
			// PEs: 25, 25 -> 24
			// srcs: (2, 1)(113) -2, (898) 1 --> (1682) -2:ND1, NW1, *, PEGB0
			10'd1 : rdata = 48'b000110110000000101000000001000000000000010000000;
			// PEs: 25, 25 -> 24
			// srcs: (3, 2)(195) 2, (980) 0 --> (1764) 0:ND2, NW2, *, PEGB0
			10'd2 : rdata = 48'b000110110000001001000000010000000000000010000000;
			// PEs: 25, 25 -> 24
			// srcs: (4, 3)(275) -3, (1060) -3 --> (1844) 9:ND3, NW3, *, PEGB0
			10'd3 : rdata = 48'b000110110000001101000000011000000000000010000000;
			// PEs: 25, 25 -> 31
			// srcs: (5, 4)(355) -2, (1140) 1 --> (1924) -2:ND4, NW4, *, PEGB7
			10'd4 : rdata = 48'b000110110000010001000000100000000000000011110000;
			// PEs: 25, 25 -> 26
			// srcs: (6, 5)(437) -3, (1222) -1 --> (2006) 3:ND5, NW5, *, PENB
			10'd5 : rdata = 48'b000110110000010101000000101000000000000100000000;
			// PEs: 25, 25 -> 27
			// srcs: (7, 6)(517) -1, (1302) -3 --> (2086) 3:ND6, NW6, *, PEGB3
			10'd6 : rdata = 48'b000110110000011001000000110000000000000010110000;
			// PEs: 25, 25 -> 25
			// srcs: (8, 7)(597) 0, (1382) -3 --> (2166) 0:ND7, NW7, *, NI0
			10'd7 : rdata = 48'b000110110000011101000000111100000000000000000000;
			// PEs: 25, 25 -> 25
			// srcs: (9, 8)(679) 1, (1464) 0 --> (2248) 0:ND8, NW8, *, NI1
			10'd8 : rdata = 48'b000110110000100001000001000100001000000000000000;
			// PEs: 25, 25 -> 25
			// srcs: (10, 9)(759) -1, (1544) 1 --> (2328) -1:ND9, NW9, *, NI2
			10'd9 : rdata = 48'b000110110000100101000001001100010000000000000000;
			// PEs: 25, 25 -> 25
			// srcs: (11, 10)(129) 2, (914) -2 --> (1698) -4:ND10, NW10, *, NI3
			10'd10 : rdata = 48'b000110110000101001000001010100011000000000000000;
			// PEs: 25, 25 -> 25
			// srcs: (12, 11)(313) -3, (1098) 0 --> (1882) 0:ND11, NW11, *, NI4
			10'd11 : rdata = 48'b000110110000101101000001011100100000000000000000;
			// PEs: 25, 25 -> 25
			// srcs: (13, 12)(493) 0, (1278) 0 --> (2062) 0:ND12, NW12, *, NI5
			10'd12 : rdata = 48'b000110110000110001000001100100101000000000000000;
			// PEs: 25, 25 -> 25
			// srcs: (14, 13)(677) -1, (1462) -1 --> (2246) 1:ND13, NW13, *, NI6
			10'd13 : rdata = 48'b000110110000110101000001101100110000000000000000;
			// PEs: 24 -> 
			// srcs: (32, 14)(1657) 1 --> (1657) 1:PENB, pass, 
			10'd14 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 24, 25 -> 24
			// srcs: (38, 15)(1656) 0, (1657) 1 --> (2436) 1:PENB, ALU, +, PEGB0
			10'd15 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 24 -> 
			// srcs: (51, 16)(1792) 0 --> (1792) 0:PENB, pass, 
			10'd16 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 24, 25 -> 24
			// srcs: (58, 17)(1791) 0, (1792) 0 --> (2571) 0:PENB, ALU, +, PEGB0
			10'd17 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 24 -> 
			// srcs: (75, 18)(1921) -6 --> (1921) -6:PENB, pass, 
			10'd18 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 24, 25 -> 25
			// srcs: (81, 19)(1920) 6, (1921) -6 --> (2700) 0:PENB, ALU, +, NI7
			10'd19 : rdata = 48'b000011101111111000111111111100111000000000000000;
			// PEs: 24 -> 
			// srcs: (87, 20)(1997) -6 --> (1997) -6:PENB, pass, 
			10'd20 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 24, 25 -> 24
			// srcs: (93, 21)(1996) 3, (1997) -6 --> (2777) -3:PENB, ALU, +, PEGB0
			10'd21 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 24 -> 
			// srcs: (95, 22)(2000) 6 --> (2000) 6:PENB, pass, 
			10'd22 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 24, 25 -> 24
			// srcs: (101, 23)(1999) 2, (2000) 6 --> (2779) 8:PENB, ALU, +, PEGB0
			10'd23 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 24 -> 
			// srcs: (103, 24)(2003) 2 --> (2003) 2:PENB, pass, 
			10'd24 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 24, 25 -> 24
			// srcs: (109, 25)(2002) -4, (2003) 2 --> (2783) -2:PENB, ALU, +, PEGB0
			10'd25 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 24 -> 
			// srcs: (111, 26)(2077) 1 --> (2077) 1:PENB, pass, 
			10'd26 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 24, 25 -> 27
			// srcs: (117, 27)(2076) 0, (2077) 1 --> (2857) 1:PENB, ALU, +, PEGB3
			10'd27 : rdata = 48'b000011101111111000111111111000000000000010110000;
			// PEs: 24 -> 
			// srcs: (119, 28)(2080) 0 --> (2080) 0:PENB, pass, 
			10'd28 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 24, 25 -> 30
			// srcs: (125, 29)(2079) 0, (2080) 0 --> (2859) 0:PENB, ALU, +, PEGB6
			10'd29 : rdata = 48'b000011101111111000111111111000000000000011100000;
			// PEs: 24 -> 
			// srcs: (127, 30)(2083) 0 --> (2083) 0:PENB, pass, 
			10'd30 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 24, 25 -> 30
			// srcs: (133, 31)(2082) 2, (2083) 0 --> (2862) 2:PENB, ALU, +, PEGB6
			10'd31 : rdata = 48'b000011101111111000111111111000000000000011100000;
			// PEs: 24 -> 
			// srcs: (135, 32)(2159) -3 --> (2159) -3:PENB, pass, 
			10'd32 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 24, 25 -> 25
			// srcs: (141, 33)(2158) 0, (2159) -3 --> (2935) -3:PENB, ALU, +, NI8
			10'd33 : rdata = 48'b000011101111111000111111111101000000000000000000;
			// PEs: 24, 25 -> 25
			// srcs: (142, 34)(2165) 0, (2166) 0 --> (2946) 0:PENB, NI0, +, NI9
			10'd34 : rdata = 48'b000011101111111010100000000101001000000000000000;
			// PEs: 24, 25 -> 26
			// srcs: (143, 35)(2247) -2, (2248) 0 --> (3026) -2:PENB, NI1, +, PENB
			10'd35 : rdata = 48'b000011101111111010100000001000000000000100000000;
			// PEs: 24, 25 -> 24
			// srcs: (144, 36)(2327) 0, (2328) -1 --> (3105) -1:PENB, NI2, +, PEGB0
			10'd36 : rdata = 48'b000011101111111010100000010000000000000010000000;
			// PEs: 25 -> 24
			// srcs: (152, 52)(1698) -4 --> (1698) -4:NI3, pass, PEGB0
			10'd37 : rdata = 48'b110001010000001100000000000000000000000010000000;
			// PEs: 25 -> 24
			// srcs: (160, 64)(1882) 0 --> (1882) 0:NI4, pass, PEGB0
			10'd38 : rdata = 48'b110001010000010000000000000000000000000010000000;
			// PEs: 25 -> 24
			// srcs: (162, 81)(2935) -3 --> (2935) -3:NI8, pass, PEGB0
			10'd39 : rdata = 48'b110001010000100000000000000000000000000010000000;
			// PEs: 25 -> 24
			// srcs: (168, 66)(2700) 0 --> (2700) 0:NI7, pass, PEGB0
			10'd40 : rdata = 48'b110001010000011100000000000000000000000010000000;
			// PEs: 25 -> 24
			// srcs: (182, 83)(2946) 0 --> (2946) 0:NI9, pass, PEGB0
			10'd41 : rdata = 48'b110001010000100100000000000000000000000010000000;
			// PEs: 24 -> 
			// srcs: (274, 37)(1917) 0 --> (1917) 0:PENB, pass, 
			10'd42 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 24, 25 -> 25
			// srcs: (280, 38)(1916) 2, (1917) 0 --> (2697) 2:PENB, ALU, +, NI0
			10'd43 : rdata = 48'b000011101111111000111111111100000000000000000000;
			// PEs: 24 -> 
			// srcs: (306, 39)(1919) 4 --> (1919) 4:PENB, pass, 
			10'd44 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 24, 25 -> 26
			// srcs: (312, 40)(1918) 1, (1919) 4 --> (2698) 5:PENB, ALU, +, PENB
			10'd45 : rdata = 48'b000011101111111000111111111000000000000100000000;
			// PEs: 25 -> 26
			// srcs: (319, 65)(2697) 2 --> (2697) 2:NI0, pass, PENB
			10'd46 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 24 -> 
			// srcs: (335, 41)(2162) 4 --> (2162) 4:PENB, pass, 
			10'd47 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 24, 25 -> 25
			// srcs: (341, 42)(2161) 0, (2162) 4 --> (2943) 4:PENB, ALU, +, NI0
			10'd48 : rdata = 48'b000011101111111000111111111100000000000000000000;
			// PEs: 24 -> 
			// srcs: (343, 43)(2164) 4 --> (2164) 4:PENB, pass, 
			10'd49 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 24, 25 -> 26
			// srcs: (349, 44)(2163) 3, (2164) 4 --> (2944) 7:PENB, ALU, +, PENB
			10'd50 : rdata = 48'b000011101111111000111111111000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (351, 45)(1606) 6 --> (1606) 6:PENB, pass, NI1
			10'd51 : rdata = 48'b110001101111111000000000000100001000000000000000;
			// PEs: 25 -> 26
			// srcs: (356, 82)(2943) 4 --> (2943) 4:NI0, pass, PENB
			10'd52 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 24, 25 -> 24
			// srcs: (357, 46)(2386) -3, (1606) 6 --> (2387) 3:PENB, NI1, +, PEGB0
			10'd53 : rdata = 48'b000011101111111010100000001000000000000010000000;
			// PEs: 26, 24 -> 24
			// srcs: (358, 47)(2417) -1, (1637) 0 --> (2418) -1:PEGB2, PENB, +, PEGB0
			10'd54 : rdata = 48'b000011110000010011011111110000000000000010000000;
			// PEs: 30, 24 -> 25
			// srcs: (359, 48)(2429) -4, (1649) 0 --> (2430) -4:PEGB6, PENB, +, NI0
			10'd55 : rdata = 48'b000011110000110011011111110100000000000000000000;
			// PEs: 24, 27 -> 25
			// srcs: (360, 49)(2454) 3, (2455) 0 --> (2456) 3:PENB, PEGB3, +, NI1
			10'd56 : rdata = 48'b000011101111111011100000110100001000000000000000;
			// PEs: 24 -> 
			// srcs: (524, 50)(1686) -1 --> (1686) -1:PENB, pass, 
			10'd57 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 24, 25 -> 24
			// srcs: (530, 51)(2466) 1, (1686) -1 --> (2467) 0:PENB, ALU, +, PEGB0
			10'd58 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 24 -> 
			// srcs: (532, 53)(1726) 6 --> (1726) 6:PENB, pass, 
			10'd59 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 24, 25 -> 24
			// srcs: (538, 54)(2505) 8, (1726) 6 --> (2506) 14:PENB, ALU, +, PEGB0
			10'd60 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 24 -> 
			// srcs: (540, 55)(1747) 0 --> (1747) 0:PENB, pass, 
			10'd61 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 24, 25 -> 24
			// srcs: (546, 56)(2526) 0, (1747) 0 --> (2527) 0:PENB, ALU, +, PEGB0
			10'd62 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 27, 24 -> 25
			// srcs: (554, 57)(2539) -5, (1762) 0 --> (2540) -5:PEGB3, PENB, +, NI2
			10'd63 : rdata = 48'b000011110000011011011111110100010000000000000000;
			// PEs: 24 -> 
			// srcs: (555, 58)(1833) 0 --> (1833) 0:PENB, pass, 
			10'd64 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 24, 25 -> 24
			// srcs: (560, 59)(2612) 6, (1833) 0 --> (2613) 6:PENB, ALU, +, PEGB0
			10'd65 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 24 -> 
			// srcs: (562, 60)(1845) 0 --> (1845) 0:PENB, pass, 
			10'd66 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 24, 25 -> 24
			// srcs: (568, 61)(2624) 10, (1845) 0 --> (2625) 10:PENB, ALU, +, PEGB0
			10'd67 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 24 -> 
			// srcs: (570, 62)(1863) 6 --> (1863) 6:PENB, pass, 
			10'd68 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 24, 25 -> 24
			// srcs: (576, 63)(2640) 1, (1863) 6 --> (2641) 7:PENB, ALU, +, PEGB0
			10'd69 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 24 -> 
			// srcs: (578, 67)(1980) 0 --> (1980) 0:PENB, pass, 
			10'd70 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 24, 25 -> 24
			// srcs: (584, 68)(2760) 0, (1980) 0 --> (2761) 0:PENB, ALU, +, PEGB0
			10'd71 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 24 -> 
			// srcs: (586, 69)(1992) 4 --> (1992) 4:PENB, pass, 
			10'd72 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 24, 25 -> 24
			// srcs: (592, 70)(2772) -1, (1992) 4 --> (2773) 3:PENB, ALU, +, PEGB0
			10'd73 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 24 -> 
			// srcs: (594, 71)(2041) 2 --> (2041) 2:PENB, pass, 
			10'd74 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 24, 25 -> 24
			// srcs: (600, 72)(2820) 3, (2041) 2 --> (2821) 5:PENB, ALU, +, PEGB0
			10'd75 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 24 -> 
			// srcs: (602, 73)(2053) 4 --> (2053) 4:PENB, pass, 
			10'd76 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 24, 25 -> 24
			// srcs: (608, 74)(2831) -4, (2053) 4 --> (2832) 0:PENB, ALU, +, PEGB0
			10'd77 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 24, 25 -> 25
			// srcs: (609, 75)(2838) -8, (2062) 0 --> (2839) -8:PENB, NI5, +, NI3
			10'd78 : rdata = 48'b000011101111111010100000101100011000000000000000;
			// PEs: 24, 26 -> 24
			// srcs: (617, 76)(2848) -1, (2069) 0 --> (2849) -1:PENB, PEGB2, +, PEGB0
			10'd79 : rdata = 48'b000011101111111011100000100000000000000010000000;
			// PEs: 24, 27 -> 25
			// srcs: (625, 77)(2851) 6, (2072) 2 --> (2852) 8:PENB, PEGB3, +, NI4
			10'd80 : rdata = 48'b000011101111111011100000110100100000000000000000;
			// PEs: 24, 28 -> 26
			// srcs: (626, 78)(2853) 6, (2075) -1 --> (2854) 5:PENB, PEGB4, +, PENB
			10'd81 : rdata = 48'b000011101111111011100001000000000000000100000000;
			// PEs: 24 -> 
			// srcs: (627, 79)(2151) 0 --> (2151) 0:PENB, pass, 
			10'd82 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 24, 25 -> 24
			// srcs: (632, 80)(2928) 5, (2151) 0 --> (2929) 5:PENB, ALU, +, PEGB0
			10'd83 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 25 -> 26
			// srcs: (633, 108)(2852) 8 --> (2852) 8:NI4, pass, PENB
			10'd84 : rdata = 48'b110001010000010000000000000000000000000100000000;
			// PEs: 24 -> 
			// srcs: (634, 84)(2206) -2 --> (2206) -2:PENB, pass, 
			10'd85 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 24, 25 -> 24
			// srcs: (640, 85)(2983) -1, (2206) -2 --> (2984) -3:PENB, ALU, +, PEGB0
			10'd86 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 24, 25 -> 29
			// srcs: (666, 86)(3022) -2, (2246) 1 --> (3023) -1:PENB, NI6, +, PEGB5
			10'd87 : rdata = 48'b000011101111111010100000110000000000000011010000;
			// PEs: 24 -> 
			// srcs: (668, 87)(2283) -6 --> (2283) -6:PENB, pass, 
			10'd88 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 24, 25 -> 24
			// srcs: (674, 88)(3059) -4, (2283) -6 --> (3060) -10:PENB, ALU, +, PEGB0
			10'd89 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 24 -> 
			// srcs: (676, 89)(2304) 1 --> (2304) 1:PENB, pass, 
			10'd90 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 24, 25 -> 24
			// srcs: (682, 90)(3080) 0, (2304) 1 --> (3081) 1:PENB, ALU, +, PEGB0
			10'd91 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 26, 24 -> 24
			// srcs: (690, 91)(3112) -4, (2335) -2 --> (3113) -6:PEGB2, PENB, +, PEGB0
			10'd92 : rdata = 48'b000011110000010011011111110000000000000010000000;
			// PEs: 24 -> 
			// srcs: (691, 92)(2347) 2 --> (2347) 2:PENB, pass, 
			10'd93 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 24, 25 -> 24
			// srcs: (696, 93)(3123) 7, (2347) 2 --> (3124) 9:PENB, ALU, +, PEGB0
			10'd94 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 24 -> 
			// srcs: (698, 94)(2409) 8 --> (2409) 8:PENB, pass, 
			10'd95 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 24, 25 -> 24
			// srcs: (704, 95)(2407) -2, (2409) 8 --> (2410) 6:PENB, ALU, +, PEGB0
			10'd96 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 25, 24 -> 24
			// srcs: (705, 96)(2430) -4, (2432) 7 --> (2433) 3:NI0, PENB, +, PEGB0
			10'd97 : rdata = 48'b000011010000000011011111110000000000000010000000;
			// PEs: 25, 24 -> 25
			// srcs: (706, 97)(2456) 3, (2458) -2 --> (2459) 1:NI1, PENB, +, NI0
			10'd98 : rdata = 48'b000011010000000111011111110100000000000000000000;
			// PEs: 24 -> 
			// srcs: (708, 98)(2492) -8 --> (2492) -8:PENB, pass, 
			10'd99 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 24, 25 -> 24
			// srcs: (714, 99)(2490) 2, (2492) -8 --> (2493) -6:PENB, ALU, +, PEGB0
			10'd100 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 24, 25 -> 24
			// srcs: (715, 100)(2538) -2, (2540) -5 --> (2541) -7:PENB, NI2, +, PEGB0
			10'd101 : rdata = 48'b000011101111111010100000010000000000000010000000;
			// PEs: 24 -> 
			// srcs: (717, 101)(2604) 3 --> (2604) 3:PENB, pass, 
			10'd102 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 24, 25 -> 24
			// srcs: (723, 102)(2602) 13, (2604) 3 --> (2605) 16:PENB, ALU, +, PEGB0
			10'd103 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 24 -> 
			// srcs: (725, 103)(2664) -4 --> (2664) -4:PENB, pass, 
			10'd104 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 24, 25 -> 24
			// srcs: (731, 104)(2662) 0, (2664) -4 --> (2665) -4:PENB, ALU, +, PEGB0
			10'd105 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 24 -> 
			// srcs: (733, 105)(2780) 8 --> (2780) 8:PENB, pass, 
			10'd106 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 24, 25 -> 24
			// srcs: (739, 106)(2778) -3, (2780) 8 --> (2781) 5:PENB, ALU, +, PEGB0
			10'd107 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 24, 25 -> 24
			// srcs: (740, 107)(2837) 0, (2839) -8 --> (2840) -8:PENB, NI3, +, PEGB0
			10'd108 : rdata = 48'b000011101111111010100000011000000000000010000000;
			// PEs: 24 -> 
			// srcs: (742, 109)(2963) -7 --> (2963) -7:PENB, pass, 
			10'd109 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 24, 25 -> 24
			// srcs: (748, 110)(2961) -1, (2963) -7 --> (2964) -8:PENB, ALU, +, PEGB0
			10'd110 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 24 -> 
			// srcs: (750, 111)(3078) -2 --> (3078) -2:PENB, pass, 
			10'd111 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 24, 25 -> 24
			// srcs: (756, 112)(3076) 4, (3078) -2 --> (3079) 2:PENB, ALU, +, PEGB0
			10'd112 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 24 -> 
			// srcs: (758, 113)(3131) -2 --> (3131) -2:PENB, pass, 
			10'd113 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 24, 25 -> 24
			// srcs: (764, 114)(3129) 9, (3131) -2 --> (3132) 7:PENB, ALU, +, PEGB0
			10'd114 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 25, 24 -> 24
			// srcs: (765, 115)(2459) 1, (2464) 0 --> (2465) 1:NI0, PENB, +, PEGB0
			10'd115 : rdata = 48'b000011010000000011011111110000000000000010000000;
			// PEs: 24 -> 
			// srcs: (778, 116)(2535) -8 --> (2535) -8:PENB, pass, 
			10'd116 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 24, 25 -> 24
			// srcs: (784, 117)(2530) -1, (2535) -8 --> (2536) -9:PENB, ALU, +, PEGB0
			10'd117 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 24 -> 
			// srcs: (786, 118)(2806) 2 --> (2806) 2:PENB, pass, 
			10'd118 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 24, 25 -> 24
			// srcs: (792, 119)(2801) 4, (2806) 2 --> (2807) 6:PENB, ALU, +, PEGB0
			10'd119 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 24 -> 
			// srcs: (794, 120)(2926) -2 --> (2926) -2:PENB, pass, 
			10'd120 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 24, 25 -> 24
			// srcs: (800, 121)(2921) -1, (2926) -2 --> (2927) -3:PENB, ALU, +, PEGB0
			10'd121 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 24 -> 
			// srcs: (802, 122)(3061) -15 --> (3061) -15:PENB, pass, 
			10'd122 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 24, 25 -> 24
			// srcs: (808, 123)(3056) -4, (3061) -15 --> (3062) -19:PENB, ALU, +, PEGB0
			10'd123 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 24 -> 
			// srcs: (810, 124)(2524) 3 --> (2524) 3:PENB, pass, 
			10'd124 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 24, 25 -> 24
			// srcs: (816, 125)(2513) 16, (2524) 3 --> (2525) 19:PENB, ALU, +, PEGB0
			10'd125 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 24 -> 
			// srcs: (1169, 126)(2841) -14 --> (2841) -14:PENB, pass, 
			10'd126 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 24, 25 -> 25
			// srcs: (1176, 127)(2830) 1, (2841) -14 --> (2842) -13:PENB, ALU, +, NI0
			10'd127 : rdata = 48'b000011101111111000111111111100000000000000000000;
			// PEs: 24 -> 
			// srcs: (1178, 128)(2403) -6 --> (2403) -6:PENB, pass, 
			10'd128 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 24, 25 -> 25
			// srcs: (1184, 129)(2380) -18, (2403) -6 --> (2404) -24:PENB, ALU, +, NI1
			10'd129 : rdata = 48'b000011101111111000111111111100001000000000000000;
			// PEs: 24, 25 -> 24
			// srcs: (1419, 130)(2819) 3, (2842) -13 --> (2843) -10:PENB, NI0, +, PEGB0
			10'd130 : rdata = 48'b000011101111111010100000000000000000000010000000;
			// PEs: 25, 24 -> 24
			// srcs: (1420, 131)(2404) -24, (2452) 14 --> (2453) -10:NI1, PENB, +, PEGB0
			10'd131 : rdata = 48'b000011010000000111011111110000000000000010000000;
			// PEs: 24 -> 
			// srcs: (1429, 132)(2940) 27 --> (2940) 27:PENB, pass, 
			10'd132 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 24, 25 -> 
			// srcs: (1435, 133)(2892) 28, (2940) 27 --> (2941) 55:PENB, ALU, +, 
			10'd133 : rdata = 48'b000011101111111000111111111000000000000000000000;
			// PEs: 24, 25 -> 24
			// srcs: (1448, 134)(2844) -31, (2941) 55 --> (2942) 24:PENB, ALU, +, PEGB0
			10'd134 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 24, 25 -> 26
			// srcs: (1540, 135)(3140) 47, (33) 2 --> (3170) 94:PENB, ND0, *, PENB
			10'd135 : rdata = 48'b000111101111111001100000000000000000000100000000;
			// PEs: 25, 26 -> 25
			// srcs: (1549, 149)(818) -2, (3954) 94 --> (4738) -96:NW0, PEGB2, -, NW0
			10'd136 : rdata = 48'b000100100000000011100000100000000100000000000000;
			// PEs: 24, 25 -> 26
			// srcs: (1620, 136)(3140) 47, (113) -2 --> (3250) -94:PENB, ND1, *, PENB
			10'd137 : rdata = 48'b000111101111111001100000001000000000000100000000;
			// PEs: 25, 26 -> 25
			// srcs: (1629, 150)(898) 1, (4034) -94 --> (4818) 95:NW1, PEGB2, -, NW1
			10'd138 : rdata = 48'b000100100000000111100000100000000100010000000000;
			// PEs: 24, 25 -> 26
			// srcs: (1636, 137)(3140) 47, (129) 2 --> (3266) 94:PENB, ND10, *, PENB
			10'd139 : rdata = 48'b000111101111111001100001010000000000000100000000;
			// PEs: 25, 26 -> 25
			// srcs: (1645, 151)(914) -2, (4050) 94 --> (4834) -96:NW10, PEGB2, -, NW10
			10'd140 : rdata = 48'b000100100000101011100000100000000110100000000000;
			// PEs: 24, 25 -> 26
			// srcs: (1702, 138)(3140) 47, (195) 2 --> (3332) 94:PENB, ND2, *, PENB
			10'd141 : rdata = 48'b000111101111111001100000010000000000000100000000;
			// PEs: 25, 26 -> 25
			// srcs: (1711, 152)(980) 0, (4116) 94 --> (4900) -94:NW2, PEGB2, -, NW2
			10'd142 : rdata = 48'b000100100000001011100000100000000100100000000000;
			// PEs: 24, 25 -> 26
			// srcs: (1782, 139)(3140) 47, (275) -3 --> (3412) -141:PENB, ND3, *, PENB
			10'd143 : rdata = 48'b000111101111111001100000011000000000000100000000;
			// PEs: 25, 26 -> 25
			// srcs: (1791, 153)(1060) -3, (4196) -141 --> (4980) 138:NW3, PEGB2, -, NW3
			10'd144 : rdata = 48'b000100100000001111100000100000000100110000000000;
			// PEs: 24, 25 -> 26
			// srcs: (1820, 140)(3140) 47, (313) -3 --> (3450) -141:PENB, ND11, *, PENB
			10'd145 : rdata = 48'b000111101111111001100001011000000000000100000000;
			// PEs: 25, 26 -> 25
			// srcs: (1829, 154)(1098) 0, (4234) -141 --> (5018) 141:NW11, PEGB2, -, NW11
			10'd146 : rdata = 48'b000100100000101111100000100000000110110000000000;
			// PEs: 24, 25 -> 26
			// srcs: (1862, 141)(3140) 47, (355) -2 --> (3492) -94:PENB, ND4, *, PENB
			10'd147 : rdata = 48'b000111101111111001100000100000000000000100000000;
			// PEs: 25, 26 -> 25
			// srcs: (1871, 155)(1140) 1, (4276) -94 --> (5060) 95:NW4, PEGB2, -, NW4
			10'd148 : rdata = 48'b000100100000010011100000100000000101000000000000;
			// PEs: 24, 25 -> 26
			// srcs: (1944, 142)(3140) 47, (437) -3 --> (3574) -141:PENB, ND5, *, PENB
			10'd149 : rdata = 48'b000111101111111001100000101000000000000100000000;
			// PEs: 25, 26 -> 25
			// srcs: (1953, 156)(1222) -1, (4358) -141 --> (5142) 140:NW5, PEGB2, -, NW5
			10'd150 : rdata = 48'b000100100000010111100000100000000101010000000000;
			// PEs: 24, 25 -> 26
			// srcs: (2000, 143)(3140) 47, (493) 0 --> (3630) 0:PENB, ND12, *, PENB
			10'd151 : rdata = 48'b000111101111111001100001100000000000000100000000;
			// PEs: 25, 26 -> 25
			// srcs: (2009, 157)(1278) 0, (4414) 0 --> (5198) 0:NW12, PEGB2, -, NW12
			10'd152 : rdata = 48'b000100100000110011100000100000000111000000000000;
			// PEs: 24, 25 -> 26
			// srcs: (2024, 144)(3140) 47, (517) -1 --> (3654) -47:PENB, ND6, *, PENB
			10'd153 : rdata = 48'b000111101111111001100000110000000000000100000000;
			// PEs: 25, 26 -> 25
			// srcs: (2033, 158)(1302) -3, (4438) -47 --> (5222) 44:NW6, PEGB2, -, NW6
			10'd154 : rdata = 48'b000100100000011011100000100000000101100000000000;
			// PEs: 24, 25 -> 26
			// srcs: (2104, 145)(3140) 47, (597) 0 --> (3734) 0:PENB, ND7, *, PENB
			10'd155 : rdata = 48'b000111101111111001100000111000000000000100000000;
			// PEs: 25, 26 -> 25
			// srcs: (2113, 159)(1382) -3, (4518) 0 --> (5302) -3:NW7, PEGB2, -, NW7
			10'd156 : rdata = 48'b000100100000011111100000100000000101110000000000;
			// PEs: 24, 25 -> 26
			// srcs: (2184, 146)(3140) 47, (677) -1 --> (3814) -47:PENB, ND13, *, PENB
			10'd157 : rdata = 48'b000111101111111001100001101000000000000100000000;
			// PEs: 24, 25 -> 26
			// srcs: (2186, 147)(3140) 47, (679) 1 --> (3816) 47:PENB, ND8, *, PENB
			10'd158 : rdata = 48'b000111101111111001100001000000000000000100000000;
			// PEs: 25, 26 -> 25
			// srcs: (2193, 160)(1462) -1, (4598) -47 --> (5382) 46:NW13, PEGB2, -, NW13
			10'd159 : rdata = 48'b000100100000110111100000100000000111010000000000;
			// PEs: 25, 26 -> 25
			// srcs: (2195, 161)(1464) 0, (4600) 47 --> (5384) -47:NW8, PEGB2, -, NW8
			10'd160 : rdata = 48'b000100100000100011100000100000000110000000000000;
			// PEs: 24, 25 -> 26
			// srcs: (2266, 148)(3140) 47, (759) -1 --> (3896) -47:PENB, ND9, *, PENB
			10'd161 : rdata = 48'b000111101111111001100001001000000000000100000000;
			// PEs: 25, 26 -> 25
			// srcs: (2275, 162)(1544) 1, (4680) -47 --> (5464) 48:NW9, PEGB2, -, NW9
			10'd162 : rdata = 48'b000100100000100111100000100000000110010000000000;
			default : rdata = 48'b000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 26) begin
	always @(*) begin
		case(address)
			// PEs: 26, 26 -> 24
			// srcs: (1, 0)(35) 1, (820) -1 --> (1604) -1:ND0, NW0, *, PEGB0
			10'd0 : rdata = 48'b000110110000000001000000000000000000000010000000;
			// PEs: 26, 26 -> 24
			// srcs: (2, 1)(115) 1, (900) 1 --> (1684) 1:ND1, NW1, *, PEGB0
			10'd1 : rdata = 48'b000110110000000101000000001000000000000010000000;
			// PEs: 26, 26 -> 24
			// srcs: (3, 2)(197) -3, (982) 1 --> (1766) -3:ND2, NW2, *, PEGB0
			10'd2 : rdata = 48'b000110110000001001000000010000000000000010000000;
			// PEs: 26, 26 -> 24
			// srcs: (4, 3)(277) 0, (1062) -3 --> (1846) 0:ND3, NW3, *, PEGB0
			10'd3 : rdata = 48'b000110110000001101000000011000000000000010000000;
			// PEs: 26, 26 -> 24
			// srcs: (5, 4)(357) -1, (1142) 2 --> (1926) -2:ND4, NW4, *, PEGB0
			10'd4 : rdata = 48'b000110110000010001000000100000000000000010000000;
			// PEs: 26, 26 -> 24
			// srcs: (6, 5)(439) 2, (1224) 0 --> (2008) 0:ND5, NW5, *, PEGB0
			10'd5 : rdata = 48'b000110110000010101000000101000000000000010000000;
			// PEs: 26, 26 -> 24
			// srcs: (7, 6)(519) 2, (1304) -1 --> (2088) -2:ND6, NW6, *, PEGB0
			10'd6 : rdata = 48'b000110110000011001000000110000000000000010000000;
			// PEs: 26, 26 -> 24
			// srcs: (8, 7)(599) 0, (1384) -1 --> (2168) 0:ND7, NW7, *, PEGB0
			10'd7 : rdata = 48'b000110110000011101000000111000000000000010000000;
			// PEs: 26, 26 -> 28
			// srcs: (9, 8)(681) 2, (1466) -1 --> (2250) -2:ND8, NW8, *, PEGB4
			10'd8 : rdata = 48'b000110110000100001000001000000000000000011000000;
			// PEs: 26, 26 -> 31
			// srcs: (10, 9)(761) 2, (1546) -3 --> (2330) -6:ND9, NW9, *, PEGB7
			10'd9 : rdata = 48'b000110110000100101000001001000000000000011110000;
			// PEs: 26, 26 -> 24
			// srcs: (11, 10)(132) -1, (917) 1 --> (1701) -1:ND10, NW10, *, PEGB0
			10'd10 : rdata = 48'b000110110000101001000001010000000000000010000000;
			// PEs: 26, 26 -> 26
			// srcs: (12, 11)(316) -1, (1101) 2 --> (1885) -2:ND11, NW11, *, NI0
			10'd11 : rdata = 48'b000110110000101101000001011100000000000000000000;
			// PEs: 26, 26 -> 26
			// srcs: (13, 12)(500) 0, (1285) 1 --> (2069) 0:ND12, NW12, *, NI1
			10'd12 : rdata = 48'b000110110000110001000001100100001000000000000000;
			// PEs: 26, 26 -> 26
			// srcs: (14, 13)(680) 2, (1465) 0 --> (2249) 0:ND13, NW13, *, NI2
			10'd13 : rdata = 48'b000110110000110101000001101100010000000000000000;
			// PEs: 29 -> 
			// srcs: (15, 19)(2334) 0 --> (2334) 0:PEGB5, pass, 
			10'd14 : rdata = 48'b110001110000101000000000000000000000000000000000;
			// PEs: 28, 26 -> 26
			// srcs: (18, 20)(2333) -4, (2334) 0 --> (3112) -4:PEGB4, ALU, +, NI3
			10'd15 : rdata = 48'b000011110000100000111111111100011000000000000000;
			// PEs: 24 -> 
			// srcs: (19, 14)(1636) 0 --> (1636) 0:PEGB0, pass, 
			10'd16 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 24, 26 -> 25
			// srcs: (28, 15)(1635) -1, (1636) 0 --> (2417) -1:PEGB0, ALU, +, PEGB1
			10'd17 : rdata = 48'b000011110000000000111111111000000000000010010000;
			// PEs: 24 -> 
			// srcs: (49, 16)(1758) 0 --> (1758) 0:PEGB0, pass, 
			10'd18 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 24, 26 -> 24
			// srcs: (58, 17)(1757) -4, (1758) 0 --> (2537) -4:PEGB0, ALU, +, PEGB0
			10'd19 : rdata = 48'b000011110000000000111111111000000000000010000000;
			// PEs: 24, 25 -> 26
			// srcs: (107, 18)(2005) 1, (2006) 3 --> (2785) 4:PEGB0, PENB, +, NI4
			10'd20 : rdata = 48'b000011110000000011011111110100100000000000000000;
			// PEs: 26 -> 24
			// srcs: (137, 21)(1885) -2 --> (1885) -2:NI0, pass, PEGB0
			10'd21 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 25, 26 -> 27
			// srcs: (146, 28)(3026) -2, (2249) 0 --> (3027) -2:PENB, NI2, +, PENB
			10'd22 : rdata = 48'b000011101111111010100000010000000000000100000000;
			// PEs: 26 -> 24
			// srcs: (154, 24)(2785) 4 --> (2785) 4:NI4, pass, PEGB0
			10'd23 : rdata = 48'b110001010000010000000000000000000000000010000000;
			// PEs: 25 -> 
			// srcs: (314, 22)(2698) 5 --> (2698) 5:PENB, pass, 
			10'd24 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 25, 26 -> 24
			// srcs: (321, 23)(2697) 2, (2698) 5 --> (2699) 7:PENB, ALU, +, PEGB0
			10'd25 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 25 -> 
			// srcs: (351, 26)(2944) 7 --> (2944) 7:PENB, pass, 
			10'd26 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 25, 26 -> 24
			// srcs: (358, 27)(2943) 4, (2944) 7 --> (2945) 11:PENB, ALU, +, PEGB0
			10'd27 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 26 -> 25
			// srcs: (612, 25)(2069) 0 --> (2069) 0:NI1, pass, PEGB1
			10'd28 : rdata = 48'b110001010000000100000000000000000000000010010000;
			// PEs: 25 -> 
			// srcs: (628, 30)(2854) 5 --> (2854) 5:PENB, pass, 
			10'd29 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 25, 26 -> 24
			// srcs: (635, 31)(2852) 8, (2854) 5 --> (2855) 13:PENB, ALU, +, PEGB0
			10'd30 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 26 -> 25
			// srcs: (685, 29)(3112) -4 --> (3112) -4:NI3, pass, PEGB1
			10'd31 : rdata = 48'b110001010000001100000000000000000000000010010000;
			// PEs: 26, 25 -> 25
			// srcs: (1543, 46)(3) 1, (3170) 94 --> (3954) 94:NM0, PENB, *, PEGB1
			10'd32 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 24, 26 -> 27
			// srcs: (1545, 32)(3140) 47, (35) 1 --> (3172) 47:PEGB0, ND0, *, PENB
			10'd33 : rdata = 48'b000111110000000001100000000000000000000100000000;
			// PEs: 26, 27 -> 26
			// srcs: (1554, 64)(820) -1, (3956) 47 --> (4740) -48:NW0, PEGB3, -, NW0
			10'd34 : rdata = 48'b000100100000000011100000110000000100000000000000;
			// PEs: 26, 25 -> 25
			// srcs: (1623, 47)(3) 1, (3250) -94 --> (4034) -94:NM0, PENB, *, PEGB1
			10'd35 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 24, 26 -> 27
			// srcs: (1625, 33)(3140) 47, (115) 1 --> (3252) 47:PEGB0, ND1, *, PENB
			10'd36 : rdata = 48'b000111110000000001100000001000000000000100000000;
			// PEs: 26, 27 -> 26
			// srcs: (1634, 65)(900) 1, (4036) 47 --> (4820) -46:NW1, PEGB3, -, NW1
			10'd37 : rdata = 48'b000100100000000111100000110000000100010000000000;
			// PEs: 26, 25 -> 25
			// srcs: (1639, 48)(3) 1, (3266) 94 --> (4050) 94:NM0, PENB, *, PEGB1
			10'd38 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 24, 26 -> 
			// srcs: (1642, 34)(3140) 47, (132) -1 --> (3269) -47:PEGB0, ND10, *, 
			10'd39 : rdata = 48'b000111110000000001100001010000000000000000000000;
			// PEs: 26, 26 -> 
			// srcs: (1645, 49)(3) 1, (3269) -47 --> (4053) -47:NM0, ALU, *, 
			10'd40 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 26, 26 -> 26
			// srcs: (1648, 66)(917) 1, (4053) -47 --> (4837) 48:NW10, ALU, -, NW10
			10'd41 : rdata = 48'b000100100000101000111111111000000110100000000000;
			// PEs: 26, 25 -> 25
			// srcs: (1705, 50)(3) 1, (3332) 94 --> (4116) 94:NM0, PENB, *, PEGB1
			10'd42 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 24, 26 -> 27
			// srcs: (1707, 35)(3140) 47, (197) -3 --> (3334) -141:PEGB0, ND2, *, PENB
			10'd43 : rdata = 48'b000111110000000001100000010000000000000100000000;
			// PEs: 26, 27 -> 26
			// srcs: (1716, 67)(982) 1, (4118) -141 --> (4902) 142:NW2, PEGB3, -, NW2
			10'd44 : rdata = 48'b000100100000001011100000110000000100100000000000;
			// PEs: 26, 25 -> 25
			// srcs: (1785, 51)(3) 1, (3412) -141 --> (4196) -141:NM0, PENB, *, PEGB1
			10'd45 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 24, 26 -> 27
			// srcs: (1787, 36)(3140) 47, (277) 0 --> (3414) 0:PEGB0, ND3, *, PENB
			10'd46 : rdata = 48'b000111110000000001100000011000000000000100000000;
			// PEs: 26, 27 -> 26
			// srcs: (1796, 68)(1062) -3, (4198) 0 --> (4982) -3:NW3, PEGB3, -, NW3
			10'd47 : rdata = 48'b000100100000001111100000110000000100110000000000;
			// PEs: 26, 25 -> 25
			// srcs: (1823, 52)(3) 1, (3450) -141 --> (4234) -141:NM0, PENB, *, PEGB1
			10'd48 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 24, 26 -> 
			// srcs: (1826, 37)(3140) 47, (316) -1 --> (3453) -47:PEGB0, ND11, *, 
			10'd49 : rdata = 48'b000111110000000001100001011000000000000000000000;
			// PEs: 26, 26 -> 
			// srcs: (1829, 53)(3) 1, (3453) -47 --> (4237) -47:NM0, ALU, *, 
			10'd50 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 26, 26 -> 26
			// srcs: (1832, 69)(1101) 2, (4237) -47 --> (5021) 49:NW11, ALU, -, NW11
			10'd51 : rdata = 48'b000100100000101100111111111000000110110000000000;
			// PEs: 26, 25 -> 25
			// srcs: (1865, 54)(3) 1, (3492) -94 --> (4276) -94:NM0, PENB, *, PEGB1
			10'd52 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 24, 26 -> 27
			// srcs: (1867, 38)(3140) 47, (357) -1 --> (3494) -47:PEGB0, ND4, *, PENB
			10'd53 : rdata = 48'b000111110000000001100000100000000000000100000000;
			// PEs: 26, 27 -> 26
			// srcs: (1876, 70)(1142) 2, (4278) -47 --> (5062) 49:NW4, PEGB3, -, NW4
			10'd54 : rdata = 48'b000100100000010011100000110000000101000000000000;
			// PEs: 26, 25 -> 25
			// srcs: (1947, 55)(3) 1, (3574) -141 --> (4358) -141:NM0, PENB, *, PEGB1
			10'd55 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 24, 26 -> 27
			// srcs: (1949, 39)(3140) 47, (439) 2 --> (3576) 94:PEGB0, ND5, *, PENB
			10'd56 : rdata = 48'b000111110000000001100000101000000000000100000000;
			// PEs: 26, 27 -> 26
			// srcs: (1958, 71)(1224) 0, (4360) 94 --> (5144) -94:NW5, PEGB3, -, NW5
			10'd57 : rdata = 48'b000100100000010111100000110000000101010000000000;
			// PEs: 26, 25 -> 25
			// srcs: (2003, 56)(3) 1, (3630) 0 --> (4414) 0:NM0, PENB, *, PEGB1
			10'd58 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 24, 26 -> 
			// srcs: (2010, 40)(3140) 47, (500) 0 --> (3637) 0:PEGB0, ND12, *, 
			10'd59 : rdata = 48'b000111110000000001100001100000000000000000000000;
			// PEs: 26, 26 -> 
			// srcs: (2013, 57)(3) 1, (3637) 0 --> (4421) 0:NM0, ALU, *, 
			10'd60 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 26, 26 -> 26
			// srcs: (2016, 72)(1285) 1, (4421) 0 --> (5205) 1:NW12, ALU, -, NW12
			10'd61 : rdata = 48'b000100100000110000111111111000000111000000000000;
			// PEs: 26, 25 -> 25
			// srcs: (2027, 58)(3) 1, (3654) -47 --> (4438) -47:NM0, PENB, *, PEGB1
			10'd62 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 24, 26 -> 27
			// srcs: (2029, 41)(3140) 47, (519) 2 --> (3656) 94:PEGB0, ND6, *, PENB
			10'd63 : rdata = 48'b000111110000000001100000110000000000000100000000;
			// PEs: 26, 27 -> 26
			// srcs: (2038, 73)(1304) -1, (4440) 94 --> (5224) -95:NW6, PEGB3, -, NW6
			10'd64 : rdata = 48'b000100100000011011100000110000000101100000000000;
			// PEs: 26, 25 -> 25
			// srcs: (2107, 59)(3) 1, (3734) 0 --> (4518) 0:NM0, PENB, *, PEGB1
			10'd65 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 24, 26 -> 27
			// srcs: (2109, 42)(3140) 47, (599) 0 --> (3736) 0:PEGB0, ND7, *, PENB
			10'd66 : rdata = 48'b000111110000000001100000111000000000000100000000;
			// PEs: 26, 27 -> 26
			// srcs: (2118, 74)(1384) -1, (4520) 0 --> (5304) -1:NW7, PEGB3, -, NW7
			10'd67 : rdata = 48'b000100100000011111100000110000000101110000000000;
			// PEs: 26, 25 -> 25
			// srcs: (2187, 60)(3) 1, (3814) -47 --> (4598) -47:NM0, PENB, *, PEGB1
			10'd68 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 26, 25 -> 25
			// srcs: (2189, 61)(3) 1, (3816) 47 --> (4600) 47:NM0, PENB, *, PEGB1
			10'd69 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 24, 26 -> 26
			// srcs: (2190, 43)(3140) 47, (680) 2 --> (3817) 94:PEGB0, ND13, *, NI0
			10'd70 : rdata = 48'b000111110000000001100001101100000000000000000000;
			// PEs: 24, 26 -> 27
			// srcs: (2191, 44)(3140) 47, (681) 2 --> (3818) 94:PEGB0, ND8, *, PENB
			10'd71 : rdata = 48'b000111110000000001100001000000000000000100000000;
			// PEs: 26, 26 -> 
			// srcs: (2193, 62)(3) 1, (3817) 94 --> (4601) 94:NM0, NI0, *, 
			10'd72 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 26, 26 -> 26
			// srcs: (2196, 75)(1465) 0, (4601) 94 --> (5385) -94:NW13, ALU, -, NW13
			10'd73 : rdata = 48'b000100100000110100111111111000000111010000000000;
			// PEs: 26, 27 -> 26
			// srcs: (2200, 76)(1466) -1, (4602) 94 --> (5386) -95:NW8, PEGB3, -, NW8
			10'd74 : rdata = 48'b000100100000100011100000110000000110000000000000;
			// PEs: 26, 25 -> 25
			// srcs: (2269, 63)(3) 1, (3896) -47 --> (4680) -47:NM0, PENB, *, PEGB1
			10'd75 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 24, 26 -> 27
			// srcs: (2271, 45)(3140) 47, (761) 2 --> (3898) 94:PEGB0, ND9, *, PENB
			10'd76 : rdata = 48'b000111110000000001100001001000000000000100000000;
			// PEs: 26, 27 -> 26
			// srcs: (2280, 77)(1546) -3, (4682) 94 --> (5466) -97:NW9, PEGB3, -, NW9
			10'd77 : rdata = 48'b000100100000100111100000110000000110010000000000;
			default : rdata = 48'b000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 27) begin
	always @(*) begin
		case(address)
			// PEs: 27, 27 -> 24
			// srcs: (1, 0)(36) 2, (821) -1 --> (1605) -2:ND0, NW0, *, PEGB0
			10'd0 : rdata = 48'b000110110000000001000000000000000000000010000000;
			// PEs: 27, 27 -> 24
			// srcs: (2, 1)(116) 2, (901) 0 --> (1685) 0:ND1, NW1, *, PEGB0
			10'd1 : rdata = 48'b000110110000000101000000001000000000000010000000;
			// PEs: 27, 27 -> 24
			// srcs: (3, 2)(198) 0, (983) 0 --> (1767) 0:ND2, NW2, *, PEGB0
			10'd2 : rdata = 48'b000110110000001001000000010000000000000010000000;
			// PEs: 27, 27 -> 24
			// srcs: (4, 3)(278) -1, (1063) 0 --> (1847) 0:ND3, NW3, *, PEGB0
			10'd3 : rdata = 48'b000110110000001101000000011000000000000010000000;
			// PEs: 27, 27 -> 24
			// srcs: (5, 4)(358) 2, (1143) -1 --> (1927) -2:ND4, NW4, *, PEGB0
			10'd4 : rdata = 48'b000110110000010001000000100000000000000010000000;
			// PEs: 27, 27 -> 24
			// srcs: (6, 5)(440) -3, (1225) 1 --> (2009) -3:ND5, NW5, *, PEGB0
			10'd5 : rdata = 48'b000110110000010101000000101000000000000010000000;
			// PEs: 27, 27 -> 24
			// srcs: (7, 6)(520) -1, (1305) 0 --> (2089) 0:ND6, NW6, *, PEGB0
			10'd6 : rdata = 48'b000110110000011001000000110000000000000010000000;
			// PEs: 27, 27 -> 24
			// srcs: (8, 7)(600) 2, (1385) -1 --> (2169) -2:ND7, NW7, *, PEGB0
			10'd7 : rdata = 48'b000110110000011101000000111000000000000010000000;
			// PEs: 27, 27 -> 28
			// srcs: (9, 8)(682) 0, (1467) -3 --> (2251) 0:ND8, NW8, *, PENB
			10'd8 : rdata = 48'b000110110000100001000001000000000000000100000000;
			// PEs: 27, 27 -> 31
			// srcs: (10, 9)(762) 0, (1547) 2 --> (2331) 0:ND9, NW9, *, PEGB7
			10'd9 : rdata = 48'b000110110000100101000001001000000000000011110000;
			// PEs: 27, 27 -> 24
			// srcs: (11, 10)(135) 2, (920) -1 --> (1704) -2:ND10, NW10, *, PEGB0
			10'd10 : rdata = 48'b000110110000101001000001010000000000000010000000;
			// PEs: 27, 27 -> 24
			// srcs: (12, 11)(319) 2, (1104) -1 --> (1888) -2:ND11, NW11, *, PEGB0
			10'd11 : rdata = 48'b000110110000101101000001011000000000000010000000;
			// PEs: 27, 27 -> 27
			// srcs: (13, 12)(503) -1, (1288) -2 --> (2072) 2:ND12, NW12, *, NI0
			10'd12 : rdata = 48'b000110110000110001000001100100000000000000000000;
			// PEs: 27, 27 -> 29
			// srcs: (14, 13)(683) -1, (1468) -2 --> (2252) 2:ND13, NW13, *, PEGB5
			10'd13 : rdata = 48'b000110110000110101000001101000000000000011010000;
			// PEs: 24 -> 
			// srcs: (21, 14)(1639) 3 --> (1639) 3:PEGB0, pass, 
			10'd14 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 24, 27 -> 24
			// srcs: (30, 15)(1638) 0, (1639) 3 --> (2419) 3:PEGB0, ALU, +, PEGB0
			10'd15 : rdata = 48'b000011110000000000111111111000000000000010000000;
			// PEs: 24 -> 
			// srcs: (51, 16)(1761) -1 --> (1761) -1:PEGB0, pass, 
			10'd16 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 24, 27 -> 27
			// srcs: (60, 17)(1760) -4, (1761) -1 --> (2539) -5:PEGB0, ALU, +, NI1
			10'd17 : rdata = 48'b000011110000000000111111111100001000000000000000;
			// PEs: 24 -> 
			// srcs: (131, 18)(2085) 0 --> (2085) 0:PEGB0, pass, 
			10'd18 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 27, 25 -> 24
			// srcs: (133, 19)(2085) 0, (2086) 3 --> (2864) 3:ALU, PEGB1, +, PEGB0
			10'd19 : rdata = 48'b000010011111111111100000010000000000000010000000;
			// PEs: 25 -> 
			// srcs: (134, 24)(2857) 1 --> (2857) 1:PEGB1, pass, 
			10'd20 : rdata = 48'b110001110000001000000000000000000000000000000000;
			// PEs: 27, 29 -> 
			// srcs: (136, 25)(2857) 1, (2078) -4 --> (2858) -3:ALU, PEGB5, +, 
			10'd21 : rdata = 48'b000010011111111111100001010000000000000000000000;
			// PEs: 27, 30 -> 24
			// srcs: (142, 26)(2858) -3, (2860) 6 --> (2861) 3:ALU, PEGB6, +, PEGB0
			10'd22 : rdata = 48'b000010011111111111100001100000000000000010000000;
			// PEs: 26, 29 -> 30
			// srcs: (152, 27)(3027) -2, (3029) 0 --> (3030) -2:PENB, PEGB5, +, PEGB6
			10'd23 : rdata = 48'b000011101111111011100001010000000000000011100000;
			// PEs: 24 -> 
			// srcs: (248, 20)(1674) 0 --> (1674) 0:PEGB0, pass, 
			10'd24 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 24, 27 -> 25
			// srcs: (257, 21)(1673) 0, (1674) 0 --> (2455) 0:PEGB0, ALU, +, PEGB1
			10'd25 : rdata = 48'b000011110000000000111111111000000000000010010000;
			// PEs: 27 -> 25
			// srcs: (549, 22)(2539) -5 --> (2539) -5:NI1, pass, PEGB1
			10'd26 : rdata = 48'b110001010000000100000000000000000000000010010000;
			// PEs: 27 -> 25
			// srcs: (620, 23)(2072) 2 --> (2072) 2:NI0, pass, PEGB1
			10'd27 : rdata = 48'b110001010000000000000000000000000000000010010000;
			// PEs: 24, 27 -> 27
			// srcs: (1546, 28)(3140) 47, (36) 2 --> (3173) 94:PEGB0, ND0, *, NI0
			10'd28 : rdata = 48'b000111110000000001100000000100000000000000000000;
			// PEs: 27, 26 -> 26
			// srcs: (1548, 42)(3) 1, (3172) 47 --> (3956) 47:NM0, PENB, *, PEGB2
			10'd29 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 27, 27 -> 
			// srcs: (1549, 43)(3) 1, (3173) 94 --> (3957) 94:NM0, NI0, *, 
			10'd30 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 27, 27 -> 27
			// srcs: (1552, 58)(821) -1, (3957) 94 --> (4741) -95:NW0, ALU, -, NW0
			10'd31 : rdata = 48'b000100100000000000111111111000000100000000000000;
			// PEs: 24, 27 -> 28
			// srcs: (1626, 29)(3140) 47, (116) 2 --> (3253) 94:PEGB0, ND1, *, PENB
			10'd32 : rdata = 48'b000111110000000001100000001000000000000100000000;
			// PEs: 27, 26 -> 26
			// srcs: (1628, 44)(3) 1, (3252) 47 --> (4036) 47:NM0, PENB, *, PEGB2
			10'd33 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 27, 28 -> 27
			// srcs: (1635, 59)(901) 0, (4037) 94 --> (4821) -94:NW1, PEGB4, -, NW1
			10'd34 : rdata = 48'b000100100000000111100001000000000100010000000000;
			// PEs: 24, 27 -> 
			// srcs: (1645, 30)(3140) 47, (135) 2 --> (3272) 94:PEGB0, ND10, *, 
			10'd35 : rdata = 48'b000111110000000001100001010000000000000000000000;
			// PEs: 27, 27 -> 
			// srcs: (1648, 45)(3) 1, (3272) 94 --> (4056) 94:NM0, ALU, *, 
			10'd36 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 27, 27 -> 27
			// srcs: (1651, 60)(920) -1, (4056) 94 --> (4840) -95:NW10, ALU, -, NW10
			10'd37 : rdata = 48'b000100100000101000111111111000000110100000000000;
			// PEs: 24, 27 -> 28
			// srcs: (1708, 31)(3140) 47, (198) 0 --> (3335) 0:PEGB0, ND2, *, PENB
			10'd38 : rdata = 48'b000111110000000001100000010000000000000100000000;
			// PEs: 27, 26 -> 26
			// srcs: (1710, 46)(3) 1, (3334) -141 --> (4118) -141:NM0, PENB, *, PEGB2
			10'd39 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 27, 28 -> 27
			// srcs: (1717, 61)(983) 0, (4119) 0 --> (4903) 0:NW2, PEGB4, -, NW2
			10'd40 : rdata = 48'b000100100000001011100001000000000100100000000000;
			// PEs: 24, 27 -> 28
			// srcs: (1788, 32)(3140) 47, (278) -1 --> (3415) -47:PEGB0, ND3, *, PENB
			10'd41 : rdata = 48'b000111110000000001100000011000000000000100000000;
			// PEs: 27, 26 -> 26
			// srcs: (1790, 47)(3) 1, (3414) 0 --> (4198) 0:NM0, PENB, *, PEGB2
			10'd42 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 27, 28 -> 27
			// srcs: (1797, 62)(1063) 0, (4199) -47 --> (4983) 47:NW3, PEGB4, -, NW3
			10'd43 : rdata = 48'b000100100000001111100001000000000100110000000000;
			// PEs: 24, 27 -> 
			// srcs: (1829, 33)(3140) 47, (319) 2 --> (3456) 94:PEGB0, ND11, *, 
			10'd44 : rdata = 48'b000111110000000001100001011000000000000000000000;
			// PEs: 27, 27 -> 
			// srcs: (1832, 48)(3) 1, (3456) 94 --> (4240) 94:NM0, ALU, *, 
			10'd45 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 27, 27 -> 27
			// srcs: (1835, 63)(1104) -1, (4240) 94 --> (5024) -95:NW11, ALU, -, NW11
			10'd46 : rdata = 48'b000100100000101100111111111000000110110000000000;
			// PEs: 24, 27 -> 28
			// srcs: (1868, 34)(3140) 47, (358) 2 --> (3495) 94:PEGB0, ND4, *, PENB
			10'd47 : rdata = 48'b000111110000000001100000100000000000000100000000;
			// PEs: 27, 26 -> 26
			// srcs: (1870, 49)(3) 1, (3494) -47 --> (4278) -47:NM0, PENB, *, PEGB2
			10'd48 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 27, 28 -> 27
			// srcs: (1877, 64)(1143) -1, (4279) 94 --> (5063) -95:NW4, PEGB4, -, NW4
			10'd49 : rdata = 48'b000100100000010011100001000000000101000000000000;
			// PEs: 24, 27 -> 28
			// srcs: (1950, 35)(3140) 47, (440) -3 --> (3577) -141:PEGB0, ND5, *, PENB
			10'd50 : rdata = 48'b000111110000000001100000101000000000000100000000;
			// PEs: 27, 26 -> 26
			// srcs: (1952, 50)(3) 1, (3576) 94 --> (4360) 94:NM0, PENB, *, PEGB2
			10'd51 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 27, 28 -> 27
			// srcs: (1959, 65)(1225) 1, (4361) -141 --> (5145) 142:NW5, PEGB4, -, NW5
			10'd52 : rdata = 48'b000100100000010111100001000000000101010000000000;
			// PEs: 24, 27 -> 
			// srcs: (2013, 36)(3140) 47, (503) -1 --> (3640) -47:PEGB0, ND12, *, 
			10'd53 : rdata = 48'b000111110000000001100001100000000000000000000000;
			// PEs: 27, 27 -> 
			// srcs: (2016, 51)(3) 1, (3640) -47 --> (4424) -47:NM0, ALU, *, 
			10'd54 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 27, 27 -> 27
			// srcs: (2019, 66)(1288) -2, (4424) -47 --> (5208) 45:NW12, ALU, -, NW12
			10'd55 : rdata = 48'b000100100000110000111111111000000111000000000000;
			// PEs: 24, 27 -> 28
			// srcs: (2030, 37)(3140) 47, (520) -1 --> (3657) -47:PEGB0, ND6, *, PENB
			10'd56 : rdata = 48'b000111110000000001100000110000000000000100000000;
			// PEs: 27, 26 -> 26
			// srcs: (2032, 52)(3) 1, (3656) 94 --> (4440) 94:NM0, PENB, *, PEGB2
			10'd57 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 27, 28 -> 27
			// srcs: (2039, 67)(1305) 0, (4441) -47 --> (5225) 47:NW6, PEGB4, -, NW6
			10'd58 : rdata = 48'b000100100000011011100001000000000101100000000000;
			// PEs: 24, 27 -> 27
			// srcs: (2110, 38)(3140) 47, (600) 2 --> (3737) 94:PEGB0, ND7, *, NI0
			10'd59 : rdata = 48'b000111110000000001100000111100000000000000000000;
			// PEs: 27, 26 -> 26
			// srcs: (2112, 53)(3) 1, (3736) 0 --> (4520) 0:NM0, PENB, *, PEGB2
			10'd60 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 27, 27 -> 
			// srcs: (2113, 54)(3) 1, (3737) 94 --> (4521) 94:NM0, NI0, *, 
			10'd61 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 27, 27 -> 27
			// srcs: (2116, 68)(1385) -1, (4521) 94 --> (5305) -95:NW7, ALU, -, NW7
			10'd62 : rdata = 48'b000100100000011100111111111000000101110000000000;
			// PEs: 24, 27 -> 28
			// srcs: (2192, 39)(3140) 47, (682) 0 --> (3819) 0:PEGB0, ND8, *, PENB
			10'd63 : rdata = 48'b000111110000000001100001000000000000000100000000;
			// PEs: 24, 27 -> 27
			// srcs: (2193, 40)(3140) 47, (683) -1 --> (3820) -47:PEGB0, ND13, *, NI0
			10'd64 : rdata = 48'b000111110000000001100001101100000000000000000000;
			// PEs: 27, 26 -> 26
			// srcs: (2194, 55)(3) 1, (3818) 94 --> (4602) 94:NM0, PENB, *, PEGB2
			10'd65 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 27, 27 -> 
			// srcs: (2196, 56)(3) 1, (3820) -47 --> (4604) -47:NM0, NI0, *, 
			10'd66 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 27, 27 -> 27
			// srcs: (2199, 70)(1468) -2, (4604) -47 --> (5388) 45:NW13, ALU, -, NW13
			10'd67 : rdata = 48'b000100100000110100111111111000000111010000000000;
			// PEs: 27, 28 -> 27
			// srcs: (2201, 69)(1467) -3, (4603) 0 --> (5387) -3:NW8, PEGB4, -, NW8
			10'd68 : rdata = 48'b000100100000100011100001000000000110000000000000;
			// PEs: 24, 27 -> 28
			// srcs: (2272, 41)(3140) 47, (762) 0 --> (3899) 0:PEGB0, ND9, *, PENB
			10'd69 : rdata = 48'b000111110000000001100001001000000000000100000000;
			// PEs: 27, 26 -> 26
			// srcs: (2274, 57)(3) 1, (3898) 94 --> (4682) 94:NM0, PENB, *, PEGB2
			10'd70 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 27, 28 -> 27
			// srcs: (2281, 71)(1547) 2, (4683) 0 --> (5467) 2:NW9, PEGB4, -, NW9
			10'd71 : rdata = 48'b000100100000100111100001000000000110010000000000;
			default : rdata = 48'b000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 28) begin
	always @(*) begin
		case(address)
			// PEs: 28, 28 -> 24
			// srcs: (1, 0)(38) 2, (823) -1 --> (1607) -2:ND0, NW0, *, PEGB0
			10'd0 : rdata = 48'b000110110000000001000000000000000000000010000000;
			// PEs: 28, 28 -> 24
			// srcs: (2, 1)(118) -2, (903) 1 --> (1687) -2:ND1, NW1, *, PEGB0
			10'd1 : rdata = 48'b000110110000000101000000001000000000000010000000;
			// PEs: 28, 28 -> 28
			// srcs: (3, 2)(200) 2, (985) -1 --> (1769) -2:ND2, NW2, *, NI0
			10'd2 : rdata = 48'b000110110000001001000000010100000000000000000000;
			// PEs: 28, 28 -> 24
			// srcs: (4, 3)(280) 0, (1065) 1 --> (1849) 0:ND3, NW3, *, PEGB0
			10'd3 : rdata = 48'b000110110000001101000000011000000000000010000000;
			// PEs: 28, 28 -> 24
			// srcs: (5, 4)(360) -1, (1145) -2 --> (1929) 2:ND4, NW4, *, PEGB0
			10'd4 : rdata = 48'b000110110000010001000000100000000000000010000000;
			// PEs: 28, 28 -> 24
			// srcs: (6, 5)(442) 2, (1227) -3 --> (2011) -6:ND5, NW5, *, PEGB0
			10'd5 : rdata = 48'b000110110000010101000000101000000000000010000000;
			// PEs: 28, 28 -> 24
			// srcs: (7, 6)(522) 0, (1307) 2 --> (2091) 0:ND6, NW6, *, PEGB0
			10'd6 : rdata = 48'b000110110000011001000000110000000000000010000000;
			// PEs: 28, 28 -> 24
			// srcs: (8, 7)(602) 2, (1387) 2 --> (2171) 4:ND7, NW7, *, PEGB0
			10'd7 : rdata = 48'b000110110000011101000000111000000000000010000000;
			// PEs: 28, 28 -> 30
			// srcs: (9, 8)(684) -1, (1469) -1 --> (2253) 1:ND8, NW8, *, PEGB6
			10'd8 : rdata = 48'b000110110000100001000001000000000000000011100000;
			// PEs: 28, 28 -> 26
			// srcs: (10, 9)(764) -2, (1549) 2 --> (2333) -4:ND9, NW9, *, PEGB2
			10'd9 : rdata = 48'b000110110000100101000001001000000000000010100000;
			// PEs: 28, 28 -> 28
			// srcs: (11, 10)(138) -3, (923) -3 --> (1707) 9:ND10, NW10, *, NI1
			10'd10 : rdata = 48'b000110110000101001000001010100001000000000000000;
			// PEs: 28, 28 -> 28
			// srcs: (12, 11)(322) 1, (1107) 2 --> (1891) 2:ND11, NW11, *, NI2
			10'd11 : rdata = 48'b000110110000101101000001011100010000000000000000;
			// PEs: 28, 28 -> 25
			// srcs: (13, 12)(506) -1, (1291) 1 --> (2075) -1:ND12, NW12, *, PEGB1
			10'd12 : rdata = 48'b000110110000110001000001100000000000000010010000;
			// PEs: 28, 28 -> 28
			// srcs: (14, 13)(686) 0, (1471) 1 --> (2255) 0:ND13, NW13, *, NI3
			10'd13 : rdata = 48'b000110110000110101000001101100011000000000000000;
			// PEs: 26, 27 -> 29
			// srcs: (15, 18)(2250) -2, (2251) 0 --> (3028) -2:PEGB2, PENB, +, PENB
			10'd14 : rdata = 48'b000011110000010011011111110000000000000100000000;
			// PEs: 31 -> 
			// srcs: (16, 19)(2337) 0 --> (2337) 0:PEGB7, pass, 
			10'd15 : rdata = 48'b110001110000111000000000000000000000000000000000;
			// PEs: 30, 28 -> 28
			// srcs: (18, 20)(2336) 4, (2337) 0 --> (3114) 4:PEGB6, ALU, +, NI4
			10'd16 : rdata = 48'b000011110000110000111111111100100000000000000000;
			// PEs: 30, 28 -> 29
			// srcs: (21, 25)(3031) 5, (2255) 0 --> (3032) 5:PEGB6, NI3, +, PENB
			10'd17 : rdata = 48'b000011110000110010100000011000000000000100000000;
			// PEs: 24 -> 
			// srcs: (23, 14)(1642) 1 --> (1642) 1:PEGB0, pass, 
			10'd18 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 24, 28 -> 24
			// srcs: (32, 15)(1641) -6, (1642) 1 --> (2422) -5:PEGB0, ALU, +, PEGB0
			10'd19 : rdata = 48'b000011110000000000111111111000000000000010000000;
			// PEs: 24 -> 
			// srcs: (56, 16)(1835) -2 --> (1835) -2:PEGB0, pass, 
			10'd20 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 24, 28 -> 28
			// srcs: (65, 17)(1834) 0, (1835) -2 --> (2614) -2:PEGB0, ALU, +, NI3
			10'd21 : rdata = 48'b000011110000000000111111111100011000000000000000;
			// PEs: 28 -> 24
			// srcs: (106, 21)(1769) -2 --> (1769) -2:NI0, pass, PEGB0
			10'd22 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 28 -> 24
			// srcs: (116, 22)(1707) 9 --> (1707) 9:NI1, pass, PEGB0
			10'd23 : rdata = 48'b110001010000000100000000000000000000000010000000;
			// PEs: 28 -> 24
			// srcs: (122, 24)(1891) 2 --> (1891) 2:NI2, pass, PEGB0
			10'd24 : rdata = 48'b110001010000001000000000000000000000000010000000;
			// PEs: 28 -> 24
			// srcs: (137, 23)(2614) -2 --> (2614) -2:NI3, pass, PEGB0
			10'd25 : rdata = 48'b110001010000001100000000000000000000000010000000;
			// PEs: 28 -> 24
			// srcs: (154, 26)(3114) 4 --> (3114) 4:NI4, pass, PEGB0
			10'd26 : rdata = 48'b110001010000010000000000000000000000000010000000;
			// PEs: 24 -> 
			// srcs: (790, 27)(3019) -11 --> (3019) -11:PEGB0, pass, 
			10'd27 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 28, 29 -> 31
			// srcs: (797, 28)(3019) -11, (3024) -2 --> (3025) -13:ALU, PEGB5, +, PEGB7
			10'd28 : rdata = 48'b000010011111111111100001010000000000000011110000;
			// PEs: 24, 28 -> 
			// srcs: (1548, 29)(3140) 47, (38) 2 --> (3175) 94:PEGB0, ND0, *, 
			10'd29 : rdata = 48'b000111110000000001100000000000000000000000000000;
			// PEs: 28, 28 -> 
			// srcs: (1551, 43)(3) 1, (3175) 94 --> (3959) 94:NM0, ALU, *, 
			10'd30 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 28, 28 -> 28
			// srcs: (1554, 58)(823) -1, (3959) 94 --> (4743) -95:NW0, ALU, -, NW0
			10'd31 : rdata = 48'b000100100000000000111111111000000100000000000000;
			// PEs: 24, 28 -> 29
			// srcs: (1628, 30)(3140) 47, (118) -2 --> (3255) -94:PEGB0, ND1, *, PENB
			10'd32 : rdata = 48'b000111110000000001100000001000000000000100000000;
			// PEs: 28, 27 -> 27
			// srcs: (1629, 44)(3) 1, (3253) 94 --> (4037) 94:NM0, PENB, *, PEGB3
			10'd33 : rdata = 48'b000111000000000011011111110000000000000010110000;
			// PEs: 28, 29 -> 28
			// srcs: (1637, 59)(903) 1, (4039) -94 --> (4823) 95:NW1, PEGB5, -, NW1
			10'd34 : rdata = 48'b000100100000000111100001010000000100010000000000;
			// PEs: 24, 28 -> 
			// srcs: (1648, 31)(3140) 47, (138) -3 --> (3275) -141:PEGB0, ND10, *, 
			10'd35 : rdata = 48'b000111110000000001100001010000000000000000000000;
			// PEs: 28, 28 -> 
			// srcs: (1651, 45)(3) 1, (3275) -141 --> (4059) -141:NM0, ALU, *, 
			10'd36 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 28, 28 -> 28
			// srcs: (1654, 60)(923) -3, (4059) -141 --> (4843) 138:NW10, ALU, -, NW10
			10'd37 : rdata = 48'b000100100000101000111111111000000110100000000000;
			// PEs: 24, 28 -> 29
			// srcs: (1710, 32)(3140) 47, (200) 2 --> (3337) 94:PEGB0, ND2, *, PENB
			10'd38 : rdata = 48'b000111110000000001100000010000000000000100000000;
			// PEs: 28, 27 -> 27
			// srcs: (1711, 46)(3) 1, (3335) 0 --> (4119) 0:NM0, PENB, *, PEGB3
			10'd39 : rdata = 48'b000111000000000011011111110000000000000010110000;
			// PEs: 28, 29 -> 28
			// srcs: (1719, 61)(985) -1, (4121) 94 --> (4905) -95:NW2, PEGB5, -, NW2
			10'd40 : rdata = 48'b000100100000001011100001010000000100100000000000;
			// PEs: 24, 28 -> 29
			// srcs: (1790, 33)(3140) 47, (280) 0 --> (3417) 0:PEGB0, ND3, *, PENB
			10'd41 : rdata = 48'b000111110000000001100000011000000000000100000000;
			// PEs: 28, 27 -> 27
			// srcs: (1791, 47)(3) 1, (3415) -47 --> (4199) -47:NM0, PENB, *, PEGB3
			10'd42 : rdata = 48'b000111000000000011011111110000000000000010110000;
			// PEs: 28, 29 -> 28
			// srcs: (1799, 62)(1065) 1, (4201) 0 --> (4985) 1:NW3, PEGB5, -, NW3
			10'd43 : rdata = 48'b000100100000001111100001010000000100110000000000;
			// PEs: 24, 28 -> 
			// srcs: (1832, 34)(3140) 47, (322) 1 --> (3459) 47:PEGB0, ND11, *, 
			10'd44 : rdata = 48'b000111110000000001100001011000000000000000000000;
			// PEs: 28, 28 -> 
			// srcs: (1835, 48)(3) 1, (3459) 47 --> (4243) 47:NM0, ALU, *, 
			10'd45 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 28, 28 -> 28
			// srcs: (1838, 63)(1107) 2, (4243) 47 --> (5027) -45:NW11, ALU, -, NW11
			10'd46 : rdata = 48'b000100100000101100111111111000000110110000000000;
			// PEs: 24, 28 -> 29
			// srcs: (1870, 35)(3140) 47, (360) -1 --> (3497) -47:PEGB0, ND4, *, PENB
			10'd47 : rdata = 48'b000111110000000001100000100000000000000100000000;
			// PEs: 28, 27 -> 27
			// srcs: (1871, 49)(3) 1, (3495) 94 --> (4279) 94:NM0, PENB, *, PEGB3
			10'd48 : rdata = 48'b000111000000000011011111110000000000000010110000;
			// PEs: 28, 29 -> 28
			// srcs: (1879, 64)(1145) -2, (4281) -47 --> (5065) 45:NW4, PEGB5, -, NW4
			10'd49 : rdata = 48'b000100100000010011100001010000000101000000000000;
			// PEs: 24, 28 -> 29
			// srcs: (1952, 36)(3140) 47, (442) 2 --> (3579) 94:PEGB0, ND5, *, PENB
			10'd50 : rdata = 48'b000111110000000001100000101000000000000100000000;
			// PEs: 28, 27 -> 27
			// srcs: (1953, 50)(3) 1, (3577) -141 --> (4361) -141:NM0, PENB, *, PEGB3
			10'd51 : rdata = 48'b000111000000000011011111110000000000000010110000;
			// PEs: 28, 29 -> 28
			// srcs: (1961, 65)(1227) -3, (4363) 94 --> (5147) -97:NW5, PEGB5, -, NW5
			10'd52 : rdata = 48'b000100100000010111100001010000000101010000000000;
			// PEs: 24, 28 -> 
			// srcs: (2016, 37)(3140) 47, (506) -1 --> (3643) -47:PEGB0, ND12, *, 
			10'd53 : rdata = 48'b000111110000000001100001100000000000000000000000;
			// PEs: 28, 28 -> 
			// srcs: (2019, 51)(3) 1, (3643) -47 --> (4427) -47:NM0, ALU, *, 
			10'd54 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 28, 28 -> 28
			// srcs: (2022, 66)(1291) 1, (4427) -47 --> (5211) 48:NW12, ALU, -, NW12
			10'd55 : rdata = 48'b000100100000110000111111111000000111000000000000;
			// PEs: 24, 28 -> 28
			// srcs: (2032, 38)(3140) 47, (522) 0 --> (3659) 0:PEGB0, ND6, *, NI0
			10'd56 : rdata = 48'b000111110000000001100000110100000000000000000000;
			// PEs: 28, 27 -> 27
			// srcs: (2033, 52)(3) 1, (3657) -47 --> (4441) -47:NM0, PENB, *, PEGB3
			10'd57 : rdata = 48'b000111000000000011011111110000000000000010110000;
			// PEs: 28, 28 -> 
			// srcs: (2035, 53)(3) 1, (3659) 0 --> (4443) 0:NM0, NI0, *, 
			10'd58 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 28, 28 -> 28
			// srcs: (2038, 67)(1307) 2, (4443) 0 --> (5227) 2:NW6, ALU, -, NW6
			10'd59 : rdata = 48'b000100100000011000111111111000000101100000000000;
			// PEs: 24, 28 -> 
			// srcs: (2112, 39)(3140) 47, (602) 2 --> (3739) 94:PEGB0, ND7, *, 
			10'd60 : rdata = 48'b000111110000000001100000111000000000000000000000;
			// PEs: 28, 28 -> 
			// srcs: (2115, 54)(3) 1, (3739) 94 --> (4523) 94:NM0, ALU, *, 
			10'd61 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 28, 28 -> 28
			// srcs: (2118, 68)(1387) 2, (4523) 94 --> (5307) -92:NW7, ALU, -, NW7
			10'd62 : rdata = 48'b000100100000011100111111111000000101110000000000;
			// PEs: 24, 28 -> 29
			// srcs: (2194, 40)(3140) 47, (684) -1 --> (3821) -47:PEGB0, ND8, *, PENB
			10'd63 : rdata = 48'b000111110000000001100001000000000000000100000000;
			// PEs: 28, 27 -> 27
			// srcs: (2195, 55)(3) 1, (3819) 0 --> (4603) 0:NM0, PENB, *, PEGB3
			10'd64 : rdata = 48'b000111000000000011011111110000000000000010110000;
			// PEs: 24, 28 -> 
			// srcs: (2196, 41)(3140) 47, (686) 0 --> (3823) 0:PEGB0, ND13, *, 
			10'd65 : rdata = 48'b000111110000000001100001101000000000000000000000;
			// PEs: 28, 28 -> 
			// srcs: (2199, 56)(3) 1, (3823) 0 --> (4607) 0:NM0, ALU, *, 
			10'd66 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 28, 28 -> 28
			// srcs: (2202, 70)(1471) 1, (4607) 0 --> (5391) 1:NW13, ALU, -, NW13
			10'd67 : rdata = 48'b000100100000110100111111111000000111010000000000;
			// PEs: 28, 29 -> 28
			// srcs: (2203, 69)(1469) -1, (4605) -47 --> (5389) 46:NW8, PEGB5, -, NW8
			10'd68 : rdata = 48'b000100100000100011100001010000000110000000000000;
			// PEs: 24, 28 -> 29
			// srcs: (2274, 42)(3140) 47, (764) -2 --> (3901) -94:PEGB0, ND9, *, PENB
			10'd69 : rdata = 48'b000111110000000001100001001000000000000100000000;
			// PEs: 28, 27 -> 27
			// srcs: (2275, 57)(3) 1, (3899) 0 --> (4683) 0:NM0, PENB, *, PEGB3
			10'd70 : rdata = 48'b000111000000000011011111110000000000000010110000;
			// PEs: 28, 29 -> 28
			// srcs: (2283, 71)(1549) 2, (4685) -94 --> (5469) 96:NW9, PEGB5, -, NW9
			10'd71 : rdata = 48'b000100100000100111100001010000000110010000000000;
			default : rdata = 48'b000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 29) begin
	always @(*) begin
		case(address)
			// PEs: 29, 29 -> 24
			// srcs: (1, 0)(39) -3, (824) 0 --> (1608) 0:ND0, NW0, *, PEGB0
			10'd0 : rdata = 48'b000110110000000001000000000000000000000010000000;
			// PEs: 29, 29 -> 24
			// srcs: (2, 1)(119) -3, (904) 1 --> (1688) -3:ND1, NW1, *, PEGB0
			10'd1 : rdata = 48'b000110110000000101000000001000000000000010000000;
			// PEs: 29, 29 -> 29
			// srcs: (3, 2)(201) 0, (986) -1 --> (1770) 0:ND2, NW2, *, NI0
			10'd2 : rdata = 48'b000110110000001001000000010100000000000000000000;
			// PEs: 29, 29 -> 24
			// srcs: (4, 3)(281) -3, (1066) -1 --> (1850) 3:ND3, NW3, *, PEGB0
			10'd3 : rdata = 48'b000110110000001101000000011000000000000010000000;
			// PEs: 29, 29 -> 24
			// srcs: (5, 4)(361) -3, (1146) 1 --> (1930) -3:ND4, NW4, *, PEGB0
			10'd4 : rdata = 48'b000110110000010001000000100000000000000010000000;
			// PEs: 29, 29 -> 24
			// srcs: (6, 5)(443) 2, (1228) -2 --> (2012) -4:ND5, NW5, *, PEGB0
			10'd5 : rdata = 48'b000110110000010101000000101000000000000010000000;
			// PEs: 29, 29 -> 24
			// srcs: (7, 6)(523) -1, (1308) 0 --> (2092) 0:ND6, NW6, *, PEGB0
			10'd6 : rdata = 48'b000110110000011001000000110000000000000010000000;
			// PEs: 29, 29 -> 24
			// srcs: (8, 7)(603) 0, (1388) 2 --> (2172) 0:ND7, NW7, *, PEGB0
			10'd7 : rdata = 48'b000110110000011101000000111000000000000010000000;
			// PEs: 29, 29 -> 30
			// srcs: (9, 8)(685) 2, (1470) 2 --> (2254) 4:ND8, NW8, *, PENB
			10'd8 : rdata = 48'b000110110000100001000001000000000000000100000000;
			// PEs: 29, 29 -> 26
			// srcs: (10, 9)(765) 0, (1550) -3 --> (2334) 0:ND9, NW9, *, PEGB2
			10'd9 : rdata = 48'b000110110000100101000001001000000000000010100000;
			// PEs: 29, 29 -> 29
			// srcs: (11, 10)(141) -2, (926) -1 --> (1710) 2:ND10, NW10, *, NI1
			10'd10 : rdata = 48'b000110110000101001000001010100001000000000000000;
			// PEs: 29, 29 -> 29
			// srcs: (12, 11)(325) -2, (1110) -2 --> (1894) 4:ND11, NW11, *, NI2
			10'd11 : rdata = 48'b000110110000101101000001011100010000000000000000;
			// PEs: 29, 29 -> 27
			// srcs: (13, 12)(509) 2, (1294) -2 --> (2078) -4:ND12, NW12, *, PEGB3
			10'd12 : rdata = 48'b000110110000110001000001100000000000000010110000;
			// PEs: 29, 29 -> 29
			// srcs: (14, 13)(689) 2, (1474) 1 --> (2258) 2:ND13, NW13, *, NI3
			10'd13 : rdata = 48'b000110110000110101000001101100011000000000000000;
			// PEs: 31 -> 
			// srcs: (15, 18)(2257) 2 --> (2257) 2:PEGB7, pass, 
			10'd14 : rdata = 48'b110001110000111000000000000000000000000000000000;
			// PEs: 30, 29 -> 
			// srcs: (17, 19)(2256) -3, (2257) 2 --> (3033) -1:PEGB6, ALU, +, 
			10'd15 : rdata = 48'b000011110000110000111111111000000000000000000000;
			// PEs: 29, 29 -> 29
			// srcs: (20, 25)(3033) -1, (2258) 2 --> (3034) 1:ALU, NI3, +, NI4
			10'd16 : rdata = 48'b000010011111111110100000011100100000000000000000;
			// PEs: 28, 27 -> 27
			// srcs: (21, 24)(3028) -2, (2252) 2 --> (3029) 0:PENB, PEGB3, +, PEGB3
			10'd17 : rdata = 48'b000011101111111011100000110000000000000010110000;
			// PEs: 28, 29 -> 30
			// srcs: (24, 28)(3032) 5, (3034) 1 --> (3035) 6:PENB, NI4, +, PENB
			10'd18 : rdata = 48'b000011101111111010100000100000000000000100000000;
			// PEs: 24 -> 
			// srcs: (25, 14)(1645) -4 --> (1645) -4:PEGB0, pass, 
			10'd19 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 24, 29 -> 24
			// srcs: (34, 15)(1644) -1, (1645) -4 --> (2424) -5:PEGB0, ALU, +, PEGB0
			10'd20 : rdata = 48'b000011110000000000111111111000000000000010000000;
			// PEs: 24 -> 
			// srcs: (63, 16)(1838) 3 --> (1838) 3:PEGB0, pass, 
			10'd21 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 24, 29 -> 29
			// srcs: (72, 17)(1837) 1, (1838) 3 --> (2617) 4:PEGB0, ALU, +, NI3
			10'd22 : rdata = 48'b000011110000000000111111111100011000000000000000;
			// PEs: 29 -> 24
			// srcs: (114, 20)(1770) 0 --> (1770) 0:NI0, pass, PEGB0
			10'd23 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 29 -> 24
			// srcs: (116, 21)(1710) 2 --> (1710) 2:NI1, pass, PEGB0
			10'd24 : rdata = 48'b110001010000000100000000000000000000000010000000;
			// PEs: 29 -> 24
			// srcs: (122, 23)(1894) 4 --> (1894) 4:NI2, pass, PEGB0
			10'd25 : rdata = 48'b110001010000001000000000000000000000000010000000;
			// PEs: 29 -> 24
			// srcs: (137, 22)(2617) 4 --> (2617) 4:NI3, pass, PEGB0
			10'd26 : rdata = 48'b110001010000001100000000000000000000000010000000;
			// PEs: 24 -> 
			// srcs: (780, 26)(3021) -1 --> (3021) -1:PEGB0, pass, 
			10'd27 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 29, 25 -> 28
			// srcs: (782, 27)(3021) -1, (3023) -1 --> (3024) -2:ALU, PEGB1, +, PEGB4
			10'd28 : rdata = 48'b000010011111111111100000010000000000000011000000;
			// PEs: 24, 29 -> 30
			// srcs: (1549, 29)(3140) 47, (39) -3 --> (3176) -141:PEGB0, ND0, *, PENB
			10'd29 : rdata = 48'b000111110000000001100000000000000000000100000000;
			// PEs: 29, 30 -> 29
			// srcs: (1558, 58)(824) 0, (3960) -141 --> (4744) 141:NW0, PEGB6, -, NW0
			10'd30 : rdata = 48'b000100100000000011100001100000000100000000000000;
			// PEs: 24, 29 -> 30
			// srcs: (1629, 30)(3140) 47, (119) -3 --> (3256) -141:PEGB0, ND1, *, PENB
			10'd31 : rdata = 48'b000111110000000001100000001000000000000100000000;
			// PEs: 29, 28 -> 28
			// srcs: (1631, 43)(3) 1, (3255) -94 --> (4039) -94:NM0, PENB, *, PEGB4
			10'd32 : rdata = 48'b000111000000000011011111110000000000000011000000;
			// PEs: 29, 30 -> 29
			// srcs: (1638, 59)(904) 1, (4040) -141 --> (4824) 142:NW1, PEGB6, -, NW1
			10'd33 : rdata = 48'b000100100000000111100001100000000100010000000000;
			// PEs: 24, 29 -> 
			// srcs: (1651, 31)(3140) 47, (141) -2 --> (3278) -94:PEGB0, ND10, *, 
			10'd34 : rdata = 48'b000111110000000001100001010000000000000000000000;
			// PEs: 29, 29 -> 
			// srcs: (1654, 44)(3) 1, (3278) -94 --> (4062) -94:NM0, ALU, *, 
			10'd35 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 29, 29 -> 29
			// srcs: (1657, 60)(926) -1, (4062) -94 --> (4846) 93:NW10, ALU, -, NW10
			10'd36 : rdata = 48'b000100100000101000111111111000000110100000000000;
			// PEs: 24, 29 -> 29
			// srcs: (1711, 32)(3140) 47, (201) 0 --> (3338) 0:PEGB0, ND2, *, NI0
			10'd37 : rdata = 48'b000111110000000001100000010100000000000000000000;
			// PEs: 29, 28 -> 28
			// srcs: (1713, 45)(3) 1, (3337) 94 --> (4121) 94:NM0, PENB, *, PEGB4
			10'd38 : rdata = 48'b000111000000000011011111110000000000000011000000;
			// PEs: 29, 29 -> 
			// srcs: (1714, 46)(3) 1, (3338) 0 --> (4122) 0:NM0, NI0, *, 
			10'd39 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 29, 29 -> 29
			// srcs: (1717, 61)(986) -1, (4122) 0 --> (4906) -1:NW2, ALU, -, NW2
			10'd40 : rdata = 48'b000100100000001000111111111000000100100000000000;
			// PEs: 24, 29 -> 30
			// srcs: (1791, 33)(3140) 47, (281) -3 --> (3418) -141:PEGB0, ND3, *, PENB
			10'd41 : rdata = 48'b000111110000000001100000011000000000000100000000;
			// PEs: 29, 28 -> 28
			// srcs: (1793, 47)(3) 1, (3417) 0 --> (4201) 0:NM0, PENB, *, PEGB4
			10'd42 : rdata = 48'b000111000000000011011111110000000000000011000000;
			// PEs: 29, 30 -> 29
			// srcs: (1800, 62)(1066) -1, (4202) -141 --> (4986) 140:NW3, PEGB6, -, NW3
			10'd43 : rdata = 48'b000100100000001111100001100000000100110000000000;
			// PEs: 24, 29 -> 
			// srcs: (1835, 34)(3140) 47, (325) -2 --> (3462) -94:PEGB0, ND11, *, 
			10'd44 : rdata = 48'b000111110000000001100001011000000000000000000000;
			// PEs: 29, 29 -> 
			// srcs: (1838, 48)(3) 1, (3462) -94 --> (4246) -94:NM0, ALU, *, 
			10'd45 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 29, 29 -> 29
			// srcs: (1841, 63)(1110) -2, (4246) -94 --> (5030) 92:NW11, ALU, -, NW11
			10'd46 : rdata = 48'b000100100000101100111111111000000110110000000000;
			// PEs: 24, 29 -> 30
			// srcs: (1871, 35)(3140) 47, (361) -3 --> (3498) -141:PEGB0, ND4, *, PENB
			10'd47 : rdata = 48'b000111110000000001100000100000000000000100000000;
			// PEs: 29, 28 -> 28
			// srcs: (1873, 49)(3) 1, (3497) -47 --> (4281) -47:NM0, PENB, *, PEGB4
			10'd48 : rdata = 48'b000111000000000011011111110000000000000011000000;
			// PEs: 29, 30 -> 29
			// srcs: (1880, 64)(1146) 1, (4282) -141 --> (5066) 142:NW4, PEGB6, -, NW4
			10'd49 : rdata = 48'b000100100000010011100001100000000101000000000000;
			// PEs: 24, 29 -> 29
			// srcs: (1953, 36)(3140) 47, (443) 2 --> (3580) 94:PEGB0, ND5, *, NI0
			10'd50 : rdata = 48'b000111110000000001100000101100000000000000000000;
			// PEs: 29, 28 -> 28
			// srcs: (1955, 50)(3) 1, (3579) 94 --> (4363) 94:NM0, PENB, *, PEGB4
			10'd51 : rdata = 48'b000111000000000011011111110000000000000011000000;
			// PEs: 29, 29 -> 
			// srcs: (1956, 51)(3) 1, (3580) 94 --> (4364) 94:NM0, NI0, *, 
			10'd52 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 29, 29 -> 29
			// srcs: (1959, 65)(1228) -2, (4364) 94 --> (5148) -96:NW5, ALU, -, NW5
			10'd53 : rdata = 48'b000100100000010100111111111000000101010000000000;
			// PEs: 24, 29 -> 
			// srcs: (2019, 37)(3140) 47, (509) 2 --> (3646) 94:PEGB0, ND12, *, 
			10'd54 : rdata = 48'b000111110000000001100001100000000000000000000000;
			// PEs: 29, 29 -> 
			// srcs: (2022, 52)(3) 1, (3646) 94 --> (4430) 94:NM0, ALU, *, 
			10'd55 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 29, 29 -> 29
			// srcs: (2025, 66)(1294) -2, (4430) 94 --> (5214) -96:NW12, ALU, -, NW12
			10'd56 : rdata = 48'b000100100000110000111111111000000111000000000000;
			// PEs: 24, 29 -> 
			// srcs: (2033, 38)(3140) 47, (523) -1 --> (3660) -47:PEGB0, ND6, *, 
			10'd57 : rdata = 48'b000111110000000001100000110000000000000000000000;
			// PEs: 29, 29 -> 
			// srcs: (2036, 53)(3) 1, (3660) -47 --> (4444) -47:NM0, ALU, *, 
			10'd58 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 29, 29 -> 29
			// srcs: (2039, 67)(1308) 0, (4444) -47 --> (5228) 47:NW6, ALU, -, NW6
			10'd59 : rdata = 48'b000100100000011000111111111000000101100000000000;
			// PEs: 24, 29 -> 
			// srcs: (2113, 39)(3140) 47, (603) 0 --> (3740) 0:PEGB0, ND7, *, 
			10'd60 : rdata = 48'b000111110000000001100000111000000000000000000000;
			// PEs: 29, 29 -> 
			// srcs: (2116, 54)(3) 1, (3740) 0 --> (4524) 0:NM0, ALU, *, 
			10'd61 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 29, 29 -> 29
			// srcs: (2119, 68)(1388) 2, (4524) 0 --> (5308) 2:NW7, ALU, -, NW7
			10'd62 : rdata = 48'b000100100000011100111111111000000101110000000000;
			// PEs: 24, 29 -> 30
			// srcs: (2195, 40)(3140) 47, (685) 2 --> (3822) 94:PEGB0, ND8, *, PENB
			10'd63 : rdata = 48'b000111110000000001100001000000000000000100000000;
			// PEs: 29, 28 -> 28
			// srcs: (2197, 55)(3) 1, (3821) -47 --> (4605) -47:NM0, PENB, *, PEGB4
			10'd64 : rdata = 48'b000111000000000011011111110000000000000011000000;
			// PEs: 24, 29 -> 
			// srcs: (2199, 41)(3140) 47, (689) 2 --> (3826) 94:PEGB0, ND13, *, 
			10'd65 : rdata = 48'b000111110000000001100001101000000000000000000000;
			// PEs: 29, 29 -> 29
			// srcs: (2202, 56)(3) 1, (3826) 94 --> (4610) 94:NM0, ALU, *, NI0
			10'd66 : rdata = 48'b000111000000000000111111111100000000000000000000;
			// PEs: 29, 30 -> 29
			// srcs: (2204, 69)(1470) 2, (4606) 94 --> (5390) -92:NW8, PEGB6, -, NW8
			10'd67 : rdata = 48'b000100100000100011100001100000000110000000000000;
			// PEs: 29, 29 -> 29
			// srcs: (2205, 70)(1474) 1, (4610) 94 --> (5394) -93:NW13, NI0, -, NW13
			10'd68 : rdata = 48'b000100100000110110100000000000000111010000000000;
			// PEs: 24, 29 -> 30
			// srcs: (2275, 42)(3140) 47, (765) 0 --> (3902) 0:PEGB0, ND9, *, PENB
			10'd69 : rdata = 48'b000111110000000001100001001000000000000100000000;
			// PEs: 29, 28 -> 28
			// srcs: (2277, 57)(3) 1, (3901) -94 --> (4685) -94:NM0, PENB, *, PEGB4
			10'd70 : rdata = 48'b000111000000000011011111110000000000000011000000;
			// PEs: 29, 30 -> 29
			// srcs: (2284, 71)(1550) -3, (4686) 0 --> (5470) -3:NW9, PEGB6, -, NW9
			10'd71 : rdata = 48'b000100100000100111100001100000000110010000000000;
			default : rdata = 48'b000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 30) begin
	always @(*) begin
		case(address)
			// PEs: 30, 30 -> 24
			// srcs: (1, 0)(41) -3, (826) 2 --> (1610) -6:ND0, NW0, *, PEGB0
			10'd0 : rdata = 48'b000110110000000001000000000000000000000010000000;
			// PEs: 30, 30 -> 24
			// srcs: (2, 1)(121) -3, (906) -3 --> (1690) 9:ND1, NW1, *, PEGB0
			10'd1 : rdata = 48'b000110110000000101000000001000000000000010000000;
			// PEs: 30, 30 -> 30
			// srcs: (3, 2)(202) 1, (987) 1 --> (1771) 1:ND2, NW2, *, NI0
			10'd2 : rdata = 48'b000110110000001001000000010100000000000000000000;
			// PEs: 30, 30 -> 24
			// srcs: (4, 3)(283) 1, (1068) 2 --> (1852) 2:ND3, NW3, *, PEGB0
			10'd3 : rdata = 48'b000110110000001101000000011000000000000010000000;
			// PEs: 30, 30 -> 24
			// srcs: (5, 4)(363) 2, (1148) -2 --> (1932) -4:ND4, NW4, *, PEGB0
			10'd4 : rdata = 48'b000110110000010001000000100000000000000010000000;
			// PEs: 30, 30 -> 30
			// srcs: (6, 5)(445) 0, (1230) 0 --> (2014) 0:ND5, NW5, *, NI1
			10'd5 : rdata = 48'b000110110000010101000000101100001000000000000000;
			// PEs: 30, 30 -> 24
			// srcs: (7, 6)(525) 2, (1310) 2 --> (2094) 4:ND6, NW6, *, PEGB0
			10'd6 : rdata = 48'b000110110000011001000000110000000000000010000000;
			// PEs: 30, 30 -> 24
			// srcs: (8, 7)(605) -3, (1390) -1 --> (2174) 3:ND7, NW7, *, PEGB0
			10'd7 : rdata = 48'b000110110000011101000000111000000000000010000000;
			// PEs: 30, 30 -> 29
			// srcs: (9, 8)(687) 1, (1472) -3 --> (2256) -3:ND8, NW8, *, PEGB5
			10'd8 : rdata = 48'b000110110000100001000001000000000000000011010000;
			// PEs: 30, 30 -> 28
			// srcs: (10, 9)(767) -2, (1552) -2 --> (2336) 4:ND9, NW9, *, PEGB4
			10'd9 : rdata = 48'b000110110000100101000001001000000000000011000000;
			// PEs: 30, 30 -> 24
			// srcs: (11, 10)(144) -2, (929) 1 --> (1713) -2:ND10, NW10, *, PEGB0
			10'd10 : rdata = 48'b000110110000101001000001010000000000000010000000;
			// PEs: 30, 30 -> 30
			// srcs: (12, 11)(328) -2, (1113) 1 --> (1897) -2:ND11, NW11, *, NI2
			10'd11 : rdata = 48'b000110110000101101000001011100010000000000000000;
			// PEs: 30, 30 -> 30
			// srcs: (13, 12)(512) -2, (1297) -3 --> (2081) 6:ND12, NW12, *, NI3
			10'd12 : rdata = 48'b000110110000110001000001100100011000000000000000;
			// PEs: 30, 30 -> 30
			// srcs: (14, 13)(696) 2, (1481) 1 --> (2265) 2:ND13, NW13, *, NI4
			10'd13 : rdata = 48'b000110110000110101000001101100100000000000000000;
			// PEs: 28, 29 -> 28
			// srcs: (15, 18)(2253) 1, (2254) 4 --> (3031) 5:PEGB4, PENB, +, PEGB4
			10'd14 : rdata = 48'b000011110000100011011111110000000000000011000000;
			// PEs: 24 -> 
			// srcs: (27, 14)(1648) -6 --> (1648) -6:PEGB0, pass, 
			10'd15 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 24, 30 -> 25
			// srcs: (36, 15)(1647) 2, (1648) -6 --> (2429) -4:PEGB0, ALU, +, PEGB1
			10'd16 : rdata = 48'b000011110000000000111111111000000000000010010000;
			// PEs: 24 -> 
			// srcs: (66, 16)(1841) -1 --> (1841) -1:PEGB0, pass, 
			10'd17 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 24, 30 -> 24
			// srcs: (75, 17)(1840) -1, (1841) -1 --> (2619) -2:PEGB0, ALU, +, PEGB0
			10'd18 : rdata = 48'b000011110000000000111111111000000000000010000000;
			// PEs: 30 -> 24
			// srcs: (122, 19)(1771) 1 --> (1771) 1:NI0, pass, PEGB0
			10'd19 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 30 -> 24
			// srcs: (123, 21)(1897) -2 --> (1897) -2:NI2, pass, PEGB0
			10'd20 : rdata = 48'b110001010000001000000000000000000000000010000000;
			// PEs: 25, 30 -> 27
			// srcs: (131, 22)(2859) 0, (2081) 6 --> (2860) 6:PEGB1, NI3, +, PEGB3
			10'd21 : rdata = 48'b000011110000001010100000011000000000000010110000;
			// PEs: 30 -> 24
			// srcs: (137, 20)(2014) 0 --> (2014) 0:NI1, pass, PEGB0
			10'd22 : rdata = 48'b110001010000000100000000000000000000000010000000;
			// PEs: 25 -> 
			// srcs: (138, 23)(2862) 2 --> (2862) 2:PEGB1, pass, 
			10'd23 : rdata = 48'b110001110000001000000000000000000000000000000000;
			// PEs: 30, 31 -> 30
			// srcs: (141, 24)(2862) 2, (2084) -2 --> (2863) 0:ALU, PEGB7, +, NI0
			10'd24 : rdata = 48'b000010011111111111100001110100000000000000000000;
			// PEs: 27, 29 -> 31
			// srcs: (158, 27)(3030) -2, (3035) 6 --> (3036) 4:PEGB3, PENB, +, PENB
			10'd25 : rdata = 48'b000011110000011011011111110000000000000100000000;
			// PEs: 30 -> 24
			// srcs: (190, 25)(2265) 2 --> (2265) 2:NI4, pass, PEGB0
			10'd26 : rdata = 48'b110001010000010000000000000000000000000010000000;
			// PEs: 30 -> 24
			// srcs: (616, 26)(2863) 0 --> (2863) 0:NI0, pass, PEGB0
			10'd27 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 24, 30 -> 31
			// srcs: (1551, 28)(3140) 47, (41) -3 --> (3178) -141:PEGB0, ND0, *, PENB
			10'd28 : rdata = 48'b000111110000000001100000000000000000000100000000;
			// PEs: 30, 29 -> 29
			// srcs: (1552, 42)(3) 1, (3176) -141 --> (3960) -141:NM0, PENB, *, PEGB5
			10'd29 : rdata = 48'b000111000000000011011111110000000000000011010000;
			// PEs: 30, 31 -> 30
			// srcs: (1560, 59)(826) 2, (3962) -141 --> (4746) 143:NW0, PEGB7, -, NW0
			10'd30 : rdata = 48'b000100100000000011100001110000000100000000000000;
			// PEs: 24, 30 -> 30
			// srcs: (1631, 29)(3140) 47, (121) -3 --> (3258) -141:PEGB0, ND1, *, NI0
			10'd31 : rdata = 48'b000111110000000001100000001100000000000000000000;
			// PEs: 30, 29 -> 29
			// srcs: (1632, 43)(3) 1, (3256) -141 --> (4040) -141:NM0, PENB, *, PEGB5
			10'd32 : rdata = 48'b000111000000000011011111110000000000000011010000;
			// PEs: 30, 30 -> 
			// srcs: (1634, 44)(3) 1, (3258) -141 --> (4042) -141:NM0, NI0, *, 
			10'd33 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 30, 30 -> 30
			// srcs: (1637, 60)(906) -3, (4042) -141 --> (4826) 138:NW1, ALU, -, NW1
			10'd34 : rdata = 48'b000100100000000100111111111000000100010000000000;
			// PEs: 24, 30 -> 
			// srcs: (1654, 30)(3140) 47, (144) -2 --> (3281) -94:PEGB0, ND10, *, 
			10'd35 : rdata = 48'b000111110000000001100001010000000000000000000000;
			// PEs: 30, 30 -> 
			// srcs: (1657, 45)(3) 1, (3281) -94 --> (4065) -94:NM0, ALU, *, 
			10'd36 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 30, 30 -> 30
			// srcs: (1660, 61)(929) 1, (4065) -94 --> (4849) 95:NW10, ALU, -, NW10
			10'd37 : rdata = 48'b000100100000101000111111111000000110100000000000;
			// PEs: 24, 30 -> 
			// srcs: (1712, 31)(3140) 47, (202) 1 --> (3339) 47:PEGB0, ND2, *, 
			10'd38 : rdata = 48'b000111110000000001100000010000000000000000000000;
			// PEs: 30, 30 -> 
			// srcs: (1715, 46)(3) 1, (3339) 47 --> (4123) 47:NM0, ALU, *, 
			10'd39 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 30, 30 -> 30
			// srcs: (1718, 62)(987) 1, (4123) 47 --> (4907) -46:NW2, ALU, -, NW2
			10'd40 : rdata = 48'b000100100000001000111111111000000100100000000000;
			// PEs: 24, 30 -> 31
			// srcs: (1793, 32)(3140) 47, (283) 1 --> (3420) 47:PEGB0, ND3, *, PENB
			10'd41 : rdata = 48'b000111110000000001100000011000000000000100000000;
			// PEs: 30, 29 -> 29
			// srcs: (1794, 47)(3) 1, (3418) -141 --> (4202) -141:NM0, PENB, *, PEGB5
			10'd42 : rdata = 48'b000111000000000011011111110000000000000011010000;
			// PEs: 30, 31 -> 30
			// srcs: (1802, 63)(1068) 2, (4204) 47 --> (4988) -45:NW3, PEGB7, -, NW3
			10'd43 : rdata = 48'b000100100000001111100001110000000100110000000000;
			// PEs: 24, 30 -> 
			// srcs: (1838, 33)(3140) 47, (328) -2 --> (3465) -94:PEGB0, ND11, *, 
			10'd44 : rdata = 48'b000111110000000001100001011000000000000000000000;
			// PEs: 30, 30 -> 
			// srcs: (1841, 48)(3) 1, (3465) -94 --> (4249) -94:NM0, ALU, *, 
			10'd45 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 30, 30 -> 30
			// srcs: (1844, 64)(1113) 1, (4249) -94 --> (5033) 95:NW11, ALU, -, NW11
			10'd46 : rdata = 48'b000100100000101100111111111000000110110000000000;
			// PEs: 24, 30 -> 30
			// srcs: (1873, 34)(3140) 47, (363) 2 --> (3500) 94:PEGB0, ND4, *, NI0
			10'd47 : rdata = 48'b000111110000000001100000100100000000000000000000;
			// PEs: 30, 29 -> 29
			// srcs: (1874, 49)(3) 1, (3498) -141 --> (4282) -141:NM0, PENB, *, PEGB5
			10'd48 : rdata = 48'b000111000000000011011111110000000000000011010000;
			// PEs: 30, 30 -> 
			// srcs: (1876, 50)(3) 1, (3500) 94 --> (4284) 94:NM0, NI0, *, 
			10'd49 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 30, 30 -> 30
			// srcs: (1879, 65)(1148) -2, (4284) 94 --> (5068) -96:NW4, ALU, -, NW4
			10'd50 : rdata = 48'b000100100000010000111111111000000101000000000000;
			// PEs: 24, 30 -> 
			// srcs: (1955, 35)(3140) 47, (445) 0 --> (3582) 0:PEGB0, ND5, *, 
			10'd51 : rdata = 48'b000111110000000001100000101000000000000000000000;
			// PEs: 30, 30 -> 
			// srcs: (1958, 51)(3) 1, (3582) 0 --> (4366) 0:NM0, ALU, *, 
			10'd52 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 30, 30 -> 30
			// srcs: (1961, 66)(1230) 0, (4366) 0 --> (5150) 0:NW5, ALU, -, NW5
			10'd53 : rdata = 48'b000100100000010100111111111000000101010000000000;
			// PEs: 24, 30 -> 
			// srcs: (2022, 36)(3140) 47, (512) -2 --> (3649) -94:PEGB0, ND12, *, 
			10'd54 : rdata = 48'b000111110000000001100001100000000000000000000000;
			// PEs: 30, 30 -> 
			// srcs: (2025, 52)(3) 1, (3649) -94 --> (4433) -94:NM0, ALU, *, 
			10'd55 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 30, 30 -> 30
			// srcs: (2028, 67)(1297) -3, (4433) -94 --> (5217) 91:NW12, ALU, -, NW12
			10'd56 : rdata = 48'b000100100000110000111111111000000111000000000000;
			// PEs: 24, 30 -> 
			// srcs: (2035, 37)(3140) 47, (525) 2 --> (3662) 94:PEGB0, ND6, *, 
			10'd57 : rdata = 48'b000111110000000001100000110000000000000000000000;
			// PEs: 30, 30 -> 
			// srcs: (2038, 53)(3) 1, (3662) 94 --> (4446) 94:NM0, ALU, *, 
			10'd58 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 30, 30 -> 30
			// srcs: (2041, 68)(1310) 2, (4446) 94 --> (5230) -92:NW6, ALU, -, NW6
			10'd59 : rdata = 48'b000100100000011000111111111000000101100000000000;
			// PEs: 24, 30 -> 
			// srcs: (2115, 38)(3140) 47, (605) -3 --> (3742) -141:PEGB0, ND7, *, 
			10'd60 : rdata = 48'b000111110000000001100000111000000000000000000000;
			// PEs: 30, 30 -> 
			// srcs: (2118, 54)(3) 1, (3742) -141 --> (4526) -141:NM0, ALU, *, 
			10'd61 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 30, 30 -> 30
			// srcs: (2121, 69)(1390) -1, (4526) -141 --> (5310) 140:NW7, ALU, -, NW7
			10'd62 : rdata = 48'b000100100000011100111111111000000101110000000000;
			// PEs: 24, 30 -> 31
			// srcs: (2197, 39)(3140) 47, (687) 1 --> (3824) 47:PEGB0, ND8, *, PENB
			10'd63 : rdata = 48'b000111110000000001100001000000000000000100000000;
			// PEs: 30, 29 -> 29
			// srcs: (2198, 55)(3) 1, (3822) 94 --> (4606) 94:NM0, PENB, *, PEGB5
			10'd64 : rdata = 48'b000111000000000011011111110000000000000011010000;
			// PEs: 24, 30 -> 30
			// srcs: (2206, 40)(3140) 47, (696) 2 --> (3833) 94:PEGB0, ND13, *, NI0
			10'd65 : rdata = 48'b000111110000000001100001101100000000000000000000;
			// PEs: 30, 31 -> 30
			// srcs: (2207, 70)(1472) -3, (4608) 47 --> (5392) -50:NW8, PEGB7, -, NW8
			10'd66 : rdata = 48'b000100100000100011100001110000000110000000000000;
			// PEs: 30, 30 -> 
			// srcs: (2209, 56)(3) 1, (3833) 94 --> (4617) 94:NM0, NI0, *, 
			10'd67 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 30, 30 -> 30
			// srcs: (2212, 71)(1481) 1, (4617) 94 --> (5401) -93:NW13, ALU, -, NW13
			10'd68 : rdata = 48'b000100100000110100111111111000000111010000000000;
			// PEs: 24, 30 -> 30
			// srcs: (2277, 41)(3140) 47, (767) -2 --> (3904) -94:PEGB0, ND9, *, NI0
			10'd69 : rdata = 48'b000111110000000001100001001100000000000000000000;
			// PEs: 30, 29 -> 29
			// srcs: (2278, 57)(3) 1, (3902) 0 --> (4686) 0:NM0, PENB, *, PEGB5
			10'd70 : rdata = 48'b000111000000000011011111110000000000000011010000;
			// PEs: 30, 30 -> 
			// srcs: (2280, 58)(3) 1, (3904) -94 --> (4688) -94:NM0, NI0, *, 
			10'd71 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 30, 30 -> 30
			// srcs: (2283, 72)(1552) -2, (4688) -94 --> (5472) 92:NW9, ALU, -, NW9
			10'd72 : rdata = 48'b000100100000100100111111111000000110010000000000;
			default : rdata = 48'b000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 31) begin
	always @(*) begin
		case(address)
			// PEs: 31, 31 -> 24
			// srcs: (1, 0)(42) 2, (827) -1 --> (1611) -2:ND0, NW0, *, PENB
			10'd0 : rdata = 48'b000110110000000001000000000000000000000100000000;
			// PEs: 31, 31 -> 24
			// srcs: (2, 1)(122) -3, (907) -2 --> (1691) 6:ND1, NW1, *, PENB
			10'd1 : rdata = 48'b000110110000000101000000001000000000000100000000;
			// PEs: 31, 31 -> 31
			// srcs: (3, 2)(203) 0, (988) -1 --> (1772) 0:ND2, NW2, *, NI0
			10'd2 : rdata = 48'b000110110000001001000000010100000000000000000000;
			// PEs: 31, 31 -> 24
			// srcs: (4, 3)(284) -2, (1069) 1 --> (1853) -2:ND3, NW3, *, PENB
			10'd3 : rdata = 48'b000110110000001101000000011000000000000100000000;
			// PEs: 31, 31 -> 24
			// srcs: (5, 4)(364) 2, (1149) 0 --> (1933) 0:ND4, NW4, *, PENB
			10'd4 : rdata = 48'b000110110000010001000000100000000000000100000000;
			// PEs: 31, 31 -> 31
			// srcs: (6, 5)(446) 2, (1231) 2 --> (2015) 4:ND5, NW5, *, NI1
			10'd5 : rdata = 48'b000110110000010101000000101100001000000000000000;
			// PEs: 31, 31 -> 24
			// srcs: (7, 6)(526) -1, (1311) 0 --> (2095) 0:ND6, NW6, *, PENB
			10'd6 : rdata = 48'b000110110000011001000000110000000000000100000000;
			// PEs: 31, 31 -> 24
			// srcs: (8, 7)(606) -3, (1391) -2 --> (2175) 6:ND7, NW7, *, PENB
			10'd7 : rdata = 48'b000110110000011101000000111000000000000100000000;
			// PEs: 31, 31 -> 29
			// srcs: (9, 8)(688) -1, (1473) -2 --> (2257) 2:ND8, NW8, *, PEGB5
			10'd8 : rdata = 48'b000110110000100001000001000000000000000011010000;
			// PEs: 31, 31 -> 28
			// srcs: (10, 9)(768) 0, (1553) -3 --> (2337) 0:ND9, NW9, *, PEGB4
			10'd9 : rdata = 48'b000110110000100101000001001000000000000011000000;
			// PEs: 31, 31 -> 31
			// srcs: (11, 10)(147) 2, (932) -1 --> (1716) -2:ND10, NW10, *, NI2
			10'd10 : rdata = 48'b000110110000101001000001010100010000000000000000;
			// PEs: 31, 31 -> 31
			// srcs: (12, 11)(331) 0, (1116) -1 --> (1900) 0:ND11, NW11, *, NI3
			10'd11 : rdata = 48'b000110110000101101000001011100011000000000000000;
			// PEs: 31, 31 -> 30
			// srcs: (13, 12)(515) 1, (1300) -2 --> (2084) -2:ND12, NW12, *, PEGB6
			10'd12 : rdata = 48'b000110110000110001000001100000000000000011100000;
			// PEs: 31, 31 -> 31
			// srcs: (14, 13)(699) 1, (1484) 1 --> (2268) 1:ND13, NW13, *, NI4
			10'd13 : rdata = 48'b000110110000110101000001101100100000000000000000;
			// PEs: 27 -> 
			// srcs: (15, 18)(2331) 0 --> (2331) 0:PEGB3, pass, 
			10'd14 : rdata = 48'b110001110000011000000000000000000000000000000000;
			// PEs: 26, 31 -> 31
			// srcs: (18, 19)(2330) -6, (2331) 0 --> (3107) -6:PEGB2, ALU, +, NI5
			10'd15 : rdata = 48'b000011110000010000111111111100101000000000000000;
			// PEs: 24 -> 
			// srcs: (31, 14)(1651) -2 --> (1651) -2:PEGB0, pass, 
			10'd16 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 24, 31 -> 24
			// srcs: (40, 15)(1650) 9, (1651) -2 --> (2431) 7:PEGB0, ALU, +, PENB
			10'd17 : rdata = 48'b000011110000000000111111111000000000000100000000;
			// PEs: 24 -> 
			// srcs: (83, 16)(1923) -6 --> (1923) -6:PEGB0, pass, 
			10'd18 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 31, 25 -> 31
			// srcs: (85, 17)(1923) -6, (1924) -2 --> (2703) -8:ALU, PEGB1, +, NI6
			10'd19 : rdata = 48'b000010011111111111100000010100110000000000000000;
			// PEs: 31 -> 24
			// srcs: (120, 22)(1716) -2 --> (1716) -2:NI2, pass, PENB
			10'd20 : rdata = 48'b110001010000001000000000000000000000000100000000;
			// PEs: 31 -> 24
			// srcs: (130, 20)(1772) 0 --> (1772) 0:NI0, pass, PENB
			10'd21 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 31 -> 24
			// srcs: (146, 21)(2015) 4 --> (2015) 4:NI1, pass, PENB
			10'd22 : rdata = 48'b110001010000000100000000000000000000000100000000;
			// PEs: 31 -> 24
			// srcs: (152, 23)(1900) 0 --> (1900) 0:NI3, pass, PENB
			10'd23 : rdata = 48'b110001010000001100000000000000000000000100000000;
			// PEs: 31 -> 24
			// srcs: (170, 25)(2268) 1 --> (2268) 1:NI4, pass, PENB
			10'd24 : rdata = 48'b110001010000010000000000000000000000000100000000;
			// PEs: 31 -> 24
			// srcs: (176, 24)(2703) -8 --> (2703) -8:NI6, pass, PENB
			10'd25 : rdata = 48'b110001010000011000000000000000000000000100000000;
			// PEs: 31 -> 24
			// srcs: (177, 26)(3107) -6 --> (3107) -6:NI5, pass, PENB
			10'd26 : rdata = 48'b110001010000010100000000000000000000000100000000;
			// PEs: 28, 30 -> 24
			// srcs: (803, 27)(3025) -13, (3036) 4 --> (3037) -9:PEGB4, PENB, +, PENB
			10'd27 : rdata = 48'b000011110000100011011111110000000000000100000000;
			// PEs: 24, 31 -> 31
			// srcs: (1552, 28)(3140) 47, (42) 2 --> (3179) 94:PEGB0, ND0, *, NI0
			10'd28 : rdata = 48'b000111110000000001100000000100000000000000000000;
			// PEs: 31, 30 -> 30
			// srcs: (1554, 42)(3) 1, (3178) -141 --> (3962) -141:NM0, PENB, *, PEGB6
			10'd29 : rdata = 48'b000111000000000011011111110000000000000011100000;
			// PEs: 31, 31 -> 
			// srcs: (1555, 43)(3) 1, (3179) 94 --> (3963) 94:NM0, NI0, *, 
			10'd30 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 31, 31 -> 31
			// srcs: (1558, 59)(827) -1, (3963) 94 --> (4747) -95:NW0, ALU, -, NW0
			10'd31 : rdata = 48'b000100100000000000111111111000000100000000000000;
			// PEs: 24, 31 -> 
			// srcs: (1632, 29)(3140) 47, (122) -3 --> (3259) -141:PEGB0, ND1, *, 
			10'd32 : rdata = 48'b000111110000000001100000001000000000000000000000;
			// PEs: 31, 31 -> 
			// srcs: (1635, 44)(3) 1, (3259) -141 --> (4043) -141:NM0, ALU, *, 
			10'd33 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 31, 31 -> 31
			// srcs: (1638, 60)(907) -2, (4043) -141 --> (4827) 139:NW1, ALU, -, NW1
			10'd34 : rdata = 48'b000100100000000100111111111000000100010000000000;
			// PEs: 24, 31 -> 
			// srcs: (1657, 30)(3140) 47, (147) 2 --> (3284) 94:PEGB0, ND10, *, 
			10'd35 : rdata = 48'b000111110000000001100001010000000000000000000000;
			// PEs: 31, 31 -> 
			// srcs: (1660, 45)(3) 1, (3284) 94 --> (4068) 94:NM0, ALU, *, 
			10'd36 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 31, 31 -> 31
			// srcs: (1663, 61)(932) -1, (4068) 94 --> (4852) -95:NW10, ALU, -, NW10
			10'd37 : rdata = 48'b000100100000101000111111111000000110100000000000;
			// PEs: 24, 31 -> 
			// srcs: (1713, 31)(3140) 47, (203) 0 --> (3340) 0:PEGB0, ND2, *, 
			10'd38 : rdata = 48'b000111110000000001100000010000000000000000000000;
			// PEs: 31, 31 -> 
			// srcs: (1716, 46)(3) 1, (3340) 0 --> (4124) 0:NM0, ALU, *, 
			10'd39 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 31, 31 -> 31
			// srcs: (1719, 62)(988) -1, (4124) 0 --> (4908) -1:NW2, ALU, -, NW2
			10'd40 : rdata = 48'b000100100000001000111111111000000100100000000000;
			// PEs: 24, 31 -> 31
			// srcs: (1794, 32)(3140) 47, (284) -2 --> (3421) -94:PEGB0, ND3, *, NI0
			10'd41 : rdata = 48'b000111110000000001100000011100000000000000000000;
			// PEs: 31, 30 -> 30
			// srcs: (1796, 47)(3) 1, (3420) 47 --> (4204) 47:NM0, PENB, *, PEGB6
			10'd42 : rdata = 48'b000111000000000011011111110000000000000011100000;
			// PEs: 31, 31 -> 
			// srcs: (1797, 48)(3) 1, (3421) -94 --> (4205) -94:NM0, NI0, *, 
			10'd43 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 31, 31 -> 31
			// srcs: (1800, 63)(1069) 1, (4205) -94 --> (4989) 95:NW3, ALU, -, NW3
			10'd44 : rdata = 48'b000100100000001100111111111000000100110000000000;
			// PEs: 24, 31 -> 
			// srcs: (1841, 33)(3140) 47, (331) 0 --> (3468) 0:PEGB0, ND11, *, 
			10'd45 : rdata = 48'b000111110000000001100001011000000000000000000000;
			// PEs: 31, 31 -> 
			// srcs: (1844, 49)(3) 1, (3468) 0 --> (4252) 0:NM0, ALU, *, 
			10'd46 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 31, 31 -> 31
			// srcs: (1847, 64)(1116) -1, (4252) 0 --> (5036) -1:NW11, ALU, -, NW11
			10'd47 : rdata = 48'b000100100000101100111111111000000110110000000000;
			// PEs: 24, 31 -> 
			// srcs: (1874, 34)(3140) 47, (364) 2 --> (3501) 94:PEGB0, ND4, *, 
			10'd48 : rdata = 48'b000111110000000001100000100000000000000000000000;
			// PEs: 31, 31 -> 
			// srcs: (1877, 50)(3) 1, (3501) 94 --> (4285) 94:NM0, ALU, *, 
			10'd49 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 31, 31 -> 31
			// srcs: (1880, 65)(1149) 0, (4285) 94 --> (5069) -94:NW4, ALU, -, NW4
			10'd50 : rdata = 48'b000100100000010000111111111000000101000000000000;
			// PEs: 24, 31 -> 
			// srcs: (1956, 35)(3140) 47, (446) 2 --> (3583) 94:PEGB0, ND5, *, 
			10'd51 : rdata = 48'b000111110000000001100000101000000000000000000000;
			// PEs: 31, 31 -> 
			// srcs: (1959, 51)(3) 1, (3583) 94 --> (4367) 94:NM0, ALU, *, 
			10'd52 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 31, 31 -> 31
			// srcs: (1962, 66)(1231) 2, (4367) 94 --> (5151) -92:NW5, ALU, -, NW5
			10'd53 : rdata = 48'b000100100000010100111111111000000101010000000000;
			// PEs: 24, 31 -> 
			// srcs: (2025, 36)(3140) 47, (515) 1 --> (3652) 47:PEGB0, ND12, *, 
			10'd54 : rdata = 48'b000111110000000001100001100000000000000000000000;
			// PEs: 31, 31 -> 
			// srcs: (2028, 52)(3) 1, (3652) 47 --> (4436) 47:NM0, ALU, *, 
			10'd55 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 31, 31 -> 31
			// srcs: (2031, 67)(1300) -2, (4436) 47 --> (5220) -49:NW12, ALU, -, NW12
			10'd56 : rdata = 48'b000100100000110000111111111000000111000000000000;
			// PEs: 24, 31 -> 
			// srcs: (2036, 37)(3140) 47, (526) -1 --> (3663) -47:PEGB0, ND6, *, 
			10'd57 : rdata = 48'b000111110000000001100000110000000000000000000000;
			// PEs: 31, 31 -> 
			// srcs: (2039, 53)(3) 1, (3663) -47 --> (4447) -47:NM0, ALU, *, 
			10'd58 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 31, 31 -> 31
			// srcs: (2042, 68)(1311) 0, (4447) -47 --> (5231) 47:NW6, ALU, -, NW6
			10'd59 : rdata = 48'b000100100000011000111111111000000101100000000000;
			// PEs: 24, 31 -> 
			// srcs: (2116, 38)(3140) 47, (606) -3 --> (3743) -141:PEGB0, ND7, *, 
			10'd60 : rdata = 48'b000111110000000001100000111000000000000000000000;
			// PEs: 31, 31 -> 
			// srcs: (2119, 54)(3) 1, (3743) -141 --> (4527) -141:NM0, ALU, *, 
			10'd61 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 31, 31 -> 31
			// srcs: (2122, 69)(1391) -2, (4527) -141 --> (5311) 139:NW7, ALU, -, NW7
			10'd62 : rdata = 48'b000100100000011100111111111000000101110000000000;
			// PEs: 24, 31 -> 31
			// srcs: (2198, 39)(3140) 47, (688) -1 --> (3825) -47:PEGB0, ND8, *, NI0
			10'd63 : rdata = 48'b000111110000000001100001000100000000000000000000;
			// PEs: 31, 30 -> 30
			// srcs: (2200, 55)(3) 1, (3824) 47 --> (4608) 47:NM0, PENB, *, PEGB6
			10'd64 : rdata = 48'b000111000000000011011111110000000000000011100000;
			// PEs: 31, 31 -> 
			// srcs: (2201, 56)(3) 1, (3825) -47 --> (4609) -47:NM0, NI0, *, 
			10'd65 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 31, 31 -> 31
			// srcs: (2204, 70)(1473) -2, (4609) -47 --> (5393) 45:NW8, ALU, -, NW8
			10'd66 : rdata = 48'b000100100000100000111111111000000110000000000000;
			// PEs: 24, 31 -> 
			// srcs: (2209, 40)(3140) 47, (699) 1 --> (3836) 47:PEGB0, ND13, *, 
			10'd67 : rdata = 48'b000111110000000001100001101000000000000000000000;
			// PEs: 31, 31 -> 
			// srcs: (2212, 57)(3) 1, (3836) 47 --> (4620) 47:NM0, ALU, *, 
			10'd68 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 31, 31 -> 31
			// srcs: (2215, 71)(1484) 1, (4620) 47 --> (5404) -46:NW13, ALU, -, NW13
			10'd69 : rdata = 48'b000100100000110100111111111000000111010000000000;
			// PEs: 24, 31 -> 
			// srcs: (2278, 41)(3140) 47, (768) 0 --> (3905) 0:PEGB0, ND9, *, 
			10'd70 : rdata = 48'b000111110000000001100001001000000000000000000000;
			// PEs: 31, 31 -> 
			// srcs: (2281, 58)(3) 1, (3905) 0 --> (4689) 0:NM0, ALU, *, 
			10'd71 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 31, 31 -> 31
			// srcs: (2284, 72)(1553) -3, (4689) 0 --> (5473) -3:NW9, ALU, -, NW9
			10'd72 : rdata = 48'b000100100000100100111111111000000110010000000000;
			default : rdata = 48'b000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 32) begin
	always @(*) begin
		case(address)
			// PEs: 39 -> 56
			// srcs: (3, 124)(1622) -6 --> (1622) -6:PENB, pass, PUGB7
			10'd0 : rdata = 48'b110001101111111000000000000000000000000000001111;
			// PEs: 39 -> 48
			// srcs: (4, 27)(1702) -4 --> (1702) -4:PENB, pass, PUGB6
			10'd1 : rdata = 48'b110001101111111000000000000000000000000000001110;
			// PEs: 39 -> 48
			// srcs: (5, 40)(1782) 3 --> (1782) 3:PENB, pass, PUGB6
			10'd2 : rdata = 48'b110001101111111000000000000000000000000000001110;
			// PEs: 33 -> 8
			// srcs: (6, 0)(1613) 0 --> (1613) 0:PEGB1, pass, PUGB1
			10'd3 : rdata = 48'b110001110000001000000000000000000000000000001001;
			// PEs: 34 -> 8
			// srcs: (7, 1)(1614) 6 --> (1614) 6:PEGB2, pass, PUGB1
			10'd4 : rdata = 48'b110001110000010000000000000000000000000000001001;
			// PEs: 35 -> 16
			// srcs: (8, 2)(1616) 0 --> (1616) 0:PEGB3, pass, PUGB2
			10'd5 : rdata = 48'b110001110000011000000000000000000000000000001010;
			// PEs: 36 -> 16
			// srcs: (9, 3)(1617) -4 --> (1617) -4:PEGB4, pass, PUGB2
			10'd6 : rdata = 48'b110001110000100000000000000000000000000000001010;
			// PEs: 37 -> 16
			// srcs: (10, 4)(1619) 0 --> (1619) 0:PEGB5, pass, PUGB2
			10'd7 : rdata = 48'b110001110000101000000000000000000000000000001010;
			// PEs: 38 -> 16
			// srcs: (11, 5)(1620) 0 --> (1620) 0:PEGB6, pass, PUGB2
			10'd8 : rdata = 48'b110001110000110000000000000000000000000000001010;
			// PEs: 33 -> 40
			// srcs: (12, 21)(1693) 0 --> (1693) 0:PEGB1, pass, PUNB
			10'd9 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 34 -> 40
			// srcs: (13, 22)(1694) -6 --> (1694) -6:PEGB2, pass, PUNB
			10'd10 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 35 -> 40
			// srcs: (14, 23)(1696) 2 --> (1696) 2:PEGB3, pass, PUNB
			10'd11 : rdata = 48'b110001110000011000000000000000000000001000000000;
			// PEs: 36 -> 40
			// srcs: (15, 24)(1697) 2 --> (1697) 2:PEGB4, pass, PUNB
			10'd12 : rdata = 48'b110001110000100000000000000000000000001000000000;
			// PEs: 37 -> 40
			// srcs: (16, 25)(1699) 0 --> (1699) 0:PEGB5, pass, PUNB
			10'd13 : rdata = 48'b110001110000101000000000000000000000001000000000;
			// PEs: 38 -> 40
			// srcs: (17, 26)(1700) -2 --> (1700) -2:PEGB6, pass, PUNB
			10'd14 : rdata = 48'b110001110000110000000000000000000000001000000000;
			// PEs: 33 -> 40
			// srcs: (18, 34)(1773) 0 --> (1773) 0:PEGB1, pass, PUNB
			10'd15 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 34 -> 40
			// srcs: (19, 35)(1774) 1 --> (1774) 1:PEGB2, pass, PUNB
			10'd16 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 35 -> 40
			// srcs: (20, 36)(1776) 9 --> (1776) 9:PEGB3, pass, PUNB
			10'd17 : rdata = 48'b110001110000011000000000000000000000001000000000;
			// PEs: 36 -> 40
			// srcs: (21, 37)(1777) 2 --> (1777) 2:PEGB4, pass, PUNB
			10'd18 : rdata = 48'b110001110000100000000000000000000000001000000000;
			// PEs: 37 -> 40
			// srcs: (22, 38)(1779) 0 --> (1779) 0:PEGB5, pass, PUNB
			10'd19 : rdata = 48'b110001110000101000000000000000000000001000000000;
			// PEs: 38 -> 40
			// srcs: (23, 39)(1780) -6 --> (1780) -6:PEGB6, pass, PUNB
			10'd20 : rdata = 48'b110001110000110000000000000000000000001000000000;
			// PEs: 33 -> 40
			// srcs: (24, 56)(1855) 4 --> (1855) 4:PEGB1, pass, PUNB
			10'd21 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 34 -> 40
			// srcs: (25, 57)(1856) 0 --> (1856) 0:PEGB2, pass, PUNB
			10'd22 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 35 -> 40
			// srcs: (26, 58)(1858) 2 --> (1858) 2:PEGB3, pass, PUNB
			10'd23 : rdata = 48'b110001110000011000000000000000000000001000000000;
			// PEs: 36 -> 40
			// srcs: (27, 59)(1859) -4 --> (1859) -4:PEGB4, pass, PUNB
			10'd24 : rdata = 48'b110001110000100000000000000000000000001000000000;
			// PEs: 37 -> 40
			// srcs: (28, 60)(1861) 1 --> (1861) 1:PEGB5, pass, PUNB
			10'd25 : rdata = 48'b110001110000101000000000000000000000001000000000;
			// PEs: 38 -> 40
			// srcs: (29, 61)(1862) 0 --> (1862) 0:PEGB6, pass, PUNB
			10'd26 : rdata = 48'b110001110000110000000000000000000000001000000000;
			// PEs: 0 -> 32
			// srcs: (30, 6)(1659) 2 --> (1659) 2:PUGB0, pass, NI0
			10'd27 : rdata = 48'b110001110000000100000000000100000000000000000000;
			// PEs: 39 -> 48
			// srcs: (31, 62)(1864) 1 --> (1864) 1:PENB, pass, PUGB6
			10'd28 : rdata = 48'b110001101111111000000000000000000000000000001110;
			// PEs: 0 -> 33
			// srcs: (32, 7)(1660) 0 --> (1660) 0:PUGB0, pass, PENB
			10'd29 : rdata = 48'b110001110000000100000000000000000000000100000000;
			// PEs: 33 -> 40
			// srcs: (33, 72)(1935) 4 --> (1935) 4:PEGB1, pass, PUNB
			10'd30 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 24 -> 32
			// srcs: (34, 10)(1682) -2 --> (1682) -2:PUNB, pass, NI1
			10'd31 : rdata = 48'b110001101111111100000000000100001000000000000000;
			// PEs: 24 -> 32
			// srcs: (35, 12)(1684) 1 --> (1684) 1:PUNB, pass, NI2
			10'd32 : rdata = 48'b110001101111111100000000000100010000000000000000;
			// PEs: 24 -> 35
			// srcs: (36, 13)(1685) 0 --> (1685) 0:PUNB, pass, PEGB3
			10'd33 : rdata = 48'b110001101111111100000000000000000000000010110000;
			// PEs: 34 -> 40
			// srcs: (37, 73)(1936) -3 --> (1936) -3:PEGB2, pass, PUNB
			10'd34 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 32 -> 33
			// srcs: (38, 8)(1659) 2 --> (1659) 2:NI0, pass, PENB
			10'd35 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 24 -> 32
			// srcs: (39, 15)(1687) -2 --> (1687) -2:PUNB, pass, NI0
			10'd36 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 24 -> 36
			// srcs: (40, 16)(1688) -3 --> (1688) -3:PUNB, pass, PEGB4
			10'd37 : rdata = 48'b110001101111111100000000000000000000000011000000;
			// PEs: 24 -> 32
			// srcs: (41, 18)(1690) 9 --> (1690) 9:PUNB, pass, NI3
			10'd38 : rdata = 48'b110001101111111100000000000100011000000000000000;
			// PEs: 24 -> 37
			// srcs: (42, 19)(1691) 6 --> (1691) 6:PUNB, pass, PEGB5
			10'd39 : rdata = 48'b110001101111111100000000000000000000000011010000;
			// PEs: 16 -> 34
			// srcs: (43, 9)(1681) 3 --> (1681) 3:PUGB2, pass, PEGB2
			10'd40 : rdata = 48'b110001110000010100000000000000000000000010100000;
			// PEs: 24 -> 32
			// srcs: (44, 29)(1764) 0 --> (1764) 0:PUNB, pass, NI4
			10'd41 : rdata = 48'b110001101111111100000000000100100000000000000000;
			// PEs: 32 -> 35
			// srcs: (45, 14)(1684) 1 --> (1684) 1:NI2, pass, PEGB3
			10'd42 : rdata = 48'b110001010000001000000000000000000000000010110000;
			// PEs: 24 -> 32
			// srcs: (46, 31)(1766) -3 --> (1766) -3:PUNB, pass, NI2
			10'd43 : rdata = 48'b110001101111111100000000000100010000000000000000;
			// PEs: 56 -> 32
			// srcs: (47, 41)(1812) 3 --> (1812) 3:PUGB7, pass, NI5
			10'd44 : rdata = 48'b110001110000111100000000000100101000000000000000;
			// PEs: 56 -> 33
			// srcs: (48, 42)(1813) 2 --> (1813) 2:PUGB7, pass, PENB
			10'd45 : rdata = 48'b110001110000111100000000000000000000000100000000;
			// PEs: 32 -> 36
			// srcs: (49, 17)(1687) -2 --> (1687) -2:NI0, pass, PEGB4
			10'd46 : rdata = 48'b110001010000000000000000000000000000000011000000;
			// PEs: 16 -> 38
			// srcs: (50, 28)(1763) 0 --> (1763) 0:PUGB2, pass, PEGB6
			10'd47 : rdata = 48'b110001110000010100000000000000000000000011100000;
			// PEs: 32 -> 37
			// srcs: (51, 20)(1690) 9 --> (1690) 9:NI3, pass, PEGB5
			10'd48 : rdata = 48'b110001010000001100000000000000000000000011010000;
			// PEs: 32 -> 34
			// srcs: (52, 11)(1682) -2 --> (1682) -2:NI1, pass, PEGB2
			10'd49 : rdata = 48'b110001010000000100000000000000000000000010100000;
			// PEs: 24 -> 39
			// srcs: (53, 32)(1767) 0 --> (1767) 0:PUNB, pass, PEGB7
			10'd50 : rdata = 48'b110001101111111100000000000000000000000011110000;
			// PEs: 32 -> 33
			// srcs: (54, 43)(1812) 3 --> (1812) 3:NI5, pass, PENB
			10'd51 : rdata = 48'b110001010000010100000000000000000000000100000000;
			// PEs: 35 -> 40
			// srcs: (55, 74)(1938) -2 --> (1938) -2:PEGB3, pass, PUNB
			10'd52 : rdata = 48'b110001110000011000000000000000000000001000000000;
			// PEs: 36 -> 40
			// srcs: (56, 75)(1939) -1 --> (1939) -1:PEGB4, pass, PUNB
			10'd53 : rdata = 48'b110001110000100000000000000000000000001000000000;
			// PEs: 37 -> 40
			// srcs: (57, 76)(1941) 0 --> (1941) 0:PEGB5, pass, PUNB
			10'd54 : rdata = 48'b110001110000101000000000000000000000001000000000;
			// PEs: 38 -> 40
			// srcs: (58, 77)(1942) 2 --> (1942) 2:PEGB6, pass, PUNB
			10'd55 : rdata = 48'b110001110000110000000000000000000000001000000000;
			// PEs: 32 -> 38
			// srcs: (59, 30)(1764) 0 --> (1764) 0:NI4, pass, PEGB6
			10'd56 : rdata = 48'b110001010000010000000000000000000000000011100000;
			// PEs: 39 -> 40
			// srcs: (60, 78)(1944) 4 --> (1944) 4:PENB, pass, PUNB
			10'd57 : rdata = 48'b110001101111111000000000000000000000001000000000;
			// PEs: 35 -> 40
			// srcs: (61, 85)(2018) -2 --> (2018) -2:PEGB3, pass, PUNB
			10'd58 : rdata = 48'b110001110000011000000000000000000000001000000000;
			// PEs: 32 -> 39
			// srcs: (62, 33)(1766) -3 --> (1766) -3:NI2, pass, PEGB7
			10'd59 : rdata = 48'b110001010000001000000000000000000000000011110000;
			// PEs: 36 -> 40
			// srcs: (63, 86)(2019) 0 --> (2019) 0:PEGB4, pass, PUNB
			10'd60 : rdata = 48'b110001110000100000000000000000000000001000000000;
			// PEs: 16 -> 32
			// srcs: (64, 44)(1843) 1 --> (1843) 1:PUGB2, pass, NI0
			10'd61 : rdata = 48'b110001110000010100000000000100000000000000000000;
			// PEs: 24 -> 34
			// srcs: (65, 45)(1844) 9 --> (1844) 9:PUNB, pass, PEGB2
			10'd62 : rdata = 48'b110001101111111100000000000000000000000010100000;
			// PEs: 24 -> 32
			// srcs: (66, 47)(1846) 0 --> (1846) 0:PUNB, pass, NI1
			10'd63 : rdata = 48'b110001101111111100000000000100001000000000000000;
			// PEs: 24 -> 35
			// srcs: (67, 48)(1847) 0 --> (1847) 0:PUNB, pass, PEGB3
			10'd64 : rdata = 48'b110001101111111100000000000000000000000010110000;
			// PEs: 24 -> 32
			// srcs: (68, 50)(1849) 0 --> (1849) 0:PUNB, pass, NI2
			10'd65 : rdata = 48'b110001101111111100000000000100010000000000000000;
			// PEs: 24 -> 36
			// srcs: (69, 51)(1850) 3 --> (1850) 3:PUNB, pass, PEGB4
			10'd66 : rdata = 48'b110001101111111100000000000000000000000011000000;
			// PEs: 24 -> 32
			// srcs: (70, 53)(1852) 2 --> (1852) 2:PUNB, pass, NI3
			10'd67 : rdata = 48'b110001101111111100000000000100011000000000000000;
			// PEs: 24 -> 37
			// srcs: (71, 54)(1853) -2 --> (1853) -2:PUNB, pass, PEGB5
			10'd68 : rdata = 48'b110001101111111100000000000000000000000011010000;
			// PEs: 24 -> 32
			// srcs: (72, 63)(1926) -2 --> (1926) -2:PUNB, pass, NI4
			10'd69 : rdata = 48'b110001101111111100000000000100100000000000000000;
			// PEs: 24 -> 33
			// srcs: (73, 64)(1927) -2 --> (1927) -2:PUNB, pass, PENB
			10'd70 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 32 -> 34
			// srcs: (74, 46)(1843) 1 --> (1843) 1:NI0, pass, PEGB2
			10'd71 : rdata = 48'b110001010000000000000000000000000000000010100000;
			// PEs: 37 -> 40
			// srcs: (75, 87)(2021) 2 --> (2021) 2:PEGB5, pass, PUNB
			10'd72 : rdata = 48'b110001110000101000000000000000000000001000000000;
			// PEs: 32 -> 35
			// srcs: (76, 49)(1846) 0 --> (1846) 0:NI1, pass, PEGB3
			10'd73 : rdata = 48'b110001010000000100000000000000000000000010110000;
			// PEs: 38 -> 40
			// srcs: (77, 88)(2022) 0 --> (2022) 0:PEGB6, pass, PUNB
			10'd74 : rdata = 48'b110001110000110000000000000000000000001000000000;
			// PEs: 32 -> 36
			// srcs: (78, 52)(1849) 0 --> (1849) 0:NI2, pass, PEGB4
			10'd75 : rdata = 48'b110001010000001000000000000000000000000011000000;
			// PEs: 32 -> 33
			// srcs: (79, 65)(1926) -2 --> (1926) -2:NI4, pass, PENB
			10'd76 : rdata = 48'b110001010000010000000000000000000000000100000000;
			// PEs: 32 -> 37
			// srcs: (80, 55)(1852) 2 --> (1852) 2:NI3, pass, PEGB5
			10'd77 : rdata = 48'b110001010000001100000000000000000000000011010000;
			// PEs: 24 -> 32
			// srcs: (81, 66)(1929) 2 --> (1929) 2:PUNB, pass, NI0
			10'd78 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 24 -> 33
			// srcs: (82, 67)(1930) -3 --> (1930) -3:PUNB, pass, PENB
			10'd79 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 39 -> 40
			// srcs: (83, 89)(2024) 0 --> (2024) 0:PENB, pass, PUNB
			10'd80 : rdata = 48'b110001101111111000000000000000000000001000000000;
			// PEs: 33 -> 40
			// srcs: (84, 99)(2097) 6 --> (2097) 6:PEGB1, pass, PUNB
			10'd81 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 34 -> 40
			// srcs: (85, 100)(2098) 0 --> (2098) 0:PEGB2, pass, PUNB
			10'd82 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 35 -> 40
			// srcs: (86, 101)(2100) -3 --> (2100) -3:PEGB3, pass, PUNB
			10'd83 : rdata = 48'b110001110000011000000000000000000000001000000000;
			// PEs: 36 -> 40
			// srcs: (87, 102)(2101) 6 --> (2101) 6:PEGB4, pass, PUNB
			10'd84 : rdata = 48'b110001110000100000000000000000000000001000000000;
			// PEs: 32 -> 33
			// srcs: (88, 68)(1929) 2 --> (1929) 2:NI0, pass, PENB
			10'd85 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 24 -> 32
			// srcs: (89, 69)(1932) -4 --> (1932) -4:PUNB, pass, NI0
			10'd86 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 24 -> 33
			// srcs: (90, 70)(1933) 0 --> (1933) 0:PUNB, pass, PENB
			10'd87 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 37 -> 40
			// srcs: (91, 103)(2103) 0 --> (2103) 0:PEGB5, pass, PUNB
			10'd88 : rdata = 48'b110001110000101000000000000000000000001000000000;
			// PEs: 38 -> 40
			// srcs: (92, 104)(2104) 0 --> (2104) 0:PEGB6, pass, PUNB
			10'd89 : rdata = 48'b110001110000110000000000000000000000001000000000;
			// PEs: 39 -> 40
			// srcs: (93, 105)(2106) -6 --> (2106) -6:PENB, pass, PUNB
			10'd90 : rdata = 48'b110001101111111000000000000000000000001000000000;
			// PEs: 33 -> 40
			// srcs: (94, 115)(2177) 0 --> (2177) 0:PEGB1, pass, PUNB
			10'd91 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 34 -> 40
			// srcs: (95, 116)(2178) 3 --> (2178) 3:PEGB2, pass, PUNB
			10'd92 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 32 -> 33
			// srcs: (96, 71)(1932) -4 --> (1932) -4:NI0, pass, PENB
			10'd93 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 24 -> 32
			// srcs: (97, 79)(2008) 0 --> (2008) 0:PUNB, pass, NI0
			10'd94 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 24 -> 33
			// srcs: (98, 80)(2009) -3 --> (2009) -3:PUNB, pass, PENB
			10'd95 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 35 -> 40
			// srcs: (99, 117)(2180) 0 --> (2180) 0:PEGB3, pass, PUNB
			10'd96 : rdata = 48'b110001110000011000000000000000000000001000000000;
			// PEs: 36 -> 40
			// srcs: (100, 118)(2181) 2 --> (2181) 2:PEGB4, pass, PUNB
			10'd97 : rdata = 48'b110001110000100000000000000000000000001000000000;
			// PEs: 37 -> 40
			// srcs: (101, 119)(2183) -2 --> (2183) -2:PEGB5, pass, PUNB
			10'd98 : rdata = 48'b110001110000101000000000000000000000001000000000;
			// PEs: 38 -> 40
			// srcs: (102, 120)(2184) -3 --> (2184) -3:PEGB6, pass, PUNB
			10'd99 : rdata = 48'b110001110000110000000000000000000000001000000000;
			// PEs: 39 -> 40
			// srcs: (103, 121)(2186) 3 --> (2186) 3:PENB, pass, PUNB
			10'd100 : rdata = 48'b110001101111111000000000000000000000001000000000;
			// PEs: 32 -> 33
			// srcs: (104, 81)(2008) 0 --> (2008) 0:NI0, pass, PENB
			10'd101 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 24 -> 32
			// srcs: (105, 82)(2011) -6 --> (2011) -6:PUNB, pass, NI0
			10'd102 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 24 -> 33
			// srcs: (106, 83)(2012) -4 --> (2012) -4:PUNB, pass, PENB
			10'd103 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 39 -> 40
			// srcs: (107, 122)(2266) -3 --> (2266) -3:PENB, pass, PUNB
			10'd104 : rdata = 48'b110001101111111000000000000000000000001000000000;
			// PEs: 39 -> 40
			// srcs: (108, 123)(2348) -2 --> (2348) -2:PENB, pass, PUNB
			10'd105 : rdata = 48'b110001101111111000000000000000000000001000000000;
			// PEs: 33 -> 48
			// srcs: (109, 145)(2440) 2 --> (2440) 2:PEGB1, pass, PUGB6
			10'd106 : rdata = 48'b110001110000001000000000000000000000000000001110;
			// PEs: 34 -> 0
			// srcs: (110, 149)(2462) 1 --> (2462) 1:PEGB2, pass, PUGB0
			10'd107 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 35 -> 24
			// srcs: (111, 150)(2466) 1 --> (2466) 1:PEGB3, pass, PUGB3
			10'd108 : rdata = 48'b110001110000011000000000000000000000000000001011;
			// PEs: 32 -> 33
			// srcs: (112, 84)(2011) -6 --> (2011) -6:NI0, pass, PENB
			10'd109 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 24 -> 32
			// srcs: (113, 90)(2088) -2 --> (2088) -2:PUNB, pass, NI0
			10'd110 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 24 -> 33
			// srcs: (114, 91)(2089) 0 --> (2089) 0:PUNB, pass, PENB
			10'd111 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 36 -> 56
			// srcs: (115, 151)(2468) -5 --> (2468) -5:PEGB4, pass, PUGB7
			10'd112 : rdata = 48'b110001110000100000000000000000000000000000001111;
			// PEs: 33 -> 40
			// srcs: (116, 134)(2016) 1 --> (2016) 1:PEGB1, pass, PUNB
			10'd113 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 37 -> 8
			// srcs: (117, 152)(2471) 15 --> (2471) 15:PEGB5, pass, PUGB1
			10'd114 : rdata = 48'b110001110000101000000000000000000000000000001001;
			// PEs: 36 -> 0
			// srcs: (118, 174)(2629) 3 --> (2629) 3:PEGB4, pass, PUGB0
			10'd115 : rdata = 48'b110001110000100000000000000000000000000000001000;
			// PEs: 32 -> 33
			// srcs: (120, 92)(2088) -2 --> (2088) -2:NI0, pass, PENB
			10'd116 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 24 -> 32
			// srcs: (121, 93)(2091) 0 --> (2091) 0:PUNB, pass, NI0
			10'd117 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 24 -> 33
			// srcs: (122, 94)(2092) 0 --> (2092) 0:PUNB, pass, PENB
			10'd118 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 34 -> 40
			// srcs: (124, 135)(2017) 0 --> (2017) 0:PEGB2, pass, PUNB
			10'd119 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 33 -> 8
			// srcs: (125, 156)(1719) 6 --> (1719) 6:PEGB1, pass, PUGB1
			10'd120 : rdata = 48'b110001110000001000000000000000000000000000001001;
			// PEs: 34 -> 24
			// srcs: (126, 157)(1726) 6 --> (1726) 6:PEGB2, pass, PUGB3
			10'd121 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 35 -> 48
			// srcs: (127, 158)(1729) -3 --> (1729) -3:PEGB3, pass, PUGB6
			10'd122 : rdata = 48'b110001110000011000000000000000000000000000001110;
			// PEs: 32 -> 33
			// srcs: (128, 95)(2091) 0 --> (2091) 0:NI0, pass, PENB
			10'd123 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 24 -> 32
			// srcs: (129, 96)(2094) 4 --> (2094) 4:PUNB, pass, NI0
			10'd124 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 24 -> 33
			// srcs: (130, 97)(2095) 0 --> (2095) 0:PUNB, pass, PENB
			10'd125 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 36 -> 16
			// srcs: (131, 159)(1732) 0 --> (1732) 0:PEGB4, pass, PUGB2
			10'd126 : rdata = 48'b110001110000100000000000000000000000000000001010;
			// PEs: 38 -> 40
			// srcs: (132, 161)(1738) 0 --> (1738) 0:PEGB6, pass, PUNB
			10'd127 : rdata = 48'b110001110000110000000000000000000000001000000000;
			// PEs: 39 -> 8
			// srcs: (133, 162)(1741) 0 --> (1741) 0:PENB, pass, PUGB1
			10'd128 : rdata = 48'b110001101111111000000000000000000000000000001001;
			// PEs: 39 -> 48
			// srcs: (134, 167)(2544) -3 --> (2544) -3:PENB, pass, PUGB6
			10'd129 : rdata = 48'b110001101111111000000000000000000000000000001110;
			// PEs: 33 -> 0
			// srcs: (135, 179)(1903) 3 --> (1903) 3:PEGB1, pass, PUGB0
			10'd130 : rdata = 48'b110001110000001000000000000000000000000000001000;
			// PEs: 32 -> 33
			// srcs: (136, 98)(2094) 4 --> (2094) 4:NI0, pass, PENB
			10'd131 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 24 -> 32
			// srcs: (137, 106)(2168) 0 --> (2168) 0:PUNB, pass, NI0
			10'd132 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 24 -> 33
			// srcs: (138, 107)(2169) -2 --> (2169) -2:PUNB, pass, PENB
			10'd133 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 33 -> 8
			// srcs: (142, 168)(2592) 5 --> (2592) 5:PEGB1, pass, PUGB1
			10'd134 : rdata = 48'b110001110000001000000000000000000000000000001001;
			// PEs: 34 -> 24
			// srcs: (143, 172)(2624) 10 --> (2624) 10:PEGB2, pass, PUGB3
			10'd135 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 32 -> 33
			// srcs: (144, 108)(2168) 0 --> (2168) 0:NI0, pass, PENB
			10'd136 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 24 -> 32
			// srcs: (145, 109)(2171) 4 --> (2171) 4:PUNB, pass, NI0
			10'd137 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 24 -> 33
			// srcs: (146, 110)(2172) 0 --> (2172) 0:PUNB, pass, PENB
			10'd138 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 36 -> 40
			// srcs: (147, 182)(1912) 3 --> (1912) 3:PEGB4, pass, PUNB
			10'd139 : rdata = 48'b110001110000100000000000000000000000001000000000;
			// PEs: 37 -> 48
			// srcs: (148, 183)(1915) 0 --> (1915) 0:PEGB5, pass, PUGB6
			10'd140 : rdata = 48'b110001110000101000000000000000000000000000001110;
			// PEs: 39 -> 0
			// srcs: (149, 229)(3119) -4 --> (3119) -4:PENB, pass, PUGB0
			10'd141 : rdata = 48'b110001101111111000000000000000000000000000001000;
			// PEs: 32 -> 33
			// srcs: (152, 111)(2171) 4 --> (2171) 4:NI0, pass, PENB
			10'd142 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 24 -> 32
			// srcs: (153, 112)(2174) 3 --> (2174) 3:PUNB, pass, NI0
			10'd143 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 24 -> 33
			// srcs: (154, 113)(2175) 6 --> (2175) 6:PUNB, pass, PENB
			10'd144 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 35 -> 8
			// srcs: (155, 173)(2626) 0 --> (2626) 0:PEGB3, pass, PUGB1
			10'd145 : rdata = 48'b110001110000011000000000000000000000000000001001;
			// PEs: 33 -> 40
			// srcs: (156, 186)(2705) -4 --> (2705) -4:PEGB1, pass, PUNB
			10'd146 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 37 -> 24
			// srcs: (157, 219)(2283) -6 --> (2283) -6:PEGB5, pass, PUGB3
			10'd147 : rdata = 48'b110001110000101000000000000000000000000000001011;
			// PEs: 33 -> 56
			// srcs: (159, 209)(2951) 4 --> (2951) 4:PEGB1, pass, PUGB7
			10'd148 : rdata = 48'b110001110000001000000000000000000000000000001111;
			// PEs: 32 -> 33
			// srcs: (160, 114)(2174) 3 --> (2174) 3:NI0, pass, PENB
			10'd149 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 34 -> 8
			// srcs: (163, 180)(1906) 6 --> (1906) 6:PEGB2, pass, PUGB1
			10'd150 : rdata = 48'b110001110000010000000000000000000000000000001001;
			// PEs: 33 -> 40
			// srcs: (164, 187)(2709) -1 --> (2709) -1:PEGB1, pass, PUNB
			10'd151 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 34 -> 24
			// srcs: (165, 230)(3123) 7 --> (3123) 7:PEGB2, pass, PUGB3
			10'd152 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 36 -> 56
			// srcs: (168, 218)(2280) 0 --> (2280) 0:PEGB4, pass, PUGB7
			10'd153 : rdata = 48'b110001110000100000000000000000000000000000001111;
			// PEs: 33 -> 40
			// srcs: (172, 188)(2711) -4 --> (2711) -4:PEGB1, pass, PUNB
			10'd154 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 39 -> 56
			// srcs: (173, 221)(2289) 0 --> (2289) 0:PENB, pass, PUGB7
			10'd155 : rdata = 48'b110001101111111000000000000000000000000000001111;
			// PEs: 33 -> 40
			// srcs: (180, 192)(2788) -3 --> (2788) -3:PEGB1, pass, PUNB
			10'd156 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 33 -> 40
			// srcs: (188, 193)(2790) -10 --> (2790) -10:PEGB1, pass, PUNB
			10'd157 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 24 -> 32
			// srcs: (214, 125)(1769) -2 --> (1769) -2:PUNB, pass, NI0
			10'd158 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 24 -> 35
			// srcs: (230, 126)(1770) 0 --> (1770) 0:PUNB, pass, PEGB3
			10'd159 : rdata = 48'b110001101111111100000000000000000000000010110000;
			// PEs: 32 -> 35
			// srcs: (239, 127)(1769) -2 --> (1769) -2:NI0, pass, PEGB3
			10'd160 : rdata = 48'b110001010000000000000000000000000000000010110000;
			// PEs: 24 -> 32
			// srcs: (246, 128)(1771) 1 --> (1771) 1:PUNB, pass, NI0
			10'd161 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 24 -> 36
			// srcs: (261, 129)(1772) 0 --> (1772) 0:PUNB, pass, PEGB4
			10'd162 : rdata = 48'b110001101111111100000000000000000000000011000000;
			// PEs: 32 -> 36
			// srcs: (270, 130)(1771) 1 --> (1771) 1:NI0, pass, PEGB4
			10'd163 : rdata = 48'b110001010000000000000000000000000000000011000000;
			// PEs: 24 -> 32
			// srcs: (274, 131)(2014) 0 --> (2014) 0:PUNB, pass, NI0
			10'd164 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 36 -> 48
			// srcs: (283, 248)(2554) -1 --> (2554) -1:PEGB4, pass, PUGB6
			10'd165 : rdata = 48'b110001110000100000000000000000000000000000001110;
			// PEs: 24 -> 33
			// srcs: (288, 132)(2015) 4 --> (2015) 4:PUNB, pass, PENB
			10'd166 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 32 -> 33
			// srcs: (294, 133)(2014) 0 --> (2014) 0:NI0, pass, PENB
			10'd167 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 0 -> 32
			// srcs: (295, 136)(2369) -1 --> (2369) -1:PUGB0, pass, NI0
			10'd168 : rdata = 48'b110001110000000100000000000100000000000000000000;
			// PEs: 48 -> 33
			// srcs: (296, 137)(1588) 2 --> (1588) 2:PUGB6, pass, PENB
			10'd169 : rdata = 48'b110001110000110100000000000000000000000100000000;
			// PEs: 33 -> 40
			// srcs: (301, 194)(2796) 4 --> (2796) 4:PEGB1, pass, PUNB
			10'd170 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 32 -> 33
			// srcs: (302, 138)(2369) -1 --> (2369) -1:NI0, pass, PENB
			10'd171 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 8 -> 32
			// srcs: (303, 139)(2388) -2 --> (2388) -2:PUGB1, pass, NI0
			10'd172 : rdata = 48'b110001110000001100000000000100000000000000000000;
			// PEs: 56 -> 33
			// srcs: (304, 140)(1609) 6 --> (1609) 6:PUGB7, pass, PENB
			10'd173 : rdata = 48'b110001110000111100000000000000000000000100000000;
			// PEs: 33 -> 0
			// srcs: (309, 234)(2370) 1 --> (2370) 1:PEGB1, pass, PUGB0
			10'd174 : rdata = 48'b110001110000001000000000000000000000000000001000;
			// PEs: 32 -> 33
			// srcs: (310, 141)(2388) -2 --> (2388) -2:NI0, pass, PENB
			10'd175 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 24 -> 32
			// srcs: (311, 142)(2419) 3 --> (2419) 3:PUNB, pass, NI0
			10'd176 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 0 -> 33
			// srcs: (312, 143)(1640) -1 --> (1640) -1:PUGB0, pass, PENB
			10'd177 : rdata = 48'b110001110000000100000000000000000000000100000000;
			// PEs: 37 -> 40
			// srcs: (313, 199)(2099) 0 --> (2099) 0:PEGB5, pass, PUNB
			10'd178 : rdata = 48'b110001110000101000000000000000000000001000000000;
			// PEs: 38 -> 40
			// srcs: (314, 200)(2102) 0 --> (2102) 0:PEGB6, pass, PUNB
			10'd179 : rdata = 48'b110001110000110000000000000000000000001000000000;
			// PEs: 32 -> 33
			// srcs: (318, 144)(2419) 3 --> (2419) 3:NI0, pass, PENB
			10'd180 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 56 -> 32
			// srcs: (319, 146)(2460) -5 --> (2460) -5:PUGB7, pass, NI0
			10'd181 : rdata = 48'b110001110000111100000000000100000000000000000000;
			// PEs: 16 -> 33
			// srcs: (320, 147)(1680) 3 --> (1680) 3:PUGB2, pass, PENB
			10'd182 : rdata = 48'b110001110000010100000000000000000000000100000000;
			// PEs: 39 -> 40
			// srcs: (321, 201)(2105) -1 --> (2105) -1:PENB, pass, PUNB
			10'd183 : rdata = 48'b110001101111111000000000000000000000001000000000;
			// PEs: 32 -> 33
			// srcs: (326, 148)(2460) -5 --> (2460) -5:NI0, pass, PENB
			10'd184 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 40 -> 32
			// srcs: (327, 153)(2478) 4 --> (2478) 4:PUGB5, pass, NI0
			10'd185 : rdata = 48'b110001110000101100000000000100000000000000000000;
			// PEs: 24 -> 33
			// srcs: (328, 154)(1698) -4 --> (1698) -4:PUNB, pass, PENB
			10'd186 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 33 -> 40
			// srcs: (329, 208)(2949) -2 --> (2949) -2:PEGB1, pass, PUNB
			10'd187 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 33 -> 56
			// srcs: (333, 240)(2461) -2 --> (2461) -2:PEGB1, pass, PUGB7
			10'd188 : rdata = 48'b110001110000001000000000000000000000000000001111;
			// PEs: 32 -> 33
			// srcs: (334, 155)(2478) 4 --> (2478) 4:NI0, pass, PENB
			10'd189 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 8 -> 33
			// srcs: (335, 160)(2514) 3 --> (2514) 3:PUGB1, pass, PENB
			10'd190 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 16 -> 32
			// srcs: (336, 163)(2528) -1 --> (2528) -1:PUGB2, pass, NI0
			10'd191 : rdata = 48'b110001110000010100000000000100000000000000000000;
			// PEs: 40 -> 33
			// srcs: (337, 164)(1750) 0 --> (1750) 0:PUGB5, pass, PENB
			10'd192 : rdata = 48'b110001110000101100000000000000000000000100000000;
			// PEs: 33 -> 40
			// srcs: (338, 215)(2271) 4 --> (2271) 4:PEGB1, pass, PUNB
			10'd193 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 32 -> 33
			// srcs: (343, 165)(2528) -1 --> (2528) -1:NI0, pass, PENB
			10'd194 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 48 -> 33
			// srcs: (344, 166)(1765) 0 --> (1765) 0:PUGB6, pass, PENB
			10'd195 : rdata = 48'b110001110000110100000000000000000000000100000000;
			// PEs: 16 -> 32
			// srcs: (345, 169)(2608) 0 --> (2608) 0:PUGB2, pass, NI0
			10'd196 : rdata = 48'b110001110000010100000000000100000000000000000000;
			// PEs: 0 -> 33
			// srcs: (346, 170)(1830) 0 --> (1830) 0:PUGB0, pass, PENB
			10'd197 : rdata = 48'b110001110000000100000000000000000000000100000000;
			// PEs: 34 -> 40
			// srcs: (347, 216)(2274) 4 --> (2274) 4:PEGB2, pass, PUNB
			10'd198 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 32 -> 33
			// srcs: (352, 171)(2608) 0 --> (2608) 0:NI0, pass, PENB
			10'd199 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 8 -> 33
			// srcs: (353, 175)(1854) 0 --> (1854) 0:PUGB1, pass, PENB
			10'd200 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 56 -> 32
			// srcs: (354, 176)(2661) 0 --> (2661) 0:PUGB7, pass, NI0
			10'd201 : rdata = 48'b110001110000111100000000000100000000000000000000;
			// PEs: 24 -> 33
			// srcs: (355, 177)(1882) 0 --> (1882) 0:PUNB, pass, PENB
			10'd202 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 35 -> 40
			// srcs: (356, 217)(2277) 0 --> (2277) 0:PEGB3, pass, PUNB
			10'd203 : rdata = 48'b110001110000011000000000000000000000001000000000;
			// PEs: 38 -> 40
			// srcs: (357, 228)(3117) -1 --> (3117) -1:PEGB6, pass, PUNB
			10'd204 : rdata = 48'b110001110000110000000000000000000000001000000000;
			// PEs: 33 -> 40
			// srcs: (358, 241)(2479) 0 --> (2479) 0:PEGB1, pass, PUNB
			10'd205 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 33 -> 40
			// srcs: (359, 245)(2515) 1 --> (2515) 1:PEGB1, pass, PUNB
			10'd206 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 33 -> 40
			// srcs: (360, 247)(2543) 0 --> (2543) 0:PEGB1, pass, PUNB
			10'd207 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 32 -> 33
			// srcs: (361, 178)(2661) 0 --> (2661) 0:NI0, pass, PENB
			10'd208 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 16 -> 33
			// srcs: (362, 181)(2686) -3 --> (2686) -3:PUGB2, pass, PENB
			10'd209 : rdata = 48'b110001110000010100000000000000000000000100000000;
			// PEs: 24 -> 33
			// srcs: (363, 184)(2700) 0 --> (2700) 0:PUNB, pass, PENB
			10'd210 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 24 -> 38
			// srcs: (364, 185)(2703) -8 --> (2703) -8:PUNB, pass, PEGB6
			10'd211 : rdata = 48'b110001101111111100000000000000000000000011100000;
			// PEs: 16 -> 32
			// srcs: (365, 189)(2774) 0 --> (2774) 0:PUGB2, pass, NI0
			10'd212 : rdata = 48'b110001110000010100000000000100000000000000000000;
			// PEs: 0 -> 33
			// srcs: (366, 190)(1995) 4 --> (1995) 4:PUGB0, pass, PENB
			10'd213 : rdata = 48'b110001110000000100000000000000000000000100000000;
			// PEs: 33 -> 8
			// srcs: (367, 250)(2632) 0 --> (2632) 0:PEGB1, pass, PUGB1
			10'd214 : rdata = 48'b110001110000001000000000000000000000000000001001;
			// PEs: 33 -> 24
			// srcs: (368, 254)(2662) 0 --> (2662) 0:PEGB1, pass, PUGB3
			10'd215 : rdata = 48'b110001110000001000000000000000000000000000001011;
			// PEs: 33 -> 0
			// srcs: (369, 255)(2687) -7 --> (2687) -7:PEGB1, pass, PUGB0
			10'd216 : rdata = 48'b110001110000001000000000000000000000000000001000;
			// PEs: 32 -> 33
			// srcs: (376, 191)(2774) 0 --> (2774) 0:NI0, pass, PENB
			10'd217 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 48 -> 32
			// srcs: (377, 195)(2813) 10 --> (2813) 10:PUGB6, pass, NI0
			10'd218 : rdata = 48'b110001110000110100000000000100000000000000000000;
			// PEs: 8 -> 33
			// srcs: (378, 196)(2035) -1 --> (2035) -1:PUGB1, pass, PENB
			10'd219 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 38 -> 40
			// srcs: (379, 257)(2704) -6 --> (2704) -6:PEGB6, pass, PUNB
			10'd220 : rdata = 48'b110001110000110000000000000000000000001000000000;
			// PEs: 32 -> 33
			// srcs: (384, 197)(2813) 10 --> (2813) 10:NI0, pass, PENB
			10'd221 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 24 -> 33
			// srcs: (385, 198)(2864) 3 --> (2864) 3:PUNB, pass, PENB
			10'd222 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 8 -> 32
			// srcs: (386, 202)(2922) 0 --> (2922) 0:PUGB1, pass, NI0
			10'd223 : rdata = 48'b110001110000001100000000000100000000000000000000;
			// PEs: 48 -> 33
			// srcs: (387, 203)(2145) 1 --> (2145) 1:PUGB6, pass, PENB
			10'd224 : rdata = 48'b110001110000110100000000000000000000000100000000;
			// PEs: 37 -> 40
			// srcs: (388, 264)(2875) 8 --> (2875) 8:PEGB5, pass, PUNB
			10'd225 : rdata = 48'b110001110000101000000000000000000000001000000000;
			// PEs: 33 -> 48
			// srcs: (391, 259)(2814) 9 --> (2814) 9:PEGB1, pass, PUGB6
			10'd226 : rdata = 48'b110001110000001000000000000000000000000000001110;
			// PEs: 32 -> 33
			// srcs: (393, 204)(2922) 0 --> (2922) 0:NI0, pass, PENB
			10'd227 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 24 -> 32
			// srcs: (394, 205)(2946) 0 --> (2946) 0:PUNB, pass, NI0
			10'd228 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 56 -> 33
			// srcs: (395, 206)(2167) -1 --> (2167) -1:PUGB7, pass, PENB
			10'd229 : rdata = 48'b110001110000111100000000000000000000000100000000;
			// PEs: 32 -> 33
			// srcs: (401, 207)(2946) 0 --> (2946) 0:NI0, pass, PENB
			10'd230 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 56 -> 33
			// srcs: (402, 210)(2176) 2 --> (2176) 2:PUGB7, pass, PENB
			10'd231 : rdata = 48'b110001110000111100000000000000000000000100000000;
			// PEs: 40 -> 32
			// srcs: (403, 211)(2960) 2 --> (2960) 2:PUGB5, pass, NI0
			10'd232 : rdata = 48'b110001110000101100000000000100000000000000000000;
			// PEs: 0 -> 33
			// srcs: (404, 212)(2182) -3 --> (2182) -3:PUGB0, pass, PENB
			10'd233 : rdata = 48'b110001110000000100000000000000000000000100000000;
			// PEs: 33 -> 8
			// srcs: (409, 267)(2956) 11 --> (2956) 11:PEGB1, pass, PUGB1
			10'd234 : rdata = 48'b110001110000001000000000000000000000000000001001;
			// PEs: 32 -> 33
			// srcs: (410, 213)(2960) 2 --> (2960) 2:NI0, pass, PENB
			10'd235 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 24 -> 33
			// srcs: (411, 214)(2265) 2 --> (2265) 2:PUNB, pass, PENB
			10'd236 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 48 -> 33
			// srcs: (412, 220)(3064) -2 --> (3064) -2:PUGB6, pass, PENB
			10'd237 : rdata = 48'b110001110000110100000000000000000000000100000000;
			// PEs: 56 -> 32
			// srcs: (413, 222)(3075) 4 --> (3075) 4:PUGB7, pass, NI0
			10'd238 : rdata = 48'b110001110000111100000000000100000000000000000000;
			// PEs: 40 -> 33
			// srcs: (414, 223)(2298) 0 --> (2298) 0:PUGB5, pass, PENB
			10'd239 : rdata = 48'b110001110000101100000000000000000000000100000000;
			// PEs: 33 -> 24
			// srcs: (417, 268)(2961) -1 --> (2961) -1:PEGB1, pass, PUGB3
			10'd240 : rdata = 48'b110001110000001000000000000000000000000000001011;
			// PEs: 32 -> 33
			// srcs: (425, 224)(3075) 4 --> (3075) 4:NI0, pass, PENB
			10'd241 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 16 -> 32
			// srcs: (426, 225)(3100) 2 --> (3100) 2:PUGB2, pass, NI0
			10'd242 : rdata = 48'b110001110000010100000000000100000000000000000000;
			// PEs: 48 -> 33
			// srcs: (427, 226)(2323) 2 --> (2323) 2:PUGB6, pass, PENB
			10'd243 : rdata = 48'b110001110000110100000000000000000000000100000000;
			// PEs: 33 -> 0
			// srcs: (428, 272)(3065) -3 --> (3065) -3:PEGB1, pass, PUGB0
			10'd244 : rdata = 48'b110001110000001000000000000000000000000000001000;
			// PEs: 33 -> 24
			// srcs: (432, 276)(3076) 4 --> (3076) 4:PEGB1, pass, PUGB3
			10'd245 : rdata = 48'b110001110000001000000000000000000000000000001011;
			// PEs: 32 -> 33
			// srcs: (433, 227)(3100) 2 --> (3100) 2:NI0, pass, PENB
			10'd246 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 40 -> 32
			// srcs: (434, 231)(3125) -2 --> (3125) -2:PUGB5, pass, NI0
			10'd247 : rdata = 48'b110001110000101100000000000100000000000000000000;
			// PEs: 33 -> 56
			// srcs: (440, 277)(3101) 4 --> (3101) 4:PEGB1, pass, PUGB7
			10'd248 : rdata = 48'b110001110000001000000000000000000000000000001111;
			// PEs: 56 -> 33
			// srcs: (562, 232)(2350) -3 --> (2350) -3:PUGB7, pass, PENB
			10'd249 : rdata = 48'b110001110000111100000000000000000000000100000000;
			// PEs: 32 -> 33
			// srcs: (568, 233)(3125) -2 --> (3125) -2:NI0, pass, PENB
			10'd250 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 24 -> 33
			// srcs: (569, 235)(2387) 3 --> (2387) 3:PUNB, pass, PENB
			10'd251 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 24 -> 33
			// srcs: (570, 236)(2418) -1 --> (2418) -1:PUNB, pass, PENB
			10'd252 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 16 -> 32
			// srcs: (571, 237)(2435) 2 --> (2435) 2:PUGB2, pass, NI0
			10'd253 : rdata = 48'b110001110000010100000000000100000000000000000000;
			// PEs: 40 -> 33
			// srcs: (572, 238)(2437) 5 --> (2437) 5:PUGB5, pass, PENB
			10'd254 : rdata = 48'b110001110000101100000000000000000000000100000000;
			// PEs: 33 -> 48
			// srcs: (576, 279)(2390) 7 --> (2390) 7:PEGB1, pass, PUGB6
			10'd255 : rdata = 48'b110001110000001000000000000000000000000000001110;
			// PEs: 33 -> 56
			// srcs: (577, 283)(2421) 1 --> (2421) 1:PEGB1, pass, PUGB7
			10'd256 : rdata = 48'b110001110000001000000000000000000000000000001111;
			// PEs: 32 -> 33
			// srcs: (578, 239)(2435) 2 --> (2435) 2:NI0, pass, PENB
			10'd257 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 0 -> 32
			// srcs: (579, 242)(2504) 1 --> (2504) 1:PUGB0, pass, NI0
			10'd258 : rdata = 48'b110001110000000100000000000100000000000000000000;
			// PEs: 24 -> 33
			// srcs: (580, 243)(2506) 14 --> (2506) 14:PUNB, pass, PENB
			10'd259 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 39 -> 48
			// srcs: (581, 300)(3045) -9 --> (3045) -9:PENB, pass, PUGB6
			10'd260 : rdata = 48'b110001101111111000000000000000000000000000001110;
			// PEs: 32 -> 33
			// srcs: (586, 244)(2504) 1 --> (2504) 1:NI0, pass, PENB
			10'd261 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 24 -> 33
			// srcs: (587, 246)(2527) 0 --> (2527) 0:PUNB, pass, PENB
			10'd262 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 16 -> 33
			// srcs: (588, 249)(2607) 2 --> (2607) 2:PUGB2, pass, PENB
			10'd263 : rdata = 48'b110001110000010100000000000000000000000100000000;
			// PEs: 16 -> 32
			// srcs: (589, 251)(2656) -4 --> (2656) -4:PUGB2, pass, NI0
			10'd264 : rdata = 48'b110001110000010100000000000100000000000000000000;
			// PEs: 48 -> 33
			// srcs: (590, 252)(2658) 2 --> (2658) 2:PUGB6, pass, PENB
			10'd265 : rdata = 48'b110001110000110100000000000000000000000100000000;
			// PEs: 33 -> 16
			// srcs: (593, 285)(2507) 15 --> (2507) 15:PEGB1, pass, PUGB2
			10'd266 : rdata = 48'b110001110000001000000000000000000000000000001010;
			// PEs: 33 -> 24
			// srcs: (594, 286)(2530) -1 --> (2530) -1:PEGB1, pass, PUGB3
			10'd267 : rdata = 48'b110001110000001000000000000000000000000000001011;
			// PEs: 32 -> 33
			// srcs: (596, 253)(2656) -4 --> (2656) -4:NI0, pass, PENB
			10'd268 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 24 -> 33
			// srcs: (597, 256)(2699) 7 --> (2699) 7:PUNB, pass, PENB
			10'd269 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 24 -> 33
			// srcs: (599, 258)(2773) 3 --> (2773) 3:PUNB, pass, PENB
			10'd270 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 33 -> 40
			// srcs: (603, 288)(2659) -2 --> (2659) -2:PEGB1, pass, PUNB
			10'd271 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 33 -> 40
			// srcs: (604, 289)(2702) 13 --> (2702) 13:PEGB1, pass, PUNB
			10'd272 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 24 -> 32
			// srcs: (607, 260)(2821) 5 --> (2821) 5:PUNB, pass, NI0
			10'd273 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 56 -> 33
			// srcs: (608, 261)(2823) 5 --> (2823) 5:PUGB7, pass, PENB
			10'd274 : rdata = 48'b110001110000111100000000000000000000000100000000;
			// PEs: 32 -> 33
			// srcs: (617, 262)(2821) 5 --> (2821) 5:NI0, pass, PENB
			10'd275 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 48 -> 33
			// srcs: (618, 265)(2925) -3 --> (2925) -3:PUGB6, pass, PENB
			10'd276 : rdata = 48'b110001110000110100000000000000000000000100000000;
			// PEs: 16 -> 32
			// srcs: (619, 269)(2973) -10 --> (2973) -10:PUGB2, pass, NI0
			10'd277 : rdata = 48'b110001110000010100000000000100000000000000000000;
			// PEs: 48 -> 33
			// srcs: (620, 270)(2975) 0 --> (2975) 0:PUGB6, pass, PENB
			10'd278 : rdata = 48'b110001110000110100000000000000000000000100000000;
			// PEs: 33 -> 40
			// srcs: (624, 294)(2824) 10 --> (2824) 10:PEGB1, pass, PUNB
			10'd279 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 33 -> 24
			// srcs: (625, 297)(2926) -2 --> (2926) -2:PEGB1, pass, PUGB3
			10'd280 : rdata = 48'b110001110000001000000000000000000000000000001011;
			// PEs: 32 -> 33
			// srcs: (626, 271)(2973) -10 --> (2973) -10:NI0, pass, PENB
			10'd281 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 48 -> 32
			// srcs: (627, 273)(3070) 4 --> (3070) 4:PUGB6, pass, NI0
			10'd282 : rdata = 48'b110001110000110100000000000100000000000000000000;
			// PEs: 8 -> 33
			// srcs: (628, 274)(3072) 0 --> (3072) 0:PUGB1, pass, PENB
			10'd283 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 35 -> 40
			// srcs: (632, 296)(2873) -2 --> (2873) -2:PEGB3, pass, PUNB
			10'd284 : rdata = 48'b110001110000011000000000000000000000001000000000;
			// PEs: 32 -> 33
			// srcs: (634, 275)(3070) 4 --> (3070) 4:NI0, pass, PENB
			10'd285 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 24 -> 38
			// srcs: (1096, 263)(2863) 0 --> (2863) 0:PUNB, pass, PEGB6
			10'd286 : rdata = 48'b110001101111111100000000000000000000000011100000;
			// PEs: 24 -> 36
			// srcs: (1097, 266)(2945) 11 --> (2945) 11:PUNB, pass, PEGB4
			10'd287 : rdata = 48'b110001101111111100000000000000000000000011000000;
			// PEs: 24 -> 33
			// srcs: (1098, 278)(3124) 9 --> (3124) 9:PUNB, pass, PENB
			10'd288 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 24 -> 32
			// srcs: (1099, 280)(2410) 6 --> (2410) 6:PUNB, pass, NI0
			10'd289 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 48 -> 33
			// srcs: (1100, 281)(2415) -3 --> (2415) -3:PUGB6, pass, PENB
			10'd290 : rdata = 48'b110001110000110100000000000000000000000100000000;
			// PEs: 32 -> 33
			// srcs: (1106, 282)(2410) 6 --> (2410) 6:NI0, pass, PENB
			10'd291 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 24 -> 33
			// srcs: (1107, 284)(2433) 3 --> (2433) 3:PUNB, pass, PENB
			10'd292 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 24 -> 33
			// srcs: (1108, 287)(2605) 16 --> (2605) 16:PUNB, pass, PENB
			10'd293 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 24 -> 33
			// srcs: (1109, 290)(2781) 5 --> (2781) 5:PUNB, pass, PENB
			10'd294 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 56 -> 32
			// srcs: (1110, 291)(2787) 0 --> (2787) 0:PUGB7, pass, NI0
			10'd295 : rdata = 48'b110001110000111100000000000100000000000000000000;
			// PEs: 40 -> 33
			// srcs: (1111, 292)(2792) -13 --> (2792) -13:PUGB5, pass, PENB
			10'd296 : rdata = 48'b110001110000101100000000000000000000000100000000;
			// PEs: 24 -> 35
			// srcs: (1112, 295)(2861) 3 --> (2861) 3:PUNB, pass, PEGB3
			10'd297 : rdata = 48'b110001101111111100000000000000000000000010110000;
			// PEs: 36 -> 8
			// srcs: (1113, 298)(2948) 10 --> (2948) 10:PEGB4, pass, PUGB1
			10'd298 : rdata = 48'b110001110000100000000000000000000000000000001001;
			// PEs: 24 -> 37
			// srcs: (1114, 302)(3132) 7 --> (3132) 7:PUNB, pass, PEGB5
			10'd299 : rdata = 48'b110001101111111100000000000000000000000011010000;
			// PEs: 33 -> 40
			// srcs: (1115, 306)(2416) 3 --> (2416) 3:PEGB1, pass, PUNB
			10'd300 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 33 -> 48
			// srcs: (1116, 307)(2439) 10 --> (2439) 10:PEGB1, pass, PUGB6
			10'd301 : rdata = 48'b110001110000001000000000000000000000000000001110;
			// PEs: 32 -> 33
			// srcs: (1117, 293)(2787) 0 --> (2787) 0:NI0, pass, PENB
			10'd302 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 56 -> 33
			// srcs: (1118, 299)(2971) 7 --> (2971) 7:PUGB7, pass, PENB
			10'd303 : rdata = 48'b110001110000111100000000000000000000000100000000;
			// PEs: 0 -> 33
			// srcs: (1119, 301)(3068) -5 --> (3068) -5:PUGB0, pass, PENB
			10'd304 : rdata = 48'b110001110000000100000000000000000000000100000000;
			// PEs: 48 -> 32
			// srcs: (1120, 303)(2391) 4 --> (2391) 4:PUGB6, pass, NI0
			10'd305 : rdata = 48'b110001110000110100000000000100000000000000000000;
			// PEs: 16 -> 33
			// srcs: (1121, 304)(2402) -10 --> (2402) -10:PUGB2, pass, PENB
			10'd306 : rdata = 48'b110001110000010100000000000000000000000100000000;
			// PEs: 33 -> 16
			// srcs: (1122, 308)(2611) 18 --> (2611) 18:PEGB1, pass, PUGB2
			10'd307 : rdata = 48'b110001110000001000000000000000000000000000001010;
			// PEs: 35 -> 40
			// srcs: (1124, 312)(2867) 2 --> (2867) 2:PEGB3, pass, PUNB
			10'd308 : rdata = 48'b110001110000011000000000000000000000001000000000;
			// PEs: 33 -> 0
			// srcs: (1125, 313)(2977) -3 --> (2977) -3:PEGB1, pass, PUGB0
			10'd309 : rdata = 48'b110001110000001000000000000000000000000000001000;
			// PEs: 33 -> 40
			// srcs: (1126, 314)(3074) -1 --> (3074) -1:PEGB1, pass, PUNB
			10'd310 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 32 -> 33
			// srcs: (1127, 305)(2391) 4 --> (2391) 4:NI0, pass, PENB
			10'd311 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 8 -> 32
			// srcs: (1128, 309)(2634) 19 --> (2634) 19:PUGB1, pass, NI0
			10'd312 : rdata = 48'b110001110000001100000000000100000000000000000000;
			// PEs: 48 -> 33
			// srcs: (1129, 310)(2645) 2 --> (2645) 2:PUGB6, pass, PENB
			10'd313 : rdata = 48'b110001110000110100000000000000000000000100000000;
			// PEs: 37 -> 8
			// srcs: (1130, 315)(3133) 11 --> (3133) 11:PEGB5, pass, PUGB1
			10'd314 : rdata = 48'b110001110000101000000000000000000000000000001001;
			// PEs: 34 -> 8
			// srcs: (1133, 321)(2794) -1 --> (2794) -1:PEGB2, pass, PUGB1
			10'd315 : rdata = 48'b110001110000010000000000000000000000000000001001;
			// PEs: 33 -> 24
			// srcs: (1134, 316)(2403) -6 --> (2403) -6:PEGB1, pass, PUGB3
			10'd316 : rdata = 48'b110001110000001000000000000000000000000000001011;
			// PEs: 32 -> 33
			// srcs: (1135, 311)(2634) 19 --> (2634) 19:NI0, pass, PENB
			10'd317 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 24 -> 32
			// srcs: (1136, 317)(2525) 19 --> (2525) 19:PUNB, pass, NI0
			10'd318 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 0 -> 33
			// srcs: (1137, 318)(2548) -21 --> (2548) -21:PUGB0, pass, PENB
			10'd319 : rdata = 48'b110001110000000100000000000000000000000100000000;
			// PEs: 33 -> 40
			// srcs: (1142, 320)(2646) 21 --> (2646) 21:PEGB1, pass, PUNB
			10'd320 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 32 -> 33
			// srcs: (1143, 319)(2525) 19 --> (2525) 19:NI0, pass, PENB
			10'd321 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 33 -> 40
			// srcs: (1150, 325)(2549) -2 --> (2549) -2:PEGB1, pass, PUNB
			10'd322 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 16 -> 32
			// srcs: (1179, 322)(2916) 16 --> (2916) 16:PUGB2, pass, NI0
			10'd323 : rdata = 48'b110001110000010100000000000100000000000000000000;
			// PEs: 56 -> 33
			// srcs: (1407, 323)(2939) 11 --> (2939) 11:PUGB7, pass, PENB
			10'd324 : rdata = 48'b110001110000111100000000000000000000000100000000;
			// PEs: 32 -> 33
			// srcs: (1414, 324)(2916) 16 --> (2916) 16:NI0, pass, PENB
			10'd325 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 33 -> 24
			// srcs: (1421, 326)(2940) 27 --> (2940) 27:PEGB1, pass, PUGB3
			10'd326 : rdata = 48'b110001110000001000000000000000000000000000001011;
			// PEs: 56 -> 32
			// srcs: (1428, 327)(2990) -1 --> (2990) -1:PUGB7, pass, NI0
			10'd327 : rdata = 48'b110001110000111100000000000100000000000000000000;
			// PEs: 16 -> 33
			// srcs: (1429, 328)(3038) -37 --> (3038) -37:PUGB2, pass, PENB
			10'd328 : rdata = 48'b110001110000010100000000000000000000000100000000;
			// PEs: 32 -> 33
			// srcs: (1435, 329)(2990) -1 --> (2990) -1:NI0, pass, PENB
			10'd329 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 33 -> 40
			// srcs: (1442, 330)(3039) -38 --> (3039) -38:PEGB1, pass, PUNB
			10'd330 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 8 -> 33
			// srcs: (1549, 331)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd331 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 34
			// srcs: (1550, 332)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd332 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 35
			// srcs: (1552, 333)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd333 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 36
			// srcs: (1553, 334)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd334 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 37
			// srcs: (1555, 335)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd335 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 38
			// srcs: (1556, 336)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd336 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 39
			// srcs: (1558, 337)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd337 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 33
			// srcs: (1629, 338)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd338 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 34
			// srcs: (1630, 339)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd339 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 35
			// srcs: (1632, 340)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd340 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 36
			// srcs: (1633, 341)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd341 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 37
			// srcs: (1635, 342)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd342 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 38
			// srcs: (1636, 343)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd343 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 39
			// srcs: (1638, 344)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd344 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 33
			// srcs: (1655, 345)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd345 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 34
			// srcs: (1662, 346)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd346 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 35
			// srcs: (1665, 347)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd347 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 36
			// srcs: (1668, 348)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd348 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 37
			// srcs: (1671, 349)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd349 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 38
			// srcs: (1674, 350)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd350 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 39
			// srcs: (1677, 351)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd351 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 33
			// srcs: (1709, 352)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd352 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 34
			// srcs: (1710, 353)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd353 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 35
			// srcs: (1712, 354)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd354 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 36
			// srcs: (1713, 355)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd355 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 37
			// srcs: (1715, 356)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd356 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 38
			// srcs: (1716, 357)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd357 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 39
			// srcs: (1718, 358)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd358 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 33
			// srcs: (1791, 359)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd359 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 34
			// srcs: (1792, 360)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd360 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 35
			// srcs: (1794, 361)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd361 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 36
			// srcs: (1795, 362)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd362 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 37
			// srcs: (1797, 363)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd363 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 38
			// srcs: (1798, 364)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd364 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 39
			// srcs: (1800, 365)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd365 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 33
			// srcs: (1839, 366)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd366 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 34
			// srcs: (1842, 367)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd367 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 35
			// srcs: (1845, 368)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd368 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 36
			// srcs: (1848, 369)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd369 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 37
			// srcs: (1851, 370)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd370 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 38
			// srcs: (1858, 371)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd371 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 39
			// srcs: (1861, 372)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd372 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 33
			// srcs: (1871, 373)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd373 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 34
			// srcs: (1872, 374)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd374 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 35
			// srcs: (1874, 375)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd375 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 36
			// srcs: (1875, 376)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd376 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 37
			// srcs: (1877, 377)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd377 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 38
			// srcs: (1878, 378)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd378 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 39
			// srcs: (1880, 379)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd379 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 33
			// srcs: (1952, 380)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd380 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 34
			// srcs: (1953, 381)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd381 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 35
			// srcs: (1954, 382)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd382 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 36
			// srcs: (1955, 383)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd383 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 37
			// srcs: (1957, 384)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd384 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 38
			// srcs: (1958, 385)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd385 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 39
			// srcs: (1960, 386)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd386 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 33
			// srcs: (2023, 387)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd387 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 34
			// srcs: (2026, 388)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd388 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 35
			// srcs: (2029, 389)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd389 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 36
			// srcs: (2032, 390)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd390 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 33
			// srcs: (2033, 391)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd391 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 34
			// srcs: (2034, 392)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd392 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 37
			// srcs: (2035, 393)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd393 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 35
			// srcs: (2036, 394)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd394 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 36
			// srcs: (2037, 395)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd395 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 38
			// srcs: (2038, 396)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd396 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 37
			// srcs: (2039, 397)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd397 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 38
			// srcs: (2040, 398)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd398 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 39
			// srcs: (2041, 399)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd399 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 39
			// srcs: (2042, 400)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd400 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 33
			// srcs: (2113, 401)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd401 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 34
			// srcs: (2114, 402)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd402 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 35
			// srcs: (2116, 403)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd403 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 36
			// srcs: (2117, 404)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd404 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 37
			// srcs: (2119, 405)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd405 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 38
			// srcs: (2120, 406)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd406 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 39
			// srcs: (2122, 407)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd407 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 33
			// srcs: (2195, 408)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd408 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 34
			// srcs: (2196, 409)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd409 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 35
			// srcs: (2197, 410)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd410 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 36
			// srcs: (2198, 411)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd411 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 37
			// srcs: (2199, 412)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd412 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 38
			// srcs: (2200, 413)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd413 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 39
			// srcs: (2202, 414)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd414 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 33
			// srcs: (2207, 415)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd415 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 34
			// srcs: (2210, 416)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd416 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 35
			// srcs: (2213, 417)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd417 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 36
			// srcs: (2216, 418)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd418 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 37
			// srcs: (2219, 419)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd419 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 38
			// srcs: (2222, 420)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd420 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 39
			// srcs: (2225, 421)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd421 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 33
			// srcs: (2275, 422)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd422 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 34
			// srcs: (2276, 423)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd423 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 35
			// srcs: (2278, 424)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd424 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 36
			// srcs: (2279, 425)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd425 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 37
			// srcs: (2281, 426)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd426 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 38
			// srcs: (2282, 427)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd427 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 39
			// srcs: (2284, 428)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd428 : rdata = 48'b110001110000001100000000000000000000000011110000;
			default : rdata = 48'b000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 33) begin
	always @(*) begin
		case(address)
			// PEs: 33, 33 -> 32
			// srcs: (1, 0)(44) -1, (829) 0 --> (1613) 0:ND0, NW0, *, PEGB0
			10'd0 : rdata = 48'b000110110000000001000000000000000000000010000000;
			// PEs: 33, 33 -> 32
			// srcs: (2, 1)(124) -1, (909) 0 --> (1693) 0:ND1, NW1, *, PEGB0
			10'd1 : rdata = 48'b000110110000000101000000001000000000000010000000;
			// PEs: 33, 33 -> 32
			// srcs: (3, 2)(204) 0, (989) 1 --> (1773) 0:ND2, NW2, *, PEGB0
			10'd2 : rdata = 48'b000110110000001001000000010000000000000010000000;
			// PEs: 33, 33 -> 32
			// srcs: (4, 3)(286) 2, (1071) 2 --> (1855) 4:ND3, NW3, *, PEGB0
			10'd3 : rdata = 48'b000110110000001101000000011000000000000010000000;
			// PEs: 33, 33 -> 32
			// srcs: (5, 4)(366) -2, (1151) -2 --> (1935) 4:ND4, NW4, *, PEGB0
			10'd4 : rdata = 48'b000110110000010001000000100000000000000010000000;
			// PEs: 33, 33 -> 33
			// srcs: (6, 5)(447) 1, (1232) 1 --> (2016) 1:ND5, NW5, *, NI0
			10'd5 : rdata = 48'b000110110000010101000000101100000000000000000000;
			// PEs: 33, 33 -> 32
			// srcs: (7, 6)(528) -2, (1313) -3 --> (2097) 6:ND6, NW6, *, PEGB0
			10'd6 : rdata = 48'b000110110000011001000000110000000000000010000000;
			// PEs: 33, 33 -> 32
			// srcs: (8, 7)(608) 0, (1393) -3 --> (2177) 0:ND7, NW7, *, PEGB0
			10'd7 : rdata = 48'b000110110000011101000000111000000000000010000000;
			// PEs: 33, 33 -> 37
			// srcs: (9, 8)(690) 0, (1475) 1 --> (2259) 0:ND8, NW8, *, PEGB5
			10'd8 : rdata = 48'b000110110000100001000001000000000000000011010000;
			// PEs: 33, 33 -> 38
			// srcs: (10, 9)(770) -1, (1555) -1 --> (2339) 1:ND9, NW9, *, PEGB6
			10'd9 : rdata = 48'b000110110000100101000001001000000000000011100000;
			// PEs: 33, 33 -> 33
			// srcs: (11, 10)(150) -2, (935) -3 --> (1719) 6:ND10, NW10, *, NI1
			10'd10 : rdata = 48'b000110110000101001000001010100001000000000000000;
			// PEs: 33, 33 -> 33
			// srcs: (12, 11)(334) -3, (1119) -1 --> (1903) 3:ND11, NW11, *, NI2
			10'd11 : rdata = 48'b000110110000101101000001011100010000000000000000;
			// PEs: 33, 33 -> 33
			// srcs: (13, 12)(518) 2, (1303) -2 --> (2087) -4:ND12, NW12, *, NI3
			10'd12 : rdata = 48'b000110110000110001000001100100011000000000000000;
			// PEs: 33, 33 -> 33
			// srcs: (14, 13)(702) 2, (1487) 2 --> (2271) 4:ND13, NW13, *, NI4
			10'd13 : rdata = 48'b000110110000110101000001101100100000000000000000;
			// PEs: 32 -> 
			// srcs: (34, 14)(1660) 0 --> (1660) 0:PENB, pass, 
			10'd14 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 32, 33 -> 32
			// srcs: (40, 15)(1659) 2, (1660) 0 --> (2440) 2:PENB, ALU, +, PEGB0
			10'd15 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 32 -> 
			// srcs: (50, 16)(1813) 2 --> (1813) 2:PENB, pass, 
			10'd16 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 32, 33 -> 33
			// srcs: (56, 17)(1812) 3, (1813) 2 --> (2592) 5:PENB, ALU, +, NI5
			10'd17 : rdata = 48'b000011101111111000111111111100101000000000000000;
			// PEs: 32 -> 
			// srcs: (75, 18)(1927) -2 --> (1927) -2:PENB, pass, 
			10'd18 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 32, 33 -> 33
			// srcs: (81, 19)(1926) -2, (1927) -2 --> (2705) -4:PENB, ALU, +, NI6
			10'd19 : rdata = 48'b000011101111111000111111111100110000000000000000;
			// PEs: 32 -> 
			// srcs: (84, 20)(1930) -3 --> (1930) -3:PENB, pass, 
			10'd20 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 32, 33 -> 33
			// srcs: (90, 21)(1929) 2, (1930) -3 --> (2709) -1:PENB, ALU, +, NI7
			10'd21 : rdata = 48'b000011101111111000111111111100111000000000000000;
			// PEs: 32 -> 
			// srcs: (92, 22)(1933) 0 --> (1933) 0:PENB, pass, 
			10'd22 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 32, 33 -> 33
			// srcs: (98, 23)(1932) -4, (1933) 0 --> (2711) -4:PENB, ALU, +, NI8
			10'd23 : rdata = 48'b000011101111111000111111111101000000000000000000;
			// PEs: 32 -> 
			// srcs: (100, 24)(2009) -3 --> (2009) -3:PENB, pass, 
			10'd24 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 32, 33 -> 33
			// srcs: (106, 25)(2008) 0, (2009) -3 --> (2788) -3:PENB, ALU, +, NI9
			10'd25 : rdata = 48'b000011101111111000111111111101001000000000000000;
			// PEs: 32 -> 33
			// srcs: (108, 26)(2012) -4 --> (2012) -4:PENB, pass, NI10
			10'd26 : rdata = 48'b110001101111111000000000000101010000000000000000;
			// PEs: 33 -> 32
			// srcs: (111, 42)(2016) 1 --> (2016) 1:NI0, pass, PEGB0
			10'd27 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 32, 33 -> 33
			// srcs: (114, 27)(2011) -6, (2012) -4 --> (2790) -10:PENB, NI10, +, NI0
			10'd28 : rdata = 48'b000011101111111010100001010100000000000000000000;
			// PEs: 32 -> 33
			// srcs: (116, 28)(2089) 0 --> (2089) 0:PENB, pass, NI10
			10'd29 : rdata = 48'b110001101111111000000000000101010000000000000000;
			// PEs: 33 -> 32
			// srcs: (120, 53)(1719) 6 --> (1719) 6:NI1, pass, PEGB0
			10'd30 : rdata = 48'b110001010000000100000000000000000000000010000000;
			// PEs: 33 -> 32
			// srcs: (121, 64)(1903) 3 --> (1903) 3:NI2, pass, PEGB0
			10'd31 : rdata = 48'b110001010000001000000000000000000000000010000000;
			// PEs: 32, 33 -> 34
			// srcs: (122, 29)(2088) -2, (2089) 0 --> (2869) -2:PENB, NI10, +, PENB
			10'd32 : rdata = 48'b000011101111111010100001010000000000000100000000;
			// PEs: 32 -> 
			// srcs: (124, 30)(2092) 0 --> (2092) 0:PENB, pass, 
			10'd33 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 32, 33 -> 39
			// srcs: (130, 31)(2091) 0, (2092) 0 --> (2871) 0:PENB, ALU, +, PEGB7
			10'd34 : rdata = 48'b000011101111111000111111111000000000000011110000;
			// PEs: 32 -> 33
			// srcs: (132, 32)(2095) 0 --> (2095) 0:PENB, pass, NI1
			10'd35 : rdata = 48'b110001101111111000000000000100001000000000000000;
			// PEs: 33 -> 32
			// srcs: (137, 58)(2592) 5 --> (2592) 5:NI5, pass, PEGB0
			10'd36 : rdata = 48'b110001010000010100000000000000000000000010000000;
			// PEs: 32, 33 -> 37
			// srcs: (138, 33)(2094) 4, (2095) 0 --> (2874) 4:PENB, NI1, +, PEGB5
			10'd37 : rdata = 48'b000011101111111010100000001000000000000011010000;
			// PEs: 32 -> 
			// srcs: (140, 34)(2169) -2 --> (2169) -2:PENB, pass, 
			10'd38 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 32, 33 -> 33
			// srcs: (146, 35)(2168) 0, (2169) -2 --> (2949) -2:PENB, ALU, +, NI1
			10'd39 : rdata = 48'b000011101111111000111111111100001000000000000000;
			// PEs: 32 -> 33
			// srcs: (148, 36)(2172) 0 --> (2172) 0:PENB, pass, NI2
			10'd40 : rdata = 48'b110001101111111000000000000100010000000000000000;
			// PEs: 33 -> 32
			// srcs: (151, 67)(2705) -4 --> (2705) -4:NI6, pass, PEGB0
			10'd41 : rdata = 48'b110001010000011000000000000000000000000010000000;
			// PEs: 32, 33 -> 32
			// srcs: (154, 37)(2171) 4, (2172) 0 --> (2951) 4:PENB, NI2, +, PEGB0
			10'd42 : rdata = 48'b000011101111111010100000010000000000000010000000;
			// PEs: 32 -> 33
			// srcs: (156, 38)(2175) 6 --> (2175) 6:PENB, pass, NI2
			10'd43 : rdata = 48'b110001101111111000000000000100010000000000000000;
			// PEs: 33 -> 32
			// srcs: (159, 68)(2709) -1 --> (2709) -1:NI7, pass, PEGB0
			10'd44 : rdata = 48'b110001010000011100000000000000000000000010000000;
			// PEs: 32, 33 -> 33
			// srcs: (162, 39)(2174) 3, (2175) 6 --> (2955) 9:PENB, NI2, +, NI5
			10'd45 : rdata = 48'b000011101111111010100000010100101000000000000000;
			// PEs: 33 -> 32
			// srcs: (167, 69)(2711) -4 --> (2711) -4:NI8, pass, PEGB0
			10'd46 : rdata = 48'b110001010000100000000000000000000000000010000000;
			// PEs: 33 -> 32
			// srcs: (175, 72)(2788) -3 --> (2788) -3:NI9, pass, PEGB0
			10'd47 : rdata = 48'b110001010000100100000000000000000000000010000000;
			// PEs: 33 -> 32
			// srcs: (183, 73)(2790) -10 --> (2790) -10:NI0, pass, PEGB0
			10'd48 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 32 -> 
			// srcs: (290, 40)(2015) 4 --> (2015) 4:PENB, pass, 
			10'd49 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 32, 33 -> 32
			// srcs: (296, 41)(2014) 0, (2015) 4 --> (2796) 4:PENB, ALU, +, PEGB0
			10'd50 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 32 -> 
			// srcs: (298, 43)(1588) 2 --> (1588) 2:PENB, pass, 
			10'd51 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 32, 33 -> 32
			// srcs: (304, 44)(2369) -1, (1588) 2 --> (2370) 1:PENB, ALU, +, PEGB0
			10'd52 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 32 -> 
			// srcs: (306, 45)(1609) 6 --> (1609) 6:PENB, pass, 
			10'd53 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 32, 33 -> 33
			// srcs: (312, 46)(2388) -2, (1609) 6 --> (2389) 4:PENB, ALU, +, NI0
			10'd54 : rdata = 48'b000011101111111000111111111100000000000000000000;
			// PEs: 32 -> 
			// srcs: (314, 47)(1640) -1 --> (1640) -1:PENB, pass, 
			10'd55 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 32, 33 -> 33
			// srcs: (320, 48)(2419) 3, (1640) -1 --> (2420) 2:PENB, ALU, +, NI2
			10'd56 : rdata = 48'b000011101111111000111111111100010000000000000000;
			// PEs: 32 -> 33
			// srcs: (322, 49)(1680) 3 --> (1680) 3:PENB, pass, NI6
			10'd57 : rdata = 48'b110001101111111000000000000100110000000000000000;
			// PEs: 33 -> 32
			// srcs: (324, 81)(2949) -2 --> (2949) -2:NI1, pass, PEGB0
			10'd58 : rdata = 48'b110001010000000100000000000000000000000010000000;
			// PEs: 32, 33 -> 32
			// srcs: (328, 50)(2460) -5, (1680) 3 --> (2461) -2:PENB, NI6, +, PEGB0
			10'd59 : rdata = 48'b000011101111111010100000110000000000000010000000;
			// PEs: 32 -> 33
			// srcs: (330, 51)(1698) -4 --> (1698) -4:PENB, pass, NI1
			10'd60 : rdata = 48'b110001101111111000000000000100001000000000000000;
			// PEs: 33 -> 32
			// srcs: (332, 86)(2271) 4 --> (2271) 4:NI4, pass, PEGB0
			10'd61 : rdata = 48'b110001010000010000000000000000000000000010000000;
			// PEs: 32, 33 -> 32
			// srcs: (336, 52)(2478) 4, (1698) -4 --> (2479) 0:PENB, NI1, +, PEGB0
			10'd62 : rdata = 48'b000011101111111010100000001000000000000010000000;
			// PEs: 32, 37 -> 32
			// srcs: (337, 54)(2514) 3, (1735) -2 --> (2515) 1:PENB, PEGB5, +, PEGB0
			10'd63 : rdata = 48'b000011101111111011100001010000000000000010000000;
			// PEs: 32 -> 
			// srcs: (339, 55)(1750) 0 --> (1750) 0:PENB, pass, 
			10'd64 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 32, 33 -> 33
			// srcs: (345, 56)(2528) -1, (1750) 0 --> (2529) -1:PENB, ALU, +, NI1
			10'd65 : rdata = 48'b000011101111111000111111111100001000000000000000;
			// PEs: 38, 32 -> 32
			// srcs: (346, 57)(2542) 0, (1765) 0 --> (2543) 0:PEGB6, PENB, +, PEGB0
			10'd66 : rdata = 48'b000011110000110011011111110000000000000010000000;
			// PEs: 32 -> 
			// srcs: (348, 59)(1830) 0 --> (1830) 0:PENB, pass, 
			10'd67 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 32, 33 -> 33
			// srcs: (354, 60)(2608) 0, (1830) 0 --> (2609) 0:PENB, ALU, +, NI4
			10'd68 : rdata = 48'b000011101111111000111111111100100000000000000000;
			// PEs: 37, 32 -> 32
			// srcs: (355, 61)(2631) 0, (1854) 0 --> (2632) 0:PEGB5, PENB, +, PEGB0
			10'd69 : rdata = 48'b000011110000101011011111110000000000000010000000;
			// PEs: 32 -> 
			// srcs: (357, 62)(1882) 0 --> (1882) 0:PENB, pass, 
			10'd70 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 32, 33 -> 32
			// srcs: (363, 63)(2661) 0, (1882) 0 --> (2662) 0:PENB, ALU, +, PEGB0
			10'd71 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 32, 35 -> 32
			// srcs: (364, 65)(2686) -3, (1909) -4 --> (2687) -7:PENB, PEGB3, +, PEGB0
			10'd72 : rdata = 48'b000011101111111011100000110000000000000010000000;
			// PEs: 32, 38 -> 33
			// srcs: (372, 66)(2700) 0, (1922) 6 --> (2701) 6:PENB, PEGB6, +, NI6
			10'd73 : rdata = 48'b000011101111111011100001100100110000000000000000;
			// PEs: 32 -> 
			// srcs: (373, 70)(1995) 4 --> (1995) 4:PENB, pass, 
			10'd74 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 32, 33 -> 33
			// srcs: (378, 71)(2774) 0, (1995) 4 --> (2775) 4:PENB, ALU, +, NI7
			10'd75 : rdata = 48'b000011101111111000111111111100111000000000000000;
			// PEs: 32 -> 
			// srcs: (380, 74)(2035) -1 --> (2035) -1:PENB, pass, 
			10'd76 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 32, 33 -> 32
			// srcs: (386, 75)(2813) 10, (2035) -1 --> (2814) 9:PENB, ALU, +, PEGB0
			10'd77 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 32, 33 -> 38
			// srcs: (387, 76)(2864) 3, (2087) -4 --> (2865) -1:PENB, NI3, +, PEGB6
			10'd78 : rdata = 48'b000011101111111010100000011000000000000011100000;
			// PEs: 32 -> 
			// srcs: (389, 77)(2145) 1 --> (2145) 1:PENB, pass, 
			10'd79 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 32, 33 -> 33
			// srcs: (395, 78)(2922) 0, (2145) 1 --> (2923) 1:PENB, ALU, +, NI3
			10'd80 : rdata = 48'b000011101111111000111111111100011000000000000000;
			// PEs: 32 -> 
			// srcs: (397, 79)(2167) -1 --> (2167) -1:PENB, pass, 
			10'd81 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 32, 33 -> 36
			// srcs: (403, 80)(2946) 0, (2167) -1 --> (2947) -1:PENB, ALU, +, PEGB4
			10'd82 : rdata = 48'b000011101111111000111111111000000000000011000000;
			// PEs: 33, 32 -> 32
			// srcs: (404, 82)(2955) 9, (2176) 2 --> (2956) 11:NI5, PENB, +, PEGB0
			10'd83 : rdata = 48'b000011010000010111011111110000000000000010000000;
			// PEs: 32 -> 
			// srcs: (406, 83)(2182) -3 --> (2182) -3:PENB, pass, 
			10'd84 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 32, 33 -> 32
			// srcs: (412, 84)(2960) 2, (2182) -3 --> (2961) -1:PENB, ALU, +, PEGB0
			10'd85 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 39, 32 -> 39
			// srcs: (413, 85)(3043) -5, (2265) 2 --> (3044) -3:PEGB7, PENB, +, PEGB7
			10'd86 : rdata = 48'b000011110000111011011111110000000000000011110000;
			// PEs: 32, 38 -> 32
			// srcs: (421, 87)(3064) -2, (2286) -1 --> (3065) -3:PENB, PEGB6, +, PEGB0
			10'd87 : rdata = 48'b000011101111111011100001100000000000000010000000;
			// PEs: 32 -> 
			// srcs: (422, 88)(2298) 0 --> (2298) 0:PENB, pass, 
			10'd88 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 32, 33 -> 32
			// srcs: (427, 89)(3075) 4, (2298) 0 --> (3076) 4:PENB, ALU, +, PEGB0
			10'd89 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 32 -> 
			// srcs: (429, 90)(2323) 2 --> (2323) 2:PENB, pass, 
			10'd90 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 32, 33 -> 32
			// srcs: (435, 91)(3100) 2, (2323) 2 --> (3101) 4:PENB, ALU, +, PEGB0
			10'd91 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 32 -> 
			// srcs: (564, 92)(2350) -3 --> (2350) -3:PENB, pass, 
			10'd92 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 32, 33 -> 33
			// srcs: (570, 93)(3125) -2, (2350) -3 --> (3126) -5:PENB, ALU, +, NI5
			10'd93 : rdata = 48'b000011101111111000111111111100101000000000000000;
			// PEs: 32, 33 -> 32
			// srcs: (571, 94)(2387) 3, (2389) 4 --> (2390) 7:PENB, NI0, +, PEGB0
			10'd94 : rdata = 48'b000011101111111010100000000000000000000010000000;
			// PEs: 32, 33 -> 32
			// srcs: (572, 95)(2418) -1, (2420) 2 --> (2421) 1:PENB, NI2, +, PEGB0
			10'd95 : rdata = 48'b000011101111111010100000010000000000000010000000;
			// PEs: 32 -> 
			// srcs: (574, 96)(2437) 5 --> (2437) 5:PENB, pass, 
			10'd96 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 32, 33 -> 33
			// srcs: (580, 97)(2435) 2, (2437) 5 --> (2438) 7:PENB, ALU, +, NI0
			10'd97 : rdata = 48'b000011101111111000111111111100000000000000000000;
			// PEs: 32 -> 
			// srcs: (582, 98)(2506) 14 --> (2506) 14:PENB, pass, 
			10'd98 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 32, 33 -> 32
			// srcs: (588, 99)(2504) 1, (2506) 14 --> (2507) 15:PENB, ALU, +, PEGB0
			10'd99 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 32, 33 -> 32
			// srcs: (589, 100)(2527) 0, (2529) -1 --> (2530) -1:PENB, NI1, +, PEGB0
			10'd100 : rdata = 48'b000011101111111010100000001000000000000010000000;
			// PEs: 32, 33 -> 33
			// srcs: (590, 101)(2607) 2, (2609) 0 --> (2610) 2:PENB, NI4, +, NI1
			10'd101 : rdata = 48'b000011101111111010100000100100001000000000000000;
			// PEs: 32 -> 
			// srcs: (592, 102)(2658) 2 --> (2658) 2:PENB, pass, 
			10'd102 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 32, 33 -> 32
			// srcs: (598, 103)(2656) -4, (2658) 2 --> (2659) -2:PENB, ALU, +, PEGB0
			10'd103 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 32, 33 -> 32
			// srcs: (599, 104)(2699) 7, (2701) 6 --> (2702) 13:PENB, NI6, +, PEGB0
			10'd104 : rdata = 48'b000011101111111010100000110000000000000010000000;
			// PEs: 32, 33 -> 33
			// srcs: (602, 105)(2773) 3, (2775) 4 --> (2776) 7:PENB, NI7, +, NI2
			10'd105 : rdata = 48'b000011101111111010100000111100010000000000000000;
			// PEs: 32 -> 
			// srcs: (610, 106)(2823) 5 --> (2823) 5:PENB, pass, 
			10'd106 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 32, 33 -> 32
			// srcs: (619, 107)(2821) 5, (2823) 5 --> (2824) 10:PENB, ALU, +, PEGB0
			10'd107 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 33, 32 -> 32
			// srcs: (620, 108)(2923) 1, (2925) -3 --> (2926) -2:NI3, PENB, +, PEGB0
			10'd108 : rdata = 48'b000011010000001111011111110000000000000010000000;
			// PEs: 32 -> 
			// srcs: (622, 109)(2975) 0 --> (2975) 0:PENB, pass, 
			10'd109 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 32, 33 -> 33
			// srcs: (628, 110)(2973) -10, (2975) 0 --> (2976) -10:PENB, ALU, +, NI3
			10'd110 : rdata = 48'b000011101111111000111111111100011000000000000000;
			// PEs: 32 -> 
			// srcs: (630, 111)(3072) 0 --> (3072) 0:PENB, pass, 
			10'd111 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 32, 33 -> 33
			// srcs: (636, 112)(3070) 4, (3072) 0 --> (3073) 4:PENB, ALU, +, NI4
			10'd112 : rdata = 48'b000011101111111000111111111100100000000000000000;
			// PEs: 32, 33 -> 37
			// srcs: (1100, 113)(3124) 9, (3126) -5 --> (3127) 4:PENB, NI5, +, PEGB5
			10'd113 : rdata = 48'b000011101111111010100000101000000000000011010000;
			// PEs: 32 -> 
			// srcs: (1102, 114)(2415) -3 --> (2415) -3:PENB, pass, 
			10'd114 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 32, 33 -> 32
			// srcs: (1108, 115)(2410) 6, (2415) -3 --> (2416) 3:PENB, ALU, +, PEGB0
			10'd115 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 32, 33 -> 32
			// srcs: (1109, 116)(2433) 3, (2438) 7 --> (2439) 10:PENB, NI0, +, PEGB0
			10'd116 : rdata = 48'b000011101111111010100000000000000000000010000000;
			// PEs: 32, 33 -> 32
			// srcs: (1110, 117)(2605) 16, (2610) 2 --> (2611) 18:PENB, NI1, +, PEGB0
			10'd117 : rdata = 48'b000011101111111010100000001000000000000010000000;
			// PEs: 33, 32 -> 33
			// srcs: (1111, 118)(2776) 7, (2781) 5 --> (2782) 12:NI2, PENB, +, NI0
			10'd118 : rdata = 48'b000011010000001011011111110100000000000000000000;
			// PEs: 32 -> 
			// srcs: (1113, 119)(2792) -13 --> (2792) -13:PENB, pass, 
			10'd119 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 32, 33 -> 34
			// srcs: (1119, 120)(2787) 0, (2792) -13 --> (2793) -13:PENB, ALU, +, PENB
			10'd120 : rdata = 48'b000011101111111000111111111000000000000100000000;
			// PEs: 32, 33 -> 32
			// srcs: (1120, 121)(2971) 7, (2976) -10 --> (2977) -3:PENB, NI3, +, PEGB0
			10'd121 : rdata = 48'b000011101111111010100000011000000000000010000000;
			// PEs: 32, 33 -> 32
			// srcs: (1121, 122)(3068) -5, (3073) 4 --> (3074) -1:PENB, NI4, +, PEGB0
			10'd122 : rdata = 48'b000011101111111010100000100000000000000010000000;
			// PEs: 32 -> 33
			// srcs: (1123, 123)(2402) -10 --> (2402) -10:PENB, pass, NI1
			10'd123 : rdata = 48'b110001101111111000000000000100001000000000000000;
			// PEs: 33 -> 34
			// srcs: (1126, 127)(2782) 12 --> (2782) 12:NI0, pass, PENB
			10'd124 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 32, 33 -> 32
			// srcs: (1129, 124)(2391) 4, (2402) -10 --> (2403) -6:PENB, NI1, +, PEGB0
			10'd125 : rdata = 48'b000011101111111010100000001000000000000010000000;
			// PEs: 32 -> 
			// srcs: (1131, 125)(2645) 2 --> (2645) 2:PENB, pass, 
			10'd126 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 32, 33 -> 32
			// srcs: (1137, 126)(2634) 19, (2645) 2 --> (2646) 21:PENB, ALU, +, PEGB0
			10'd127 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 32 -> 
			// srcs: (1139, 128)(2548) -21 --> (2548) -21:PENB, pass, 
			10'd128 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 32, 33 -> 32
			// srcs: (1145, 129)(2525) 19, (2548) -21 --> (2549) -2:PENB, ALU, +, PEGB0
			10'd129 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 32 -> 
			// srcs: (1409, 130)(2939) 11 --> (2939) 11:PENB, pass, 
			10'd130 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 32, 33 -> 32
			// srcs: (1416, 131)(2916) 16, (2939) 11 --> (2940) 27:PENB, ALU, +, PEGB0
			10'd131 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 32 -> 
			// srcs: (1431, 132)(3038) -37 --> (3038) -37:PENB, pass, 
			10'd132 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 32, 33 -> 32
			// srcs: (1437, 133)(2990) -1, (3038) -37 --> (3039) -38:PENB, ALU, +, PEGB0
			10'd133 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 32, 33 -> 34
			// srcs: (1551, 134)(3140) 47, (44) -1 --> (3181) -47:PENB, ND0, *, PENB
			10'd134 : rdata = 48'b000111101111111001100000000000000000000100000000;
			// PEs: 33, 34 -> 33
			// srcs: (1560, 148)(829) 0, (3965) -47 --> (4749) 47:NW0, PEGB2, -, NW0
			10'd135 : rdata = 48'b000100100000000011100000100000000100000000000000;
			// PEs: 32, 33 -> 34
			// srcs: (1631, 135)(3140) 47, (124) -1 --> (3261) -47:PENB, ND1, *, PENB
			10'd136 : rdata = 48'b000111101111111001100000001000000000000100000000;
			// PEs: 33, 34 -> 33
			// srcs: (1640, 149)(909) 0, (4045) -47 --> (4829) 47:NW1, PEGB2, -, NW1
			10'd137 : rdata = 48'b000100100000000111100000100000000100010000000000;
			// PEs: 32, 33 -> 34
			// srcs: (1657, 136)(3140) 47, (150) -2 --> (3287) -94:PENB, ND10, *, PENB
			10'd138 : rdata = 48'b000111101111111001100001010000000000000100000000;
			// PEs: 33, 34 -> 33
			// srcs: (1666, 150)(935) -3, (4071) -94 --> (4855) 91:NW10, PEGB2, -, NW10
			10'd139 : rdata = 48'b000100100000101011100000100000000110100000000000;
			// PEs: 32, 33 -> 34
			// srcs: (1711, 137)(3140) 47, (204) 0 --> (3341) 0:PENB, ND2, *, PENB
			10'd140 : rdata = 48'b000111101111111001100000010000000000000100000000;
			// PEs: 33, 34 -> 33
			// srcs: (1720, 151)(989) 1, (4125) 0 --> (4909) 1:NW2, PEGB2, -, NW2
			10'd141 : rdata = 48'b000100100000001011100000100000000100100000000000;
			// PEs: 32, 33 -> 34
			// srcs: (1793, 138)(3140) 47, (286) 2 --> (3423) 94:PENB, ND3, *, PENB
			10'd142 : rdata = 48'b000111101111111001100000011000000000000100000000;
			// PEs: 33, 34 -> 33
			// srcs: (1802, 152)(1071) 2, (4207) 94 --> (4991) -92:NW3, PEGB2, -, NW3
			10'd143 : rdata = 48'b000100100000001111100000100000000100110000000000;
			// PEs: 32, 33 -> 34
			// srcs: (1841, 139)(3140) 47, (334) -3 --> (3471) -141:PENB, ND11, *, PENB
			10'd144 : rdata = 48'b000111101111111001100001011000000000000100000000;
			// PEs: 33, 34 -> 33
			// srcs: (1850, 153)(1119) -1, (4255) -141 --> (5039) 140:NW11, PEGB2, -, NW11
			10'd145 : rdata = 48'b000100100000101111100000100000000110110000000000;
			// PEs: 32, 33 -> 34
			// srcs: (1873, 140)(3140) 47, (366) -2 --> (3503) -94:PENB, ND4, *, PENB
			10'd146 : rdata = 48'b000111101111111001100000100000000000000100000000;
			// PEs: 33, 34 -> 33
			// srcs: (1882, 154)(1151) -2, (4287) -94 --> (5071) 92:NW4, PEGB2, -, NW4
			10'd147 : rdata = 48'b000100100000010011100000100000000101000000000000;
			// PEs: 32, 33 -> 34
			// srcs: (1954, 141)(3140) 47, (447) 1 --> (3584) 47:PENB, ND5, *, PENB
			10'd148 : rdata = 48'b000111101111111001100000101000000000000100000000;
			// PEs: 33, 34 -> 33
			// srcs: (1963, 155)(1232) 1, (4368) 47 --> (5152) -46:NW5, PEGB2, -, NW5
			10'd149 : rdata = 48'b000100100000010111100000100000000101010000000000;
			// PEs: 32, 33 -> 34
			// srcs: (2025, 142)(3140) 47, (518) 2 --> (3655) 94:PENB, ND12, *, PENB
			10'd150 : rdata = 48'b000111101111111001100001100000000000000100000000;
			// PEs: 33, 34 -> 33
			// srcs: (2034, 156)(1303) -2, (4439) 94 --> (5223) -96:NW12, PEGB2, -, NW12
			10'd151 : rdata = 48'b000100100000110011100000100000000111000000000000;
			// PEs: 32, 33 -> 34
			// srcs: (2035, 143)(3140) 47, (528) -2 --> (3665) -94:PENB, ND6, *, PENB
			10'd152 : rdata = 48'b000111101111111001100000110000000000000100000000;
			// PEs: 33, 34 -> 33
			// srcs: (2044, 157)(1313) -3, (4449) -94 --> (5233) 91:NW6, PEGB2, -, NW6
			10'd153 : rdata = 48'b000100100000011011100000100000000101100000000000;
			// PEs: 32, 33 -> 34
			// srcs: (2115, 144)(3140) 47, (608) 0 --> (3745) 0:PENB, ND7, *, PENB
			10'd154 : rdata = 48'b000111101111111001100000111000000000000100000000;
			// PEs: 33, 34 -> 33
			// srcs: (2124, 158)(1393) -3, (4529) 0 --> (5313) -3:NW7, PEGB2, -, NW7
			10'd155 : rdata = 48'b000100100000011111100000100000000101110000000000;
			// PEs: 32, 33 -> 34
			// srcs: (2197, 145)(3140) 47, (690) 0 --> (3827) 0:PENB, ND8, *, PENB
			10'd156 : rdata = 48'b000111101111111001100001000000000000000100000000;
			// PEs: 33, 34 -> 33
			// srcs: (2206, 159)(1475) 1, (4611) 0 --> (5395) 1:NW8, PEGB2, -, NW8
			10'd157 : rdata = 48'b000100100000100011100000100000000110000000000000;
			// PEs: 32, 33 -> 34
			// srcs: (2209, 146)(3140) 47, (702) 2 --> (3839) 94:PENB, ND13, *, PENB
			10'd158 : rdata = 48'b000111101111111001100001101000000000000100000000;
			// PEs: 33, 34 -> 33
			// srcs: (2218, 160)(1487) 2, (4623) 94 --> (5407) -92:NW13, PEGB2, -, NW13
			10'd159 : rdata = 48'b000100100000110111100000100000000111010000000000;
			// PEs: 32, 33 -> 34
			// srcs: (2277, 147)(3140) 47, (770) -1 --> (3907) -47:PENB, ND9, *, PENB
			10'd160 : rdata = 48'b000111101111111001100001001000000000000100000000;
			// PEs: 33, 34 -> 33
			// srcs: (2286, 161)(1555) -1, (4691) -47 --> (5475) 46:NW9, PEGB2, -, NW9
			10'd161 : rdata = 48'b000100100000100111100000100000000110010000000000;
			default : rdata = 48'b000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 34) begin
	always @(*) begin
		case(address)
			// PEs: 34, 34 -> 32
			// srcs: (1, 0)(45) -2, (830) -3 --> (1614) 6:ND0, NW0, *, PEGB0
			10'd0 : rdata = 48'b000110110000000001000000000000000000000010000000;
			// PEs: 34, 34 -> 32
			// srcs: (2, 1)(125) -3, (910) 2 --> (1694) -6:ND1, NW1, *, PEGB0
			10'd1 : rdata = 48'b000110110000000101000000001000000000000010000000;
			// PEs: 34, 34 -> 32
			// srcs: (3, 2)(205) -1, (990) -1 --> (1774) 1:ND2, NW2, *, PEGB0
			10'd2 : rdata = 48'b000110110000001001000000010000000000000010000000;
			// PEs: 34, 34 -> 32
			// srcs: (4, 3)(287) 0, (1072) -2 --> (1856) 0:ND3, NW3, *, PEGB0
			10'd3 : rdata = 48'b000110110000001101000000011000000000000010000000;
			// PEs: 34, 34 -> 32
			// srcs: (5, 4)(367) 1, (1152) -3 --> (1936) -3:ND4, NW4, *, PEGB0
			10'd4 : rdata = 48'b000110110000010001000000100000000000000010000000;
			// PEs: 34, 34 -> 34
			// srcs: (6, 5)(448) 0, (1233) 0 --> (2017) 0:ND5, NW5, *, NI0
			10'd5 : rdata = 48'b000110110000010101000000101100000000000000000000;
			// PEs: 34, 34 -> 32
			// srcs: (7, 6)(529) 0, (1314) -1 --> (2098) 0:ND6, NW6, *, PEGB0
			10'd6 : rdata = 48'b000110110000011001000000110000000000000010000000;
			// PEs: 34, 34 -> 32
			// srcs: (8, 7)(609) -1, (1394) -3 --> (2178) 3:ND7, NW7, *, PEGB0
			10'd7 : rdata = 48'b000110110000011101000000111000000000000010000000;
			// PEs: 34, 34 -> 37
			// srcs: (9, 8)(691) 1, (1476) -1 --> (2260) -1:ND8, NW8, *, PEGB5
			10'd8 : rdata = 48'b000110110000100001000001000000000000000011010000;
			// PEs: 34, 34 -> 38
			// srcs: (10, 9)(771) 1, (1556) -2 --> (2340) -2:ND9, NW9, *, PEGB6
			10'd9 : rdata = 48'b000110110000100101000001001000000000000011100000;
			// PEs: 34, 34 -> 34
			// srcs: (11, 10)(157) -3, (942) -2 --> (1726) 6:ND10, NW10, *, NI1
			10'd10 : rdata = 48'b000110110000101001000001010100001000000000000000;
			// PEs: 34, 34 -> 34
			// srcs: (12, 11)(337) -3, (1122) -2 --> (1906) 6:ND11, NW11, *, NI2
			10'd11 : rdata = 48'b000110110000101101000001011100010000000000000000;
			// PEs: 34, 34 -> 34
			// srcs: (13, 12)(521) 1, (1306) -2 --> (2090) -2:ND12, NW12, *, NI3
			10'd12 : rdata = 48'b000110110000110001000001100100011000000000000000;
			// PEs: 34, 34 -> 34
			// srcs: (14, 13)(705) -2, (1490) -2 --> (2274) 4:ND13, NW13, *, NI4
			10'd13 : rdata = 48'b000110110000110101000001101100100000000000000000;
			// PEs: 38 -> 
			// srcs: (15, 18)(2346) 1 --> (2346) 1:PEGB6, pass, 
			10'd14 : rdata = 48'b110001110000110000000000000000000000000000000000;
			// PEs: 37, 34 -> 34
			// srcs: (18, 19)(2345) 6, (2346) 1 --> (3123) 7:PEGB5, ALU, +, NI5
			10'd15 : rdata = 48'b000011110000101000111111111100101000000000000000;
			// PEs: 32 -> 
			// srcs: (48, 14)(1681) 3 --> (1681) 3:PEGB0, pass, 
			10'd16 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 34, 32 -> 32
			// srcs: (57, 15)(1681) 3, (1682) -2 --> (2462) 1:ALU, PEGB0, +, PEGB0
			10'd17 : rdata = 48'b000010011111111111100000000000000000000010000000;
			// PEs: 32 -> 
			// srcs: (70, 16)(1844) 9 --> (1844) 9:PEGB0, pass, 
			10'd18 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 32, 34 -> 34
			// srcs: (79, 17)(1843) 1, (1844) 9 --> (2624) 10:PEGB0, ALU, +, NI6
			10'd19 : rdata = 48'b000011110000000000111111111100110000000000000000;
			// PEs: 34 -> 32
			// srcs: (119, 20)(2017) 0 --> (2017) 0:NI0, pass, PEGB0
			10'd20 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 34 -> 32
			// srcs: (120, 21)(1726) 6 --> (1726) 6:NI1, pass, PEGB0
			10'd21 : rdata = 48'b110001010000000100000000000000000000000010000000;
			// PEs: 33, 34 -> 35
			// srcs: (125, 24)(2869) -2, (2090) -2 --> (2870) -4:PENB, NI3, +, PENB
			10'd22 : rdata = 48'b000011101111111010100000011000000000000100000000;
			// PEs: 34 -> 32
			// srcs: (137, 22)(2624) 10 --> (2624) 10:NI6, pass, PEGB0
			10'd23 : rdata = 48'b110001010000011000000000000000000000000010000000;
			// PEs: 34 -> 32
			// srcs: (158, 23)(1906) 6 --> (1906) 6:NI2, pass, PEGB0
			10'd24 : rdata = 48'b110001010000001000000000000000000000000010000000;
			// PEs: 34 -> 32
			// srcs: (160, 26)(3123) 7 --> (3123) 7:NI5, pass, PEGB0
			10'd25 : rdata = 48'b110001010000010100000000000000000000000010000000;
			// PEs: 34 -> 32
			// srcs: (341, 25)(2274) 4 --> (2274) 4:NI4, pass, PEGB0
			10'd26 : rdata = 48'b110001010000010000000000000000000000000010000000;
			// PEs: 33 -> 
			// srcs: (1121, 27)(2793) -13 --> (2793) -13:PENB, pass, 
			10'd27 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 33, 34 -> 32
			// srcs: (1128, 28)(2782) 12, (2793) -13 --> (2794) -1:PENB, ALU, +, PEGB0
			10'd28 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 34, 33 -> 33
			// srcs: (1554, 43)(3) 1, (3181) -47 --> (3965) -47:NM0, PENB, *, PEGB1
			10'd29 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 32, 34 -> 35
			// srcs: (1555, 29)(3140) 47, (45) -2 --> (3182) -94:PEGB0, ND0, *, PENB
			10'd30 : rdata = 48'b000111110000000001100000000000000000000100000000;
			// PEs: 34, 35 -> 34
			// srcs: (1564, 61)(830) -3, (3966) -94 --> (4750) 91:NW0, PEGB3, -, NW0
			10'd31 : rdata = 48'b000100100000000011100000110000000100000000000000;
			// PEs: 34, 33 -> 33
			// srcs: (1634, 44)(3) 1, (3261) -47 --> (4045) -47:NM0, PENB, *, PEGB1
			10'd32 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 32, 34 -> 35
			// srcs: (1635, 30)(3140) 47, (125) -3 --> (3262) -141:PEGB0, ND1, *, PENB
			10'd33 : rdata = 48'b000111110000000001100000001000000000000100000000;
			// PEs: 34, 35 -> 34
			// srcs: (1644, 62)(910) 2, (4046) -141 --> (4830) 143:NW1, PEGB3, -, NW1
			10'd34 : rdata = 48'b000100100000000111100000110000000100010000000000;
			// PEs: 34, 33 -> 33
			// srcs: (1660, 45)(3) 1, (3287) -94 --> (4071) -94:NM0, PENB, *, PEGB1
			10'd35 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 32, 34 -> 
			// srcs: (1667, 31)(3140) 47, (157) -3 --> (3294) -141:PEGB0, ND10, *, 
			10'd36 : rdata = 48'b000111110000000001100001010000000000000000000000;
			// PEs: 34, 34 -> 
			// srcs: (1670, 46)(3) 1, (3294) -141 --> (4078) -141:NM0, ALU, *, 
			10'd37 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 34, 34 -> 34
			// srcs: (1673, 63)(942) -2, (4078) -141 --> (4862) 139:NW10, ALU, -, NW10
			10'd38 : rdata = 48'b000100100000101000111111111000000110100000000000;
			// PEs: 34, 33 -> 33
			// srcs: (1714, 47)(3) 1, (3341) 0 --> (4125) 0:NM0, PENB, *, PEGB1
			10'd39 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 32, 34 -> 35
			// srcs: (1715, 32)(3140) 47, (205) -1 --> (3342) -47:PEGB0, ND2, *, PENB
			10'd40 : rdata = 48'b000111110000000001100000010000000000000100000000;
			// PEs: 34, 35 -> 34
			// srcs: (1724, 64)(990) -1, (4126) -47 --> (4910) 46:NW2, PEGB3, -, NW2
			10'd41 : rdata = 48'b000100100000001011100000110000000100100000000000;
			// PEs: 34, 33 -> 33
			// srcs: (1796, 48)(3) 1, (3423) 94 --> (4207) 94:NM0, PENB, *, PEGB1
			10'd42 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 32, 34 -> 35
			// srcs: (1797, 33)(3140) 47, (287) 0 --> (3424) 0:PEGB0, ND3, *, PENB
			10'd43 : rdata = 48'b000111110000000001100000011000000000000100000000;
			// PEs: 34, 35 -> 34
			// srcs: (1806, 65)(1072) -2, (4208) 0 --> (4992) -2:NW3, PEGB3, -, NW3
			10'd44 : rdata = 48'b000100100000001111100000110000000100110000000000;
			// PEs: 34, 33 -> 33
			// srcs: (1844, 49)(3) 1, (3471) -141 --> (4255) -141:NM0, PENB, *, PEGB1
			10'd45 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 32, 34 -> 
			// srcs: (1847, 34)(3140) 47, (337) -3 --> (3474) -141:PEGB0, ND11, *, 
			10'd46 : rdata = 48'b000111110000000001100001011000000000000000000000;
			// PEs: 34, 34 -> 
			// srcs: (1850, 50)(3) 1, (3474) -141 --> (4258) -141:NM0, ALU, *, 
			10'd47 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 34, 34 -> 34
			// srcs: (1853, 66)(1122) -2, (4258) -141 --> (5042) 139:NW11, ALU, -, NW11
			10'd48 : rdata = 48'b000100100000101100111111111000000110110000000000;
			// PEs: 34, 33 -> 33
			// srcs: (1876, 51)(3) 1, (3503) -94 --> (4287) -94:NM0, PENB, *, PEGB1
			10'd49 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 32, 34 -> 35
			// srcs: (1877, 35)(3140) 47, (367) 1 --> (3504) 47:PEGB0, ND4, *, PENB
			10'd50 : rdata = 48'b000111110000000001100000100000000000000100000000;
			// PEs: 34, 35 -> 34
			// srcs: (1886, 67)(1152) -3, (4288) 47 --> (5072) -50:NW4, PEGB3, -, NW4
			10'd51 : rdata = 48'b000100100000010011100000110000000101000000000000;
			// PEs: 34, 33 -> 33
			// srcs: (1957, 52)(3) 1, (3584) 47 --> (4368) 47:NM0, PENB, *, PEGB1
			10'd52 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 32, 34 -> 35
			// srcs: (1958, 36)(3140) 47, (448) 0 --> (3585) 0:PEGB0, ND5, *, PENB
			10'd53 : rdata = 48'b000111110000000001100000101000000000000100000000;
			// PEs: 34, 35 -> 34
			// srcs: (1967, 68)(1233) 0, (4369) 0 --> (5153) 0:NW5, PEGB3, -, NW5
			10'd54 : rdata = 48'b000100100000010111100000110000000101010000000000;
			// PEs: 34, 33 -> 33
			// srcs: (2028, 53)(3) 1, (3655) 94 --> (4439) 94:NM0, PENB, *, PEGB1
			10'd55 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 32, 34 -> 
			// srcs: (2031, 37)(3140) 47, (521) 1 --> (3658) 47:PEGB0, ND12, *, 
			10'd56 : rdata = 48'b000111110000000001100001100000000000000000000000;
			// PEs: 34, 34 -> 
			// srcs: (2034, 54)(3) 1, (3658) 47 --> (4442) 47:NM0, ALU, *, 
			10'd57 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 34, 34 -> 34
			// srcs: (2037, 69)(1306) -2, (4442) 47 --> (5226) -49:NW12, ALU, -, NW12
			10'd58 : rdata = 48'b000100100000110000111111111000000111000000000000;
			// PEs: 34, 33 -> 33
			// srcs: (2038, 55)(3) 1, (3665) -94 --> (4449) -94:NM0, PENB, *, PEGB1
			10'd59 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 32, 34 -> 35
			// srcs: (2039, 38)(3140) 47, (529) 0 --> (3666) 0:PEGB0, ND6, *, PENB
			10'd60 : rdata = 48'b000111110000000001100000110000000000000100000000;
			// PEs: 34, 35 -> 34
			// srcs: (2048, 70)(1314) -1, (4450) 0 --> (5234) -1:NW6, PEGB3, -, NW6
			10'd61 : rdata = 48'b000100100000011011100000110000000101100000000000;
			// PEs: 34, 33 -> 33
			// srcs: (2118, 56)(3) 1, (3745) 0 --> (4529) 0:NM0, PENB, *, PEGB1
			10'd62 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 32, 34 -> 35
			// srcs: (2119, 39)(3140) 47, (609) -1 --> (3746) -47:PEGB0, ND7, *, PENB
			10'd63 : rdata = 48'b000111110000000001100000111000000000000100000000;
			// PEs: 34, 35 -> 34
			// srcs: (2128, 71)(1394) -3, (4530) -47 --> (5314) 44:NW7, PEGB3, -, NW7
			10'd64 : rdata = 48'b000100100000011111100000110000000101110000000000;
			// PEs: 34, 33 -> 33
			// srcs: (2200, 57)(3) 1, (3827) 0 --> (4611) 0:NM0, PENB, *, PEGB1
			10'd65 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 32, 34 -> 35
			// srcs: (2201, 40)(3140) 47, (691) 1 --> (3828) 47:PEGB0, ND8, *, PENB
			10'd66 : rdata = 48'b000111110000000001100001000000000000000100000000;
			// PEs: 34, 35 -> 34
			// srcs: (2210, 72)(1476) -1, (4612) 47 --> (5396) -48:NW8, PEGB3, -, NW8
			10'd67 : rdata = 48'b000100100000100011100000110000000110000000000000;
			// PEs: 34, 33 -> 33
			// srcs: (2212, 58)(3) 1, (3839) 94 --> (4623) 94:NM0, PENB, *, PEGB1
			10'd68 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 32, 34 -> 
			// srcs: (2215, 41)(3140) 47, (705) -2 --> (3842) -94:PEGB0, ND13, *, 
			10'd69 : rdata = 48'b000111110000000001100001101000000000000000000000;
			// PEs: 34, 34 -> 
			// srcs: (2218, 59)(3) 1, (3842) -94 --> (4626) -94:NM0, ALU, *, 
			10'd70 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 34, 34 -> 34
			// srcs: (2221, 73)(1490) -2, (4626) -94 --> (5410) 92:NW13, ALU, -, NW13
			10'd71 : rdata = 48'b000100100000110100111111111000000111010000000000;
			// PEs: 34, 33 -> 33
			// srcs: (2280, 60)(3) 1, (3907) -47 --> (4691) -47:NM0, PENB, *, PEGB1
			10'd72 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 32, 34 -> 35
			// srcs: (2281, 42)(3140) 47, (771) 1 --> (3908) 47:PEGB0, ND9, *, PENB
			10'd73 : rdata = 48'b000111110000000001100001001000000000000100000000;
			// PEs: 34, 35 -> 34
			// srcs: (2290, 74)(1556) -2, (4692) 47 --> (5476) -49:NW9, PEGB3, -, NW9
			10'd74 : rdata = 48'b000100100000100111100000110000000110010000000000;
			default : rdata = 48'b000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 35) begin
	always @(*) begin
		case(address)
			// PEs: 35, 35 -> 32
			// srcs: (1, 0)(47) 2, (832) 0 --> (1616) 0:ND0, NW0, *, PEGB0
			10'd0 : rdata = 48'b000110110000000001000000000000000000000010000000;
			// PEs: 35, 35 -> 32
			// srcs: (2, 1)(127) -1, (912) -2 --> (1696) 2:ND1, NW1, *, PEGB0
			10'd1 : rdata = 48'b000110110000000101000000001000000000000010000000;
			// PEs: 35, 35 -> 32
			// srcs: (3, 2)(207) -3, (992) -3 --> (1776) 9:ND2, NW2, *, PEGB0
			10'd2 : rdata = 48'b000110110000001001000000010000000000000010000000;
			// PEs: 35, 35 -> 32
			// srcs: (4, 3)(289) -2, (1074) -1 --> (1858) 2:ND3, NW3, *, PEGB0
			10'd3 : rdata = 48'b000110110000001101000000011000000000000010000000;
			// PEs: 35, 35 -> 32
			// srcs: (5, 4)(369) -1, (1154) 2 --> (1938) -2:ND4, NW4, *, PEGB0
			10'd4 : rdata = 48'b000110110000010001000000100000000000000010000000;
			// PEs: 35, 35 -> 32
			// srcs: (6, 5)(449) -1, (1234) 2 --> (2018) -2:ND5, NW5, *, PEGB0
			10'd5 : rdata = 48'b000110110000010101000000101000000000000010000000;
			// PEs: 35, 35 -> 32
			// srcs: (7, 6)(531) -3, (1316) 1 --> (2100) -3:ND6, NW6, *, PEGB0
			10'd6 : rdata = 48'b000110110000011001000000110000000000000010000000;
			// PEs: 35, 35 -> 32
			// srcs: (8, 7)(611) 1, (1396) 0 --> (2180) 0:ND7, NW7, *, PEGB0
			10'd7 : rdata = 48'b000110110000011101000000111000000000000010000000;
			// PEs: 35, 35 -> 35
			// srcs: (9, 8)(692) 2, (1477) -3 --> (2261) -6:ND8, NW8, *, NI0
			10'd8 : rdata = 48'b000110110000100001000001000100000000000000000000;
			// PEs: 35, 35 -> 39
			// srcs: (10, 9)(773) -2, (1558) 2 --> (2342) -4:ND9, NW9, *, PEGB7
			10'd9 : rdata = 48'b000110110000100101000001001000000000000011110000;
			// PEs: 35, 35 -> 35
			// srcs: (11, 10)(160) 1, (945) -3 --> (1729) -3:ND10, NW10, *, NI1
			10'd10 : rdata = 48'b000110110000101001000001010100001000000000000000;
			// PEs: 35, 35 -> 33
			// srcs: (12, 11)(340) -2, (1125) 2 --> (1909) -4:ND11, NW11, *, PEGB1
			10'd11 : rdata = 48'b000110110000101101000001011000000000000010010000;
			// PEs: 35, 35 -> 39
			// srcs: (13, 12)(524) 2, (1309) 1 --> (2093) 2:ND12, NW12, *, PEGB7
			10'd12 : rdata = 48'b000110110000110001000001100000000000000011110000;
			// PEs: 35, 35 -> 35
			// srcs: (14, 13)(708) 0, (1493) -2 --> (2277) 0:ND13, NW13, *, NI2
			10'd13 : rdata = 48'b000110110000110101000001101100010000000000000000;
			// PEs: 35, 36 -> 38
			// srcs: (15, 20)(2261) -6, (2262) 1 --> (3041) -5:NI0, PEGB4, +, PEGB6
			10'd14 : rdata = 48'b000011010000000011100001000000000000000011100000;
			// PEs: 32 -> 
			// srcs: (41, 14)(1685) 0 --> (1685) 0:PEGB0, pass, 
			10'd15 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 32, 35 -> 32
			// srcs: (50, 15)(1684) 1, (1685) 0 --> (2466) 1:PEGB0, ALU, +, PEGB0
			10'd16 : rdata = 48'b000011110000000000111111111000000000000010000000;
			// PEs: 32 -> 
			// srcs: (72, 16)(1847) 0 --> (1847) 0:PEGB0, pass, 
			10'd17 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 32, 35 -> 35
			// srcs: (81, 17)(1846) 0, (1847) 0 --> (2626) 0:PEGB0, ALU, +, NI0
			10'd18 : rdata = 48'b000011110000000000111111111100000000000000000000;
			// PEs: 35 -> 32
			// srcs: (120, 21)(1729) -3 --> (1729) -3:NI1, pass, PEGB0
			10'd19 : rdata = 48'b110001010000000100000000000000000000000010000000;
			// PEs: 34, 39 -> 35
			// srcs: (144, 24)(2870) -4, (2872) 2 --> (2873) -2:PENB, PEGB7, +, NI1
			10'd20 : rdata = 48'b000011101111111011100001110100001000000000000000;
			// PEs: 35 -> 32
			// srcs: (149, 22)(2626) 0 --> (2626) 0:NI0, pass, PEGB0
			10'd21 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 32 -> 
			// srcs: (235, 18)(1770) 0 --> (1770) 0:PEGB0, pass, 
			10'd22 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 32, 35 -> 36
			// srcs: (244, 19)(1769) -2, (1770) 0 --> (2552) -2:PEGB0, ALU, +, PENB
			10'd23 : rdata = 48'b000011110000000000111111111000000000000100000000;
			// PEs: 35 -> 32
			// srcs: (350, 23)(2277) 0 --> (2277) 0:NI2, pass, PEGB0
			10'd24 : rdata = 48'b110001010000001000000000000000000000000010000000;
			// PEs: 35 -> 32
			// srcs: (627, 27)(2873) -2 --> (2873) -2:NI1, pass, PEGB0
			10'd25 : rdata = 48'b110001010000000100000000000000000000000010000000;
			// PEs: 32 -> 
			// srcs: (1117, 25)(2861) 3 --> (2861) 3:PEGB0, pass, 
			10'd26 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 35, 38 -> 32
			// srcs: (1119, 26)(2861) 3, (2866) -1 --> (2867) 2:ALU, PEGB6, +, PEGB0
			10'd27 : rdata = 48'b000010011111111111100001100000000000000010000000;
			// PEs: 32, 35 -> 36
			// srcs: (1557, 28)(3140) 47, (47) 2 --> (3184) 94:PEGB0, ND0, *, PENB
			10'd28 : rdata = 48'b000111110000000001100000000000000000000100000000;
			// PEs: 35, 34 -> 34
			// srcs: (1558, 42)(3) 1, (3182) -94 --> (3966) -94:NM0, PENB, *, PEGB2
			10'd29 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 35, 36 -> 35
			// srcs: (1566, 56)(832) 0, (3968) 94 --> (4752) -94:NW0, PEGB4, -, NW0
			10'd30 : rdata = 48'b000100100000000011100001000000000100000000000000;
			// PEs: 32, 35 -> 36
			// srcs: (1637, 29)(3140) 47, (127) -1 --> (3264) -47:PEGB0, ND1, *, PENB
			10'd31 : rdata = 48'b000111110000000001100000001000000000000100000000;
			// PEs: 35, 34 -> 34
			// srcs: (1638, 43)(3) 1, (3262) -141 --> (4046) -141:NM0, PENB, *, PEGB2
			10'd32 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 35, 36 -> 35
			// srcs: (1646, 57)(912) -2, (4048) -47 --> (4832) 45:NW1, PEGB4, -, NW1
			10'd33 : rdata = 48'b000100100000000111100001000000000100010000000000;
			// PEs: 32, 35 -> 
			// srcs: (1670, 30)(3140) 47, (160) 1 --> (3297) 47:PEGB0, ND10, *, 
			10'd34 : rdata = 48'b000111110000000001100001010000000000000000000000;
			// PEs: 35, 35 -> 
			// srcs: (1673, 44)(3) 1, (3297) 47 --> (4081) 47:NM0, ALU, *, 
			10'd35 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 35, 35 -> 35
			// srcs: (1676, 58)(945) -3, (4081) 47 --> (4865) -50:NW10, ALU, -, NW10
			10'd36 : rdata = 48'b000100100000101000111111111000000110100000000000;
			// PEs: 32, 35 -> 36
			// srcs: (1717, 31)(3140) 47, (207) -3 --> (3344) -141:PEGB0, ND2, *, PENB
			10'd37 : rdata = 48'b000111110000000001100000010000000000000100000000;
			// PEs: 35, 34 -> 34
			// srcs: (1718, 45)(3) 1, (3342) -47 --> (4126) -47:NM0, PENB, *, PEGB2
			10'd38 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 35, 36 -> 35
			// srcs: (1726, 59)(992) -3, (4128) -141 --> (4912) 138:NW2, PEGB4, -, NW2
			10'd39 : rdata = 48'b000100100000001011100001000000000100100000000000;
			// PEs: 32, 35 -> 36
			// srcs: (1799, 32)(3140) 47, (289) -2 --> (3426) -94:PEGB0, ND3, *, PENB
			10'd40 : rdata = 48'b000111110000000001100000011000000000000100000000;
			// PEs: 35, 34 -> 34
			// srcs: (1800, 46)(3) 1, (3424) 0 --> (4208) 0:NM0, PENB, *, PEGB2
			10'd41 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 35, 36 -> 35
			// srcs: (1808, 60)(1074) -1, (4210) -94 --> (4994) 93:NW3, PEGB4, -, NW3
			10'd42 : rdata = 48'b000100100000001111100001000000000100110000000000;
			// PEs: 32, 35 -> 
			// srcs: (1850, 33)(3140) 47, (340) -2 --> (3477) -94:PEGB0, ND11, *, 
			10'd43 : rdata = 48'b000111110000000001100001011000000000000000000000;
			// PEs: 35, 35 -> 
			// srcs: (1853, 47)(3) 1, (3477) -94 --> (4261) -94:NM0, ALU, *, 
			10'd44 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 35, 35 -> 35
			// srcs: (1856, 61)(1125) 2, (4261) -94 --> (5045) 96:NW11, ALU, -, NW11
			10'd45 : rdata = 48'b000100100000101100111111111000000110110000000000;
			// PEs: 32, 35 -> 36
			// srcs: (1879, 34)(3140) 47, (369) -1 --> (3506) -47:PEGB0, ND4, *, PENB
			10'd46 : rdata = 48'b000111110000000001100000100000000000000100000000;
			// PEs: 35, 34 -> 34
			// srcs: (1880, 48)(3) 1, (3504) 47 --> (4288) 47:NM0, PENB, *, PEGB2
			10'd47 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 35, 36 -> 35
			// srcs: (1888, 62)(1154) 2, (4290) -47 --> (5074) 49:NW4, PEGB4, -, NW4
			10'd48 : rdata = 48'b000100100000010011100001000000000101000000000000;
			// PEs: 32, 35 -> 36
			// srcs: (1959, 35)(3140) 47, (449) -1 --> (3586) -47:PEGB0, ND5, *, PENB
			10'd49 : rdata = 48'b000111110000000001100000101000000000000100000000;
			// PEs: 35, 34 -> 34
			// srcs: (1961, 49)(3) 1, (3585) 0 --> (4369) 0:NM0, PENB, *, PEGB2
			10'd50 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 35, 36 -> 35
			// srcs: (1968, 63)(1234) 2, (4370) -47 --> (5154) 49:NW5, PEGB4, -, NW5
			10'd51 : rdata = 48'b000100100000010111100001000000000101010000000000;
			// PEs: 32, 35 -> 
			// srcs: (2034, 36)(3140) 47, (524) 2 --> (3661) 94:PEGB0, ND12, *, 
			10'd52 : rdata = 48'b000111110000000001100001100000000000000000000000;
			// PEs: 35, 35 -> 
			// srcs: (2037, 50)(3) 1, (3661) 94 --> (4445) 94:NM0, ALU, *, 
			10'd53 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 35, 35 -> 35
			// srcs: (2040, 64)(1309) 1, (4445) 94 --> (5229) -93:NW12, ALU, -, NW12
			10'd54 : rdata = 48'b000100100000110000111111111000000111000000000000;
			// PEs: 32, 35 -> 36
			// srcs: (2041, 37)(3140) 47, (531) -3 --> (3668) -141:PEGB0, ND6, *, PENB
			10'd55 : rdata = 48'b000111110000000001100000110000000000000100000000;
			// PEs: 35, 34 -> 34
			// srcs: (2042, 51)(3) 1, (3666) 0 --> (4450) 0:NM0, PENB, *, PEGB2
			10'd56 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 35, 36 -> 35
			// srcs: (2050, 65)(1316) 1, (4452) -141 --> (5236) 142:NW6, PEGB4, -, NW6
			10'd57 : rdata = 48'b000100100000011011100001000000000101100000000000;
			// PEs: 32, 35 -> 36
			// srcs: (2121, 38)(3140) 47, (611) 1 --> (3748) 47:PEGB0, ND7, *, PENB
			10'd58 : rdata = 48'b000111110000000001100000111000000000000100000000;
			// PEs: 35, 34 -> 34
			// srcs: (2122, 52)(3) 1, (3746) -47 --> (4530) -47:NM0, PENB, *, PEGB2
			10'd59 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 35, 36 -> 35
			// srcs: (2130, 66)(1396) 0, (4532) 47 --> (5316) -47:NW7, PEGB4, -, NW7
			10'd60 : rdata = 48'b000100100000011111100001000000000101110000000000;
			// PEs: 32, 35 -> 36
			// srcs: (2202, 39)(3140) 47, (692) 2 --> (3829) 94:PEGB0, ND8, *, PENB
			10'd61 : rdata = 48'b000111110000000001100001000000000000000100000000;
			// PEs: 35, 34 -> 34
			// srcs: (2204, 53)(3) 1, (3828) 47 --> (4612) 47:NM0, PENB, *, PEGB2
			10'd62 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 35, 36 -> 35
			// srcs: (2211, 67)(1477) -3, (4613) 94 --> (5397) -97:NW8, PEGB4, -, NW8
			10'd63 : rdata = 48'b000100100000100011100001000000000110000000000000;
			// PEs: 32, 35 -> 
			// srcs: (2218, 40)(3140) 47, (708) 0 --> (3845) 0:PEGB0, ND13, *, 
			10'd64 : rdata = 48'b000111110000000001100001101000000000000000000000;
			// PEs: 35, 35 -> 
			// srcs: (2221, 54)(3) 1, (3845) 0 --> (4629) 0:NM0, ALU, *, 
			10'd65 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 35, 35 -> 35
			// srcs: (2224, 68)(1493) -2, (4629) 0 --> (5413) -2:NW13, ALU, -, NW13
			10'd66 : rdata = 48'b000100100000110100111111111000000111010000000000;
			// PEs: 32, 35 -> 36
			// srcs: (2283, 41)(3140) 47, (773) -2 --> (3910) -94:PEGB0, ND9, *, PENB
			10'd67 : rdata = 48'b000111110000000001100001001000000000000100000000;
			// PEs: 35, 34 -> 34
			// srcs: (2284, 55)(3) 1, (3908) 47 --> (4692) 47:NM0, PENB, *, PEGB2
			10'd68 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 35, 36 -> 35
			// srcs: (2292, 69)(1558) 2, (4694) -94 --> (5478) 96:NW9, PEGB4, -, NW9
			10'd69 : rdata = 48'b000100100000100111100001000000000110010000000000;
			default : rdata = 48'b000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 36) begin
	always @(*) begin
		case(address)
			// PEs: 36, 36 -> 32
			// srcs: (1, 0)(48) -2, (833) 2 --> (1617) -4:ND0, NW0, *, PEGB0
			10'd0 : rdata = 48'b000110110000000001000000000000000000000010000000;
			// PEs: 36, 36 -> 32
			// srcs: (2, 1)(128) -2, (913) -1 --> (1697) 2:ND1, NW1, *, PEGB0
			10'd1 : rdata = 48'b000110110000000101000000001000000000000010000000;
			// PEs: 36, 36 -> 32
			// srcs: (3, 2)(208) -2, (993) -1 --> (1777) 2:ND2, NW2, *, PEGB0
			10'd2 : rdata = 48'b000110110000001001000000010000000000000010000000;
			// PEs: 36, 36 -> 32
			// srcs: (4, 3)(290) 2, (1075) -2 --> (1859) -4:ND3, NW3, *, PEGB0
			10'd3 : rdata = 48'b000110110000001101000000011000000000000010000000;
			// PEs: 36, 36 -> 32
			// srcs: (5, 4)(370) 1, (1155) -1 --> (1939) -1:ND4, NW4, *, PEGB0
			10'd4 : rdata = 48'b000110110000010001000000100000000000000010000000;
			// PEs: 36, 36 -> 32
			// srcs: (6, 5)(450) 0, (1235) 2 --> (2019) 0:ND5, NW5, *, PEGB0
			10'd5 : rdata = 48'b000110110000010101000000101000000000000010000000;
			// PEs: 36, 36 -> 32
			// srcs: (7, 6)(532) -3, (1317) -2 --> (2101) 6:ND6, NW6, *, PEGB0
			10'd6 : rdata = 48'b000110110000011001000000110000000000000010000000;
			// PEs: 36, 36 -> 32
			// srcs: (8, 7)(612) -2, (1397) -1 --> (2181) 2:ND7, NW7, *, PEGB0
			10'd7 : rdata = 48'b000110110000011101000000111000000000000010000000;
			// PEs: 36, 36 -> 35
			// srcs: (9, 8)(693) 1, (1478) 1 --> (2262) 1:ND8, NW8, *, PEGB3
			10'd8 : rdata = 48'b000110110000100001000001000000000000000010110000;
			// PEs: 36, 36 -> 39
			// srcs: (10, 9)(774) -2, (1559) 0 --> (2343) 0:ND9, NW9, *, PEGB7
			10'd9 : rdata = 48'b000110110000100101000001001000000000000011110000;
			// PEs: 36, 36 -> 36
			// srcs: (11, 10)(163) -3, (948) 0 --> (1732) 0:ND10, NW10, *, NI0
			10'd10 : rdata = 48'b000110110000101001000001010100000000000000000000;
			// PEs: 36, 36 -> 36
			// srcs: (12, 11)(343) -3, (1128) -1 --> (1912) 3:ND11, NW11, *, NI1
			10'd11 : rdata = 48'b000110110000101101000001011100001000000000000000;
			// PEs: 36, 36 -> 37
			// srcs: (13, 12)(527) 2, (1312) 2 --> (2096) 4:ND12, NW12, *, PENB
			10'd12 : rdata = 48'b000110110000110001000001100000000000000100000000;
			// PEs: 36, 36 -> 36
			// srcs: (14, 13)(711) 0, (1496) 2 --> (2280) 0:ND13, NW13, *, NI2
			10'd13 : rdata = 48'b000110110000110101000001101100010000000000000000;
			// PEs: 32 -> 
			// srcs: (45, 14)(1688) -3 --> (1688) -3:PEGB0, pass, 
			10'd14 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 32, 36 -> 32
			// srcs: (54, 15)(1687) -2, (1688) -3 --> (2468) -5:PEGB0, ALU, +, PEGB0
			10'd15 : rdata = 48'b000011110000000000111111111000000000000010000000;
			// PEs: 32 -> 
			// srcs: (74, 16)(1850) 3 --> (1850) 3:PEGB0, pass, 
			10'd16 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 32, 36 -> 32
			// srcs: (83, 17)(1849) 0, (1850) 3 --> (2629) 3:PEGB0, ALU, +, PEGB0
			10'd17 : rdata = 48'b000011110000000000111111111000000000000010000000;
			// PEs: 36 -> 32
			// srcs: (120, 20)(1732) 0 --> (1732) 0:NI0, pass, PEGB0
			10'd18 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 36 -> 32
			// srcs: (141, 22)(1912) 3 --> (1912) 3:NI1, pass, PEGB0
			10'd19 : rdata = 48'b110001010000000100000000000000000000000010000000;
			// PEs: 36 -> 32
			// srcs: (163, 23)(2280) 0 --> (2280) 0:NI2, pass, PEGB0
			10'd20 : rdata = 48'b110001010000001000000000000000000000000010000000;
			// PEs: 32 -> 
			// srcs: (266, 18)(1772) 0 --> (1772) 0:PEGB0, pass, 
			10'd21 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 32, 36 -> 
			// srcs: (275, 19)(1771) 1, (1772) 0 --> (2553) 1:PEGB0, ALU, +, 
			10'd22 : rdata = 48'b000011110000000000111111111000000000000000000000;
			// PEs: 35, 36 -> 32
			// srcs: (278, 21)(2552) -2, (2553) 1 --> (2554) -1:PENB, ALU, +, PEGB0
			10'd23 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 32 -> 
			// srcs: (1102, 24)(2945) 11 --> (2945) 11:PEGB0, pass, 
			10'd24 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 36, 33 -> 32
			// srcs: (1104, 25)(2945) 11, (2947) -1 --> (2948) 10:ALU, PEGB1, +, PEGB0
			10'd25 : rdata = 48'b000010011111111111100000010000000000000010000000;
			// PEs: 32, 36 -> 36
			// srcs: (1558, 26)(3140) 47, (48) -2 --> (3185) -94:PEGB0, ND0, *, NI0
			10'd26 : rdata = 48'b000111110000000001100000000100000000000000000000;
			// PEs: 36, 35 -> 35
			// srcs: (1560, 40)(3) 1, (3184) 94 --> (3968) 94:NM0, PENB, *, PEGB3
			10'd27 : rdata = 48'b000111000000000011011111110000000000000010110000;
			// PEs: 36, 36 -> 
			// srcs: (1561, 41)(3) 1, (3185) -94 --> (3969) -94:NM0, NI0, *, 
			10'd28 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 36, 36 -> 36
			// srcs: (1564, 56)(833) 2, (3969) -94 --> (4753) 96:NW0, ALU, -, NW0
			10'd29 : rdata = 48'b000100100000000000111111111000000100000000000000;
			// PEs: 32, 36 -> 37
			// srcs: (1638, 27)(3140) 47, (128) -2 --> (3265) -94:PEGB0, ND1, *, PENB
			10'd30 : rdata = 48'b000111110000000001100000001000000000000100000000;
			// PEs: 36, 35 -> 35
			// srcs: (1640, 42)(3) 1, (3264) -47 --> (4048) -47:NM0, PENB, *, PEGB3
			10'd31 : rdata = 48'b000111000000000011011111110000000000000010110000;
			// PEs: 36, 37 -> 36
			// srcs: (1647, 57)(913) -1, (4049) -94 --> (4833) 93:NW1, PEGB5, -, NW1
			10'd32 : rdata = 48'b000100100000000111100001010000000100010000000000;
			// PEs: 32, 36 -> 
			// srcs: (1673, 28)(3140) 47, (163) -3 --> (3300) -141:PEGB0, ND10, *, 
			10'd33 : rdata = 48'b000111110000000001100001010000000000000000000000;
			// PEs: 36, 36 -> 
			// srcs: (1676, 43)(3) 1, (3300) -141 --> (4084) -141:NM0, ALU, *, 
			10'd34 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 36, 36 -> 36
			// srcs: (1679, 58)(948) 0, (4084) -141 --> (4868) 141:NW10, ALU, -, NW10
			10'd35 : rdata = 48'b000100100000101000111111111000000110100000000000;
			// PEs: 32, 36 -> 37
			// srcs: (1718, 29)(3140) 47, (208) -2 --> (3345) -94:PEGB0, ND2, *, PENB
			10'd36 : rdata = 48'b000111110000000001100000010000000000000100000000;
			// PEs: 36, 35 -> 35
			// srcs: (1720, 44)(3) 1, (3344) -141 --> (4128) -141:NM0, PENB, *, PEGB3
			10'd37 : rdata = 48'b000111000000000011011111110000000000000010110000;
			// PEs: 36, 37 -> 36
			// srcs: (1727, 59)(993) -1, (4129) -94 --> (4913) 93:NW2, PEGB5, -, NW2
			10'd38 : rdata = 48'b000100100000001011100001010000000100100000000000;
			// PEs: 32, 36 -> 37
			// srcs: (1800, 30)(3140) 47, (290) 2 --> (3427) 94:PEGB0, ND3, *, PENB
			10'd39 : rdata = 48'b000111110000000001100000011000000000000100000000;
			// PEs: 36, 35 -> 35
			// srcs: (1802, 45)(3) 1, (3426) -94 --> (4210) -94:NM0, PENB, *, PEGB3
			10'd40 : rdata = 48'b000111000000000011011111110000000000000010110000;
			// PEs: 36, 37 -> 36
			// srcs: (1809, 60)(1075) -2, (4211) 94 --> (4995) -96:NW3, PEGB5, -, NW3
			10'd41 : rdata = 48'b000100100000001111100001010000000100110000000000;
			// PEs: 32, 36 -> 
			// srcs: (1853, 31)(3140) 47, (343) -3 --> (3480) -141:PEGB0, ND11, *, 
			10'd42 : rdata = 48'b000111110000000001100001011000000000000000000000;
			// PEs: 36, 36 -> 
			// srcs: (1856, 46)(3) 1, (3480) -141 --> (4264) -141:NM0, ALU, *, 
			10'd43 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 36, 36 -> 36
			// srcs: (1859, 61)(1128) -1, (4264) -141 --> (5048) 140:NW11, ALU, -, NW11
			10'd44 : rdata = 48'b000100100000101100111111111000000110110000000000;
			// PEs: 32, 36 -> 37
			// srcs: (1880, 32)(3140) 47, (370) 1 --> (3507) 47:PEGB0, ND4, *, PENB
			10'd45 : rdata = 48'b000111110000000001100000100000000000000100000000;
			// PEs: 36, 35 -> 35
			// srcs: (1882, 47)(3) 1, (3506) -47 --> (4290) -47:NM0, PENB, *, PEGB3
			10'd46 : rdata = 48'b000111000000000011011111110000000000000010110000;
			// PEs: 36, 37 -> 36
			// srcs: (1889, 62)(1155) -1, (4291) 47 --> (5075) -48:NW4, PEGB5, -, NW4
			10'd47 : rdata = 48'b000100100000010011100001010000000101000000000000;
			// PEs: 32, 36 -> 37
			// srcs: (1960, 33)(3140) 47, (450) 0 --> (3587) 0:PEGB0, ND5, *, PENB
			10'd48 : rdata = 48'b000111110000000001100000101000000000000100000000;
			// PEs: 36, 35 -> 35
			// srcs: (1962, 48)(3) 1, (3586) -47 --> (4370) -47:NM0, PENB, *, PEGB3
			10'd49 : rdata = 48'b000111000000000011011111110000000000000010110000;
			// PEs: 36, 37 -> 36
			// srcs: (1969, 63)(1235) 2, (4371) 0 --> (5155) 2:NW5, PEGB5, -, NW5
			10'd50 : rdata = 48'b000100100000010111100001010000000101010000000000;
			// PEs: 32, 36 -> 
			// srcs: (2037, 34)(3140) 47, (527) 2 --> (3664) 94:PEGB0, ND12, *, 
			10'd51 : rdata = 48'b000111110000000001100001100000000000000000000000;
			// PEs: 36, 36 -> 36
			// srcs: (2040, 49)(3) 1, (3664) 94 --> (4448) 94:NM0, ALU, *, NI0
			10'd52 : rdata = 48'b000111000000000000111111111100000000000000000000;
			// PEs: 32, 36 -> 37
			// srcs: (2042, 35)(3140) 47, (532) -3 --> (3669) -141:PEGB0, ND6, *, PENB
			10'd53 : rdata = 48'b000111110000000001100000110000000000000100000000;
			// PEs: 36, 36 -> 36
			// srcs: (2043, 64)(1312) 2, (4448) 94 --> (5232) -92:NW12, NI0, -, NW12
			10'd54 : rdata = 48'b000100100000110010100000000000000111000000000000;
			// PEs: 36, 35 -> 35
			// srcs: (2044, 50)(3) 1, (3668) -141 --> (4452) -141:NM0, PENB, *, PEGB3
			10'd55 : rdata = 48'b000111000000000011011111110000000000000010110000;
			// PEs: 36, 37 -> 36
			// srcs: (2051, 65)(1317) -2, (4453) -141 --> (5237) 139:NW6, PEGB5, -, NW6
			10'd56 : rdata = 48'b000100100000011011100001010000000101100000000000;
			// PEs: 32, 36 -> 37
			// srcs: (2122, 36)(3140) 47, (612) -2 --> (3749) -94:PEGB0, ND7, *, PENB
			10'd57 : rdata = 48'b000111110000000001100000111000000000000100000000;
			// PEs: 36, 35 -> 35
			// srcs: (2124, 51)(3) 1, (3748) 47 --> (4532) 47:NM0, PENB, *, PEGB3
			10'd58 : rdata = 48'b000111000000000011011111110000000000000010110000;
			// PEs: 36, 37 -> 36
			// srcs: (2131, 66)(1397) -1, (4533) -94 --> (5317) 93:NW7, PEGB5, -, NW7
			10'd59 : rdata = 48'b000100100000011111100001010000000101110000000000;
			// PEs: 32, 36 -> 37
			// srcs: (2203, 37)(3140) 47, (693) 1 --> (3830) 47:PEGB0, ND8, *, PENB
			10'd60 : rdata = 48'b000111110000000001100001000000000000000100000000;
			// PEs: 36, 35 -> 35
			// srcs: (2205, 52)(3) 1, (3829) 94 --> (4613) 94:NM0, PENB, *, PEGB3
			10'd61 : rdata = 48'b000111000000000011011111110000000000000010110000;
			// PEs: 36, 37 -> 36
			// srcs: (2212, 67)(1478) 1, (4614) 47 --> (5398) -46:NW8, PEGB5, -, NW8
			10'd62 : rdata = 48'b000100100000100011100001010000000110000000000000;
			// PEs: 32, 36 -> 
			// srcs: (2221, 38)(3140) 47, (711) 0 --> (3848) 0:PEGB0, ND13, *, 
			10'd63 : rdata = 48'b000111110000000001100001101000000000000000000000;
			// PEs: 36, 36 -> 
			// srcs: (2224, 53)(3) 1, (3848) 0 --> (4632) 0:NM0, ALU, *, 
			10'd64 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 36, 36 -> 36
			// srcs: (2227, 68)(1496) 2, (4632) 0 --> (5416) 2:NW13, ALU, -, NW13
			10'd65 : rdata = 48'b000100100000110100111111111000000111010000000000;
			// PEs: 32, 36 -> 36
			// srcs: (2284, 39)(3140) 47, (774) -2 --> (3911) -94:PEGB0, ND9, *, NI0
			10'd66 : rdata = 48'b000111110000000001100001001100000000000000000000;
			// PEs: 36, 35 -> 35
			// srcs: (2286, 54)(3) 1, (3910) -94 --> (4694) -94:NM0, PENB, *, PEGB3
			10'd67 : rdata = 48'b000111000000000011011111110000000000000010110000;
			// PEs: 36, 36 -> 
			// srcs: (2287, 55)(3) 1, (3911) -94 --> (4695) -94:NM0, NI0, *, 
			10'd68 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 36, 36 -> 36
			// srcs: (2290, 69)(1559) 0, (4695) -94 --> (5479) 94:NW9, ALU, -, NW9
			10'd69 : rdata = 48'b000100100000100100111111111000000110010000000000;
			default : rdata = 48'b000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 37) begin
	always @(*) begin
		case(address)
			// PEs: 37, 37 -> 32
			// srcs: (1, 0)(50) -2, (835) 0 --> (1619) 0:ND0, NW0, *, PEGB0
			10'd0 : rdata = 48'b000110110000000001000000000000000000000010000000;
			// PEs: 37, 37 -> 32
			// srcs: (2, 1)(130) 1, (915) 0 --> (1699) 0:ND1, NW1, *, PEGB0
			10'd1 : rdata = 48'b000110110000000101000000001000000000000010000000;
			// PEs: 37, 37 -> 32
			// srcs: (3, 2)(210) 1, (995) 0 --> (1779) 0:ND2, NW2, *, PEGB0
			10'd2 : rdata = 48'b000110110000001001000000010000000000000010000000;
			// PEs: 37, 37 -> 32
			// srcs: (4, 3)(292) -1, (1077) -1 --> (1861) 1:ND3, NW3, *, PEGB0
			10'd3 : rdata = 48'b000110110000001101000000011000000000000010000000;
			// PEs: 37, 37 -> 32
			// srcs: (5, 4)(372) 0, (1157) -3 --> (1941) 0:ND4, NW4, *, PEGB0
			10'd4 : rdata = 48'b000110110000010001000000100000000000000010000000;
			// PEs: 37, 37 -> 32
			// srcs: (6, 5)(452) -2, (1237) -1 --> (2021) 2:ND5, NW5, *, PEGB0
			10'd5 : rdata = 48'b000110110000010101000000101000000000000010000000;
			// PEs: 37, 37 -> 32
			// srcs: (7, 6)(534) 1, (1319) 0 --> (2103) 0:ND6, NW6, *, PEGB0
			10'd6 : rdata = 48'b000110110000011001000000110000000000000010000000;
			// PEs: 37, 37 -> 32
			// srcs: (8, 7)(614) -1, (1399) 2 --> (2183) -2:ND7, NW7, *, PEGB0
			10'd7 : rdata = 48'b000110110000011101000000111000000000000010000000;
			// PEs: 37, 37 -> 39
			// srcs: (9, 8)(694) 2, (1479) -2 --> (2263) -4:ND8, NW8, *, PEGB7
			10'd8 : rdata = 48'b000110110000100001000001000000000000000011110000;
			// PEs: 37, 37 -> 34
			// srcs: (10, 9)(776) -3, (1561) -2 --> (2345) 6:ND9, NW9, *, PEGB2
			10'd9 : rdata = 48'b000110110000100101000001001000000000000010100000;
			// PEs: 37, 37 -> 33
			// srcs: (11, 10)(166) 2, (951) -1 --> (1735) -2:ND10, NW10, *, PEGB1
			10'd10 : rdata = 48'b000110110000101001000001010000000000000010010000;
			// PEs: 37, 37 -> 37
			// srcs: (12, 11)(346) -2, (1131) 0 --> (1915) 0:ND11, NW11, *, NI0
			10'd11 : rdata = 48'b000110110000101101000001011100000000000000000000;
			// PEs: 37, 37 -> 37
			// srcs: (13, 12)(530) 1, (1315) 0 --> (2099) 0:ND12, NW12, *, NI1
			10'd12 : rdata = 48'b000110110000110001000001100100001000000000000000;
			// PEs: 37, 37 -> 37
			// srcs: (14, 13)(714) -3, (1499) 2 --> (2283) -6:ND13, NW13, *, NI2
			10'd13 : rdata = 48'b000110110000110101000001101100010000000000000000;
			// PEs: 34 -> 
			// srcs: (15, 18)(2260) -1 --> (2260) -1:PEGB2, pass, 
			10'd14 : rdata = 48'b110001110000010000000000000000000000000000000000;
			// PEs: 33, 37 -> 38
			// srcs: (17, 19)(2259) 0, (2260) -1 --> (3040) -1:PEGB1, ALU, +, PENB
			10'd15 : rdata = 48'b000011110000001000111111111000000000000100000000;
			// PEs: 32 -> 
			// srcs: (47, 14)(1691) 6 --> (1691) 6:PEGB0, pass, 
			10'd16 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 32, 37 -> 32
			// srcs: (56, 15)(1690) 9, (1691) 6 --> (2471) 15:PEGB0, ALU, +, PEGB0
			10'd17 : rdata = 48'b000011110000000000111111111000000000000010000000;
			// PEs: 32 -> 
			// srcs: (76, 16)(1853) -2 --> (1853) -2:PEGB0, pass, 
			10'd18 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 32, 37 -> 33
			// srcs: (85, 17)(1852) 2, (1853) -2 --> (2631) 0:PEGB0, ALU, +, PEGB1
			10'd19 : rdata = 48'b000011110000000000111111111000000000000010010000;
			// PEs: 37 -> 32
			// srcs: (141, 20)(1915) 0 --> (1915) 0:NI0, pass, PEGB0
			10'd20 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 33, 36 -> 37
			// srcs: (144, 21)(2874) 4, (2096) 4 --> (2875) 8:PEGB1, PENB, +, NI0
			10'd21 : rdata = 48'b000011110000001011011111110100000000000000000000;
			// PEs: 37 -> 32
			// srcs: (151, 23)(2283) -6 --> (2283) -6:NI2, pass, PEGB0
			10'd22 : rdata = 48'b110001010000001000000000000000000000000010000000;
			// PEs: 37 -> 32
			// srcs: (307, 22)(2099) 0 --> (2099) 0:NI1, pass, PEGB0
			10'd23 : rdata = 48'b110001010000000100000000000000000000000010000000;
			// PEs: 37 -> 32
			// srcs: (382, 24)(2875) 8 --> (2875) 8:NI0, pass, PEGB0
			10'd24 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 32 -> 
			// srcs: (1119, 25)(3132) 7 --> (3132) 7:PEGB0, pass, 
			10'd25 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 33, 37 -> 32
			// srcs: (1121, 26)(3127) 4, (3132) 7 --> (3133) 11:PEGB1, ALU, +, PEGB0
			10'd26 : rdata = 48'b000011110000001000111111111000000000000010000000;
			// PEs: 32, 37 -> 38
			// srcs: (1560, 27)(3140) 47, (50) -2 --> (3187) -94:PEGB0, ND0, *, PENB
			10'd27 : rdata = 48'b000111110000000001100000000000000000000100000000;
			// PEs: 37, 38 -> 37
			// srcs: (1569, 56)(835) 0, (3971) -94 --> (4755) 94:NW0, PEGB6, -, NW0
			10'd28 : rdata = 48'b000100100000000011100001100000000100000000000000;
			// PEs: 32, 37 -> 38
			// srcs: (1640, 28)(3140) 47, (130) 1 --> (3267) 47:PEGB0, ND1, *, PENB
			10'd29 : rdata = 48'b000111110000000001100000001000000000000100000000;
			// PEs: 37, 36 -> 36
			// srcs: (1641, 41)(3) 1, (3265) -94 --> (4049) -94:NM0, PENB, *, PEGB4
			10'd30 : rdata = 48'b000111000000000011011111110000000000000011000000;
			// PEs: 37, 38 -> 37
			// srcs: (1649, 57)(915) 0, (4051) 47 --> (4835) -47:NW1, PEGB6, -, NW1
			10'd31 : rdata = 48'b000100100000000111100001100000000100010000000000;
			// PEs: 32, 37 -> 
			// srcs: (1676, 29)(3140) 47, (166) 2 --> (3303) 94:PEGB0, ND10, *, 
			10'd32 : rdata = 48'b000111110000000001100001010000000000000000000000;
			// PEs: 37, 37 -> 
			// srcs: (1679, 42)(3) 1, (3303) 94 --> (4087) 94:NM0, ALU, *, 
			10'd33 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 37, 37 -> 37
			// srcs: (1682, 58)(951) -1, (4087) 94 --> (4871) -95:NW10, ALU, -, NW10
			10'd34 : rdata = 48'b000100100000101000111111111000000110100000000000;
			// PEs: 32, 37 -> 38
			// srcs: (1720, 30)(3140) 47, (210) 1 --> (3347) 47:PEGB0, ND2, *, PENB
			10'd35 : rdata = 48'b000111110000000001100000010000000000000100000000;
			// PEs: 37, 36 -> 36
			// srcs: (1721, 43)(3) 1, (3345) -94 --> (4129) -94:NM0, PENB, *, PEGB4
			10'd36 : rdata = 48'b000111000000000011011111110000000000000011000000;
			// PEs: 37, 38 -> 37
			// srcs: (1729, 59)(995) 0, (4131) 47 --> (4915) -47:NW2, PEGB6, -, NW2
			10'd37 : rdata = 48'b000100100000001011100001100000000100100000000000;
			// PEs: 32, 37 -> 38
			// srcs: (1802, 31)(3140) 47, (292) -1 --> (3429) -47:PEGB0, ND3, *, PENB
			10'd38 : rdata = 48'b000111110000000001100000011000000000000100000000;
			// PEs: 37, 36 -> 36
			// srcs: (1803, 44)(3) 1, (3427) 94 --> (4211) 94:NM0, PENB, *, PEGB4
			10'd39 : rdata = 48'b000111000000000011011111110000000000000011000000;
			// PEs: 37, 38 -> 37
			// srcs: (1811, 60)(1077) -1, (4213) -47 --> (4997) 46:NW3, PEGB6, -, NW3
			10'd40 : rdata = 48'b000100100000001111100001100000000100110000000000;
			// PEs: 32, 37 -> 
			// srcs: (1856, 32)(3140) 47, (346) -2 --> (3483) -94:PEGB0, ND11, *, 
			10'd41 : rdata = 48'b000111110000000001100001011000000000000000000000;
			// PEs: 37, 37 -> 
			// srcs: (1859, 45)(3) 1, (3483) -94 --> (4267) -94:NM0, ALU, *, 
			10'd42 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 37, 37 -> 37
			// srcs: (1862, 61)(1131) 0, (4267) -94 --> (5051) 94:NW11, ALU, -, NW11
			10'd43 : rdata = 48'b000100100000101100111111111000000110110000000000;
			// PEs: 32, 37 -> 37
			// srcs: (1882, 33)(3140) 47, (372) 0 --> (3509) 0:PEGB0, ND4, *, NI0
			10'd44 : rdata = 48'b000111110000000001100000100100000000000000000000;
			// PEs: 37, 36 -> 36
			// srcs: (1883, 46)(3) 1, (3507) 47 --> (4291) 47:NM0, PENB, *, PEGB4
			10'd45 : rdata = 48'b000111000000000011011111110000000000000011000000;
			// PEs: 37, 37 -> 
			// srcs: (1885, 47)(3) 1, (3509) 0 --> (4293) 0:NM0, NI0, *, 
			10'd46 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 37, 37 -> 37
			// srcs: (1888, 62)(1157) -3, (4293) 0 --> (5077) -3:NW4, ALU, -, NW4
			10'd47 : rdata = 48'b000100100000010000111111111000000101000000000000;
			// PEs: 32, 37 -> 38
			// srcs: (1962, 34)(3140) 47, (452) -2 --> (3589) -94:PEGB0, ND5, *, PENB
			10'd48 : rdata = 48'b000111110000000001100000101000000000000100000000;
			// PEs: 37, 36 -> 36
			// srcs: (1963, 48)(3) 1, (3587) 0 --> (4371) 0:NM0, PENB, *, PEGB4
			10'd49 : rdata = 48'b000111000000000011011111110000000000000011000000;
			// PEs: 37, 38 -> 37
			// srcs: (1971, 63)(1237) -1, (4373) -94 --> (5157) 93:NW5, PEGB6, -, NW5
			10'd50 : rdata = 48'b000100100000010111100001100000000101010000000000;
			// PEs: 32, 37 -> 
			// srcs: (2040, 35)(3140) 47, (530) 1 --> (3667) 47:PEGB0, ND12, *, 
			10'd51 : rdata = 48'b000111110000000001100001100000000000000000000000;
			// PEs: 37, 37 -> 37
			// srcs: (2043, 49)(3) 1, (3667) 47 --> (4451) 47:NM0, ALU, *, NI0
			10'd52 : rdata = 48'b000111000000000000111111111100000000000000000000;
			// PEs: 32, 37 -> 38
			// srcs: (2044, 36)(3140) 47, (534) 1 --> (3671) 47:PEGB0, ND6, *, PENB
			10'd53 : rdata = 48'b000111110000000001100000110000000000000100000000;
			// PEs: 37, 36 -> 36
			// srcs: (2045, 50)(3) 1, (3669) -141 --> (4453) -141:NM0, PENB, *, PEGB4
			10'd54 : rdata = 48'b000111000000000011011111110000000000000011000000;
			// PEs: 37, 37 -> 37
			// srcs: (2046, 64)(1315) 0, (4451) 47 --> (5235) -47:NW12, NI0, -, NW12
			10'd55 : rdata = 48'b000100100000110010100000000000000111000000000000;
			// PEs: 37, 38 -> 37
			// srcs: (2053, 65)(1319) 0, (4455) 47 --> (5239) -47:NW6, PEGB6, -, NW6
			10'd56 : rdata = 48'b000100100000011011100001100000000101100000000000;
			// PEs: 32, 37 -> 38
			// srcs: (2124, 37)(3140) 47, (614) -1 --> (3751) -47:PEGB0, ND7, *, PENB
			10'd57 : rdata = 48'b000111110000000001100000111000000000000100000000;
			// PEs: 37, 36 -> 36
			// srcs: (2125, 51)(3) 1, (3749) -94 --> (4533) -94:NM0, PENB, *, PEGB4
			10'd58 : rdata = 48'b000111000000000011011111110000000000000011000000;
			// PEs: 37, 38 -> 37
			// srcs: (2133, 66)(1399) 2, (4535) -47 --> (5319) 49:NW7, PEGB6, -, NW7
			10'd59 : rdata = 48'b000100100000011111100001100000000101110000000000;
			// PEs: 32, 37 -> 37
			// srcs: (2204, 38)(3140) 47, (694) 2 --> (3831) 94:PEGB0, ND8, *, NI0
			10'd60 : rdata = 48'b000111110000000001100001000100000000000000000000;
			// PEs: 37, 36 -> 36
			// srcs: (2206, 52)(3) 1, (3830) 47 --> (4614) 47:NM0, PENB, *, PEGB4
			10'd61 : rdata = 48'b000111000000000011011111110000000000000011000000;
			// PEs: 37, 37 -> 
			// srcs: (2207, 53)(3) 1, (3831) 94 --> (4615) 94:NM0, NI0, *, 
			10'd62 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 37, 37 -> 37
			// srcs: (2210, 67)(1479) -2, (4615) 94 --> (5399) -96:NW8, ALU, -, NW8
			10'd63 : rdata = 48'b000100100000100000111111111000000110000000000000;
			// PEs: 32, 37 -> 
			// srcs: (2224, 39)(3140) 47, (714) -3 --> (3851) -141:PEGB0, ND13, *, 
			10'd64 : rdata = 48'b000111110000000001100001101000000000000000000000;
			// PEs: 37, 37 -> 
			// srcs: (2227, 54)(3) 1, (3851) -141 --> (4635) -141:NM0, ALU, *, 
			10'd65 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 37, 37 -> 37
			// srcs: (2230, 68)(1499) 2, (4635) -141 --> (5419) 143:NW13, ALU, -, NW13
			10'd66 : rdata = 48'b000100100000110100111111111000000111010000000000;
			// PEs: 32, 37 -> 
			// srcs: (2286, 40)(3140) 47, (776) -3 --> (3913) -141:PEGB0, ND9, *, 
			10'd67 : rdata = 48'b000111110000000001100001001000000000000000000000;
			// PEs: 37, 37 -> 
			// srcs: (2289, 55)(3) 1, (3913) -141 --> (4697) -141:NM0, ALU, *, 
			10'd68 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 37, 37 -> 37
			// srcs: (2292, 69)(1561) -2, (4697) -141 --> (5481) 139:NW9, ALU, -, NW9
			10'd69 : rdata = 48'b000100100000100100111111111000000110010000000000;
			default : rdata = 48'b000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 38) begin
	always @(*) begin
		case(address)
			// PEs: 38, 38 -> 32
			// srcs: (1, 0)(51) 0, (836) -2 --> (1620) 0:ND0, NW0, *, PEGB0
			10'd0 : rdata = 48'b000110110000000001000000000000000000000010000000;
			// PEs: 38, 38 -> 32
			// srcs: (2, 1)(131) -2, (916) 1 --> (1700) -2:ND1, NW1, *, PEGB0
			10'd1 : rdata = 48'b000110110000000101000000001000000000000010000000;
			// PEs: 38, 38 -> 32
			// srcs: (3, 2)(211) -3, (996) 2 --> (1780) -6:ND2, NW2, *, PEGB0
			10'd2 : rdata = 48'b000110110000001001000000010000000000000010000000;
			// PEs: 38, 38 -> 32
			// srcs: (4, 3)(293) 1, (1078) 0 --> (1862) 0:ND3, NW3, *, PEGB0
			10'd3 : rdata = 48'b000110110000001101000000011000000000000010000000;
			// PEs: 38, 38 -> 32
			// srcs: (5, 4)(373) -1, (1158) -2 --> (1942) 2:ND4, NW4, *, PEGB0
			10'd4 : rdata = 48'b000110110000010001000000100000000000000010000000;
			// PEs: 38, 38 -> 32
			// srcs: (6, 5)(453) 0, (1238) -1 --> (2022) 0:ND5, NW5, *, PEGB0
			10'd5 : rdata = 48'b000110110000010101000000101000000000000010000000;
			// PEs: 38, 38 -> 32
			// srcs: (7, 6)(535) 2, (1320) 0 --> (2104) 0:ND6, NW6, *, PEGB0
			10'd6 : rdata = 48'b000110110000011001000000110000000000000010000000;
			// PEs: 38, 38 -> 32
			// srcs: (8, 7)(615) 1, (1400) -3 --> (2184) -3:ND7, NW7, *, PEGB0
			10'd7 : rdata = 48'b000110110000011101000000111000000000000010000000;
			// PEs: 38, 38 -> 39
			// srcs: (9, 8)(695) 1, (1480) -1 --> (2264) -1:ND8, NW8, *, PENB
			10'd8 : rdata = 48'b000110110000100001000001000000000000000100000000;
			// PEs: 38, 38 -> 34
			// srcs: (10, 9)(777) 1, (1562) 1 --> (2346) 1:ND9, NW9, *, PEGB2
			10'd9 : rdata = 48'b000110110000100101000001001000000000000010100000;
			// PEs: 38, 38 -> 32
			// srcs: (11, 10)(169) -2, (954) 0 --> (1738) 0:ND10, NW10, *, PEGB0
			10'd10 : rdata = 48'b000110110000101001000001010000000000000010000000;
			// PEs: 38, 38 -> 38
			// srcs: (12, 11)(353) -2, (1138) -3 --> (1922) 6:ND11, NW11, *, NI0
			10'd11 : rdata = 48'b000110110000101101000001011100000000000000000000;
			// PEs: 38, 38 -> 32
			// srcs: (13, 12)(533) 0, (1318) -2 --> (2102) 0:ND12, NW12, *, PEGB0
			10'd12 : rdata = 48'b000110110000110001000001100000000000000010000000;
			// PEs: 38, 38 -> 38
			// srcs: (14, 13)(717) 1, (1502) -1 --> (2286) -1:ND13, NW13, *, NI1
			10'd13 : rdata = 48'b000110110000110101000001101100001000000000000000;
			// PEs: 34 -> 
			// srcs: (15, 16)(2340) -2 --> (2340) -2:PEGB2, pass, 
			10'd14 : rdata = 48'b110001110000010000000000000000000000000000000000;
			// PEs: 33, 38 -> 32
			// srcs: (18, 17)(2339) 1, (2340) -2 --> (3117) -1:PEGB1, ALU, +, PEGB0
			10'd15 : rdata = 48'b000011110000001000111111111000000000000010000000;
			// PEs: 37, 35 -> 39
			// srcs: (23, 21)(3040) -1, (3041) -5 --> (3042) -6:PENB, PEGB3, +, PENB
			10'd16 : rdata = 48'b000011101111111011100000110000000000000100000000;
			// PEs: 32 -> 
			// srcs: (55, 14)(1763) 0 --> (1763) 0:PEGB0, pass, 
			10'd17 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 38, 32 -> 33
			// srcs: (64, 15)(1763) 0, (1764) 0 --> (2542) 0:ALU, PEGB0, +, PEGB1
			10'd18 : rdata = 48'b000010011111111111100000000000000000000010010000;
			// PEs: 38 -> 33
			// srcs: (367, 18)(1922) 6 --> (1922) 6:NI0, pass, PEGB1
			10'd19 : rdata = 48'b110001010000000000000000000000000000000010010000;
			// PEs: 32 -> 
			// srcs: (369, 19)(2703) -8 --> (2703) -8:PEGB0, pass, 
			10'd20 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 38, 39 -> 32
			// srcs: (371, 20)(2703) -8, (1925) 2 --> (2704) -6:ALU, PEGB7, +, PEGB0
			10'd21 : rdata = 48'b000010011111111111100001110000000000000010000000;
			// PEs: 38 -> 33
			// srcs: (416, 22)(2286) -1 --> (2286) -1:NI1, pass, PEGB1
			10'd22 : rdata = 48'b110001010000000100000000000000000000000010010000;
			// PEs: 32 -> 
			// srcs: (1101, 23)(2863) 0 --> (2863) 0:PEGB0, pass, 
			10'd23 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 38, 33 -> 35
			// srcs: (1103, 24)(2863) 0, (2865) -1 --> (2866) -1:ALU, PEGB1, +, PEGB3
			10'd24 : rdata = 48'b000010011111111111100000010000000000000010110000;
			// PEs: 32, 38 -> 39
			// srcs: (1561, 25)(3140) 47, (51) 0 --> (3188) 0:PEGB0, ND0, *, PENB
			10'd25 : rdata = 48'b000111110000000001100000000000000000000100000000;
			// PEs: 38, 37 -> 37
			// srcs: (1563, 39)(3) 1, (3187) -94 --> (3971) -94:NM0, PENB, *, PEGB5
			10'd26 : rdata = 48'b000111000000000011011111110000000000000011010000;
			// PEs: 38, 39 -> 38
			// srcs: (1570, 56)(836) -2, (3972) 0 --> (4756) -2:NW0, PEGB7, -, NW0
			10'd27 : rdata = 48'b000100100000000011100001110000000100000000000000;
			// PEs: 32, 38 -> 38
			// srcs: (1641, 26)(3140) 47, (131) -2 --> (3268) -94:PEGB0, ND1, *, NI0
			10'd28 : rdata = 48'b000111110000000001100000001100000000000000000000;
			// PEs: 38, 37 -> 37
			// srcs: (1643, 40)(3) 1, (3267) 47 --> (4051) 47:NM0, PENB, *, PEGB5
			10'd29 : rdata = 48'b000111000000000011011111110000000000000011010000;
			// PEs: 38, 38 -> 
			// srcs: (1644, 41)(3) 1, (3268) -94 --> (4052) -94:NM0, NI0, *, 
			10'd30 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 38, 38 -> 38
			// srcs: (1647, 57)(916) 1, (4052) -94 --> (4836) 95:NW1, ALU, -, NW1
			10'd31 : rdata = 48'b000100100000000100111111111000000100010000000000;
			// PEs: 32, 38 -> 
			// srcs: (1679, 27)(3140) 47, (169) -2 --> (3306) -94:PEGB0, ND10, *, 
			10'd32 : rdata = 48'b000111110000000001100001010000000000000000000000;
			// PEs: 38, 38 -> 
			// srcs: (1682, 42)(3) 1, (3306) -94 --> (4090) -94:NM0, ALU, *, 
			10'd33 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 38, 38 -> 38
			// srcs: (1685, 58)(954) 0, (4090) -94 --> (4874) 94:NW10, ALU, -, NW10
			10'd34 : rdata = 48'b000100100000101000111111111000000110100000000000;
			// PEs: 32, 38 -> 39
			// srcs: (1721, 28)(3140) 47, (211) -3 --> (3348) -141:PEGB0, ND2, *, PENB
			10'd35 : rdata = 48'b000111110000000001100000010000000000000100000000;
			// PEs: 38, 37 -> 37
			// srcs: (1723, 43)(3) 1, (3347) 47 --> (4131) 47:NM0, PENB, *, PEGB5
			10'd36 : rdata = 48'b000111000000000011011111110000000000000011010000;
			// PEs: 38, 39 -> 38
			// srcs: (1730, 59)(996) 2, (4132) -141 --> (4916) 143:NW2, PEGB7, -, NW2
			10'd37 : rdata = 48'b000100100000001011100001110000000100100000000000;
			// PEs: 32, 38 -> 38
			// srcs: (1803, 29)(3140) 47, (293) 1 --> (3430) 47:PEGB0, ND3, *, NI0
			10'd38 : rdata = 48'b000111110000000001100000011100000000000000000000;
			// PEs: 38, 37 -> 37
			// srcs: (1805, 44)(3) 1, (3429) -47 --> (4213) -47:NM0, PENB, *, PEGB5
			10'd39 : rdata = 48'b000111000000000011011111110000000000000011010000;
			// PEs: 38, 38 -> 
			// srcs: (1806, 45)(3) 1, (3430) 47 --> (4214) 47:NM0, NI0, *, 
			10'd40 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 38, 38 -> 38
			// srcs: (1809, 60)(1078) 0, (4214) 47 --> (4998) -47:NW3, ALU, -, NW3
			10'd41 : rdata = 48'b000100100000001100111111111000000100110000000000;
			// PEs: 32, 38 -> 
			// srcs: (1863, 30)(3140) 47, (353) -2 --> (3490) -94:PEGB0, ND11, *, 
			10'd42 : rdata = 48'b000111110000000001100001011000000000000000000000;
			// PEs: 38, 38 -> 
			// srcs: (1866, 46)(3) 1, (3490) -94 --> (4274) -94:NM0, ALU, *, 
			10'd43 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 38, 38 -> 38
			// srcs: (1869, 61)(1138) -3, (4274) -94 --> (5058) 91:NW11, ALU, -, NW11
			10'd44 : rdata = 48'b000100100000101100111111111000000110110000000000;
			// PEs: 32, 38 -> 
			// srcs: (1883, 31)(3140) 47, (373) -1 --> (3510) -47:PEGB0, ND4, *, 
			10'd45 : rdata = 48'b000111110000000001100000100000000000000000000000;
			// PEs: 38, 38 -> 
			// srcs: (1886, 47)(3) 1, (3510) -47 --> (4294) -47:NM0, ALU, *, 
			10'd46 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 38, 38 -> 38
			// srcs: (1889, 62)(1158) -2, (4294) -47 --> (5078) 45:NW4, ALU, -, NW4
			10'd47 : rdata = 48'b000100100000010000111111111000000101000000000000;
			// PEs: 32, 38 -> 39
			// srcs: (1963, 32)(3140) 47, (453) 0 --> (3590) 0:PEGB0, ND5, *, PENB
			10'd48 : rdata = 48'b000111110000000001100000101000000000000100000000;
			// PEs: 38, 37 -> 37
			// srcs: (1965, 48)(3) 1, (3589) -94 --> (4373) -94:NM0, PENB, *, PEGB5
			10'd49 : rdata = 48'b000111000000000011011111110000000000000011010000;
			// PEs: 38, 39 -> 38
			// srcs: (1972, 63)(1238) -1, (4374) 0 --> (5158) -1:NW5, PEGB7, -, NW5
			10'd50 : rdata = 48'b000100100000010111100001110000000101010000000000;
			// PEs: 32, 38 -> 38
			// srcs: (2043, 33)(3140) 47, (533) 0 --> (3670) 0:PEGB0, ND12, *, NI0
			10'd51 : rdata = 48'b000111110000000001100001100100000000000000000000;
			// PEs: 32, 38 -> 39
			// srcs: (2045, 34)(3140) 47, (535) 2 --> (3672) 94:PEGB0, ND6, *, PENB
			10'd52 : rdata = 48'b000111110000000001100000110000000000000100000000;
			// PEs: 38, 38 -> 38
			// srcs: (2046, 49)(3) 1, (3670) 0 --> (4454) 0:NM0, NI0, *, NI1
			10'd53 : rdata = 48'b000111000000000010100000000100001000000000000000;
			// PEs: 38, 37 -> 37
			// srcs: (2047, 50)(3) 1, (3671) 47 --> (4455) 47:NM0, PENB, *, PEGB5
			10'd54 : rdata = 48'b000111000000000011011111110000000000000011010000;
			// PEs: 38, 38 -> 38
			// srcs: (2049, 64)(1318) -2, (4454) 0 --> (5238) -2:NW12, NI1, -, NW12
			10'd55 : rdata = 48'b000100100000110010100000001000000111000000000000;
			// PEs: 38, 39 -> 38
			// srcs: (2054, 65)(1320) 0, (4456) 94 --> (5240) -94:NW6, PEGB7, -, NW6
			10'd56 : rdata = 48'b000100100000011011100001110000000101100000000000;
			// PEs: 32, 38 -> 38
			// srcs: (2125, 35)(3140) 47, (615) 1 --> (3752) 47:PEGB0, ND7, *, NI0
			10'd57 : rdata = 48'b000111110000000001100000111100000000000000000000;
			// PEs: 38, 37 -> 37
			// srcs: (2127, 51)(3) 1, (3751) -47 --> (4535) -47:NM0, PENB, *, PEGB5
			10'd58 : rdata = 48'b000111000000000011011111110000000000000011010000;
			// PEs: 38, 38 -> 
			// srcs: (2128, 52)(3) 1, (3752) 47 --> (4536) 47:NM0, NI0, *, 
			10'd59 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 38, 38 -> 38
			// srcs: (2131, 66)(1400) -3, (4536) 47 --> (5320) -50:NW7, ALU, -, NW7
			10'd60 : rdata = 48'b000100100000011100111111111000000101110000000000;
			// PEs: 32, 38 -> 
			// srcs: (2205, 36)(3140) 47, (695) 1 --> (3832) 47:PEGB0, ND8, *, 
			10'd61 : rdata = 48'b000111110000000001100001000000000000000000000000;
			// PEs: 38, 38 -> 
			// srcs: (2208, 53)(3) 1, (3832) 47 --> (4616) 47:NM0, ALU, *, 
			10'd62 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 38, 38 -> 38
			// srcs: (2211, 67)(1480) -1, (4616) 47 --> (5400) -48:NW8, ALU, -, NW8
			10'd63 : rdata = 48'b000100100000100000111111111000000110000000000000;
			// PEs: 32, 38 -> 
			// srcs: (2227, 37)(3140) 47, (717) 1 --> (3854) 47:PEGB0, ND13, *, 
			10'd64 : rdata = 48'b000111110000000001100001101000000000000000000000;
			// PEs: 38, 38 -> 
			// srcs: (2230, 54)(3) 1, (3854) 47 --> (4638) 47:NM0, ALU, *, 
			10'd65 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 38, 38 -> 38
			// srcs: (2233, 68)(1502) -1, (4638) 47 --> (5422) -48:NW13, ALU, -, NW13
			10'd66 : rdata = 48'b000100100000110100111111111000000111010000000000;
			// PEs: 32, 38 -> 
			// srcs: (2287, 38)(3140) 47, (777) 1 --> (3914) 47:PEGB0, ND9, *, 
			10'd67 : rdata = 48'b000111110000000001100001001000000000000000000000;
			// PEs: 38, 38 -> 
			// srcs: (2290, 55)(3) 1, (3914) 47 --> (4698) 47:NM0, ALU, *, 
			10'd68 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 38, 38 -> 38
			// srcs: (2293, 69)(1562) 1, (4698) 47 --> (5482) -46:NW9, ALU, -, NW9
			10'd69 : rdata = 48'b000100100000100100111111111000000110010000000000;
			default : rdata = 48'b000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 39) begin
	always @(*) begin
		case(address)
			// PEs: 39, 39 -> 32
			// srcs: (1, 0)(53) -3, (838) 2 --> (1622) -6:ND0, NW0, *, PENB
			10'd0 : rdata = 48'b000110110000000001000000000000000000000100000000;
			// PEs: 39, 39 -> 32
			// srcs: (2, 1)(133) -2, (918) 2 --> (1702) -4:ND1, NW1, *, PENB
			10'd1 : rdata = 48'b000110110000000101000000001000000000000100000000;
			// PEs: 39, 39 -> 32
			// srcs: (3, 2)(213) -1, (998) -3 --> (1782) 3:ND2, NW2, *, PENB
			10'd2 : rdata = 48'b000110110000001001000000010000000000000100000000;
			// PEs: 39, 39 -> 32
			// srcs: (4, 3)(295) 1, (1080) 1 --> (1864) 1:ND3, NW3, *, PENB
			10'd3 : rdata = 48'b000110110000001101000000011000000000000100000000;
			// PEs: 39, 39 -> 32
			// srcs: (5, 4)(375) -2, (1160) -2 --> (1944) 4:ND4, NW4, *, PENB
			10'd4 : rdata = 48'b000110110000010001000000100000000000000100000000;
			// PEs: 39, 39 -> 32
			// srcs: (6, 5)(455) 2, (1240) 0 --> (2024) 0:ND5, NW5, *, PENB
			10'd5 : rdata = 48'b000110110000010101000000101000000000000100000000;
			// PEs: 39, 39 -> 32
			// srcs: (7, 6)(537) -3, (1322) 2 --> (2106) -6:ND6, NW6, *, PENB
			10'd6 : rdata = 48'b000110110000011001000000110000000000000100000000;
			// PEs: 39, 39 -> 32
			// srcs: (8, 7)(617) -1, (1402) -3 --> (2186) 3:ND7, NW7, *, PENB
			10'd7 : rdata = 48'b000110110000011101000000111000000000000100000000;
			// PEs: 39, 39 -> 32
			// srcs: (9, 8)(697) -3, (1482) 1 --> (2266) -3:ND8, NW8, *, PENB
			10'd8 : rdata = 48'b000110110000100001000001000000000000000100000000;
			// PEs: 39, 39 -> 32
			// srcs: (10, 9)(779) 1, (1564) -2 --> (2348) -2:ND9, NW9, *, PENB
			10'd9 : rdata = 48'b000110110000100101000001001000000000000100000000;
			// PEs: 39, 39 -> 32
			// srcs: (11, 10)(172) 1, (957) 0 --> (1741) 0:ND10, NW10, *, PENB
			10'd10 : rdata = 48'b000110110000101001000001010000000000000100000000;
			// PEs: 39, 39 -> 38
			// srcs: (12, 11)(356) -1, (1141) -2 --> (1925) 2:ND11, NW11, *, PEGB6
			10'd11 : rdata = 48'b000110110000101101000001011000000000000011100000;
			// PEs: 39, 39 -> 39
			// srcs: (13, 12)(536) 1, (1321) -1 --> (2105) -1:ND12, NW12, *, NI0
			10'd12 : rdata = 48'b000110110000110001000001100100000000000000000000;
			// PEs: 39, 39 -> 39
			// srcs: (14, 13)(720) 0, (1505) -2 --> (2289) 0:ND13, NW13, *, NI1
			10'd13 : rdata = 48'b000110110000110101000001101100001000000000000000;
			// PEs: 37, 38 -> 33
			// srcs: (15, 16)(2263) -4, (2264) -1 --> (3043) -5:PEGB5, PENB, +, PEGB1
			10'd14 : rdata = 48'b000011110000101011011111110000000000000010010000;
			// PEs: 36 -> 
			// srcs: (16, 17)(2343) 0 --> (2343) 0:PEGB4, pass, 
			10'd15 : rdata = 48'b110001110000100000000000000000000000000000000000;
			// PEs: 35, 39 -> 39
			// srcs: (18, 18)(2342) -4, (2343) 0 --> (3119) -4:PEGB3, ALU, +, NI2
			10'd16 : rdata = 48'b000011110000011000111111111100010000000000000000;
			// PEs: 32 -> 
			// srcs: (58, 14)(1767) 0 --> (1767) 0:PEGB0, pass, 
			10'd17 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 32, 39 -> 32
			// srcs: (67, 15)(1766) -3, (1767) 0 --> (2544) -3:PEGB0, ALU, +, PENB
			10'd18 : rdata = 48'b000011110000000000111111111000000000000100000000;
			// PEs: 33 -> 
			// srcs: (135, 19)(2871) 0 --> (2871) 0:PEGB1, pass, 
			10'd19 : rdata = 48'b110001110000001000000000000000000000000000000000;
			// PEs: 39, 35 -> 35
			// srcs: (138, 20)(2871) 0, (2093) 2 --> (2872) 2:ALU, PEGB3, +, PEGB3
			10'd20 : rdata = 48'b000010011111111111100000110000000000000010110000;
			// PEs: 39 -> 32
			// srcs: (141, 23)(3119) -4 --> (3119) -4:NI2, pass, PENB
			10'd21 : rdata = 48'b110001010000001000000000000000000000000100000000;
			// PEs: 39 -> 32
			// srcs: (171, 22)(2289) 0 --> (2289) 0:NI1, pass, PENB
			10'd22 : rdata = 48'b110001010000000100000000000000000000000100000000;
			// PEs: 39 -> 32
			// srcs: (317, 21)(2105) -1 --> (2105) -1:NI0, pass, PENB
			10'd23 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 38, 33 -> 32
			// srcs: (419, 24)(3042) -6, (3044) -3 --> (3045) -9:PENB, PEGB1, +, PENB
			10'd24 : rdata = 48'b000011101111111011100000010000000000000100000000;
			// PEs: 32, 39 -> 39
			// srcs: (1563, 25)(3140) 47, (53) -3 --> (3190) -141:PEGB0, ND0, *, NI0
			10'd25 : rdata = 48'b000111110000000001100000000100000000000000000000;
			// PEs: 39, 38 -> 38
			// srcs: (1564, 39)(3) 1, (3188) 0 --> (3972) 0:NM0, PENB, *, PEGB6
			10'd26 : rdata = 48'b000111000000000011011111110000000000000011100000;
			// PEs: 39, 39 -> 
			// srcs: (1566, 40)(3) 1, (3190) -141 --> (3974) -141:NM0, NI0, *, 
			10'd27 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 39, 39 -> 39
			// srcs: (1569, 57)(838) 2, (3974) -141 --> (4758) 143:NW0, ALU, -, NW0
			10'd28 : rdata = 48'b000100100000000000111111111000000100000000000000;
			// PEs: 32, 39 -> 
			// srcs: (1643, 26)(3140) 47, (133) -2 --> (3270) -94:PEGB0, ND1, *, 
			10'd29 : rdata = 48'b000111110000000001100000001000000000000000000000;
			// PEs: 39, 39 -> 
			// srcs: (1646, 41)(3) 1, (3270) -94 --> (4054) -94:NM0, ALU, *, 
			10'd30 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 39, 39 -> 39
			// srcs: (1649, 58)(918) 2, (4054) -94 --> (4838) 96:NW1, ALU, -, NW1
			10'd31 : rdata = 48'b000100100000000100111111111000000100010000000000;
			// PEs: 32, 39 -> 
			// srcs: (1682, 27)(3140) 47, (172) 1 --> (3309) 47:PEGB0, ND10, *, 
			10'd32 : rdata = 48'b000111110000000001100001010000000000000000000000;
			// PEs: 39, 39 -> 
			// srcs: (1685, 42)(3) 1, (3309) 47 --> (4093) 47:NM0, ALU, *, 
			10'd33 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 39, 39 -> 39
			// srcs: (1688, 59)(957) 0, (4093) 47 --> (4877) -47:NW10, ALU, -, NW10
			10'd34 : rdata = 48'b000100100000101000111111111000000110100000000000;
			// PEs: 32, 39 -> 39
			// srcs: (1723, 28)(3140) 47, (213) -1 --> (3350) -47:PEGB0, ND2, *, NI0
			10'd35 : rdata = 48'b000111110000000001100000010100000000000000000000;
			// PEs: 39, 38 -> 38
			// srcs: (1724, 43)(3) 1, (3348) -141 --> (4132) -141:NM0, PENB, *, PEGB6
			10'd36 : rdata = 48'b000111000000000011011111110000000000000011100000;
			// PEs: 39, 39 -> 
			// srcs: (1726, 44)(3) 1, (3350) -47 --> (4134) -47:NM0, NI0, *, 
			10'd37 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 39, 39 -> 39
			// srcs: (1729, 60)(998) -3, (4134) -47 --> (4918) 44:NW2, ALU, -, NW2
			10'd38 : rdata = 48'b000100100000001000111111111000000100100000000000;
			// PEs: 32, 39 -> 
			// srcs: (1805, 29)(3140) 47, (295) 1 --> (3432) 47:PEGB0, ND3, *, 
			10'd39 : rdata = 48'b000111110000000001100000011000000000000000000000;
			// PEs: 39, 39 -> 
			// srcs: (1808, 45)(3) 1, (3432) 47 --> (4216) 47:NM0, ALU, *, 
			10'd40 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 39, 39 -> 39
			// srcs: (1811, 61)(1080) 1, (4216) 47 --> (5000) -46:NW3, ALU, -, NW3
			10'd41 : rdata = 48'b000100100000001100111111111000000100110000000000;
			// PEs: 32, 39 -> 
			// srcs: (1866, 30)(3140) 47, (356) -1 --> (3493) -47:PEGB0, ND11, *, 
			10'd42 : rdata = 48'b000111110000000001100001011000000000000000000000;
			// PEs: 39, 39 -> 
			// srcs: (1869, 46)(3) 1, (3493) -47 --> (4277) -47:NM0, ALU, *, 
			10'd43 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 39, 39 -> 39
			// srcs: (1872, 62)(1141) -2, (4277) -47 --> (5061) 45:NW11, ALU, -, NW11
			10'd44 : rdata = 48'b000100100000101100111111111000000110110000000000;
			// PEs: 32, 39 -> 
			// srcs: (1885, 31)(3140) 47, (375) -2 --> (3512) -94:PEGB0, ND4, *, 
			10'd45 : rdata = 48'b000111110000000001100000100000000000000000000000;
			// PEs: 39, 39 -> 
			// srcs: (1888, 47)(3) 1, (3512) -94 --> (4296) -94:NM0, ALU, *, 
			10'd46 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 39, 39 -> 39
			// srcs: (1891, 63)(1160) -2, (4296) -94 --> (5080) 92:NW4, ALU, -, NW4
			10'd47 : rdata = 48'b000100100000010000111111111000000101000000000000;
			// PEs: 32, 39 -> 39
			// srcs: (1965, 32)(3140) 47, (455) 2 --> (3592) 94:PEGB0, ND5, *, NI0
			10'd48 : rdata = 48'b000111110000000001100000101100000000000000000000;
			// PEs: 39, 38 -> 38
			// srcs: (1966, 48)(3) 1, (3590) 0 --> (4374) 0:NM0, PENB, *, PEGB6
			10'd49 : rdata = 48'b000111000000000011011111110000000000000011100000;
			// PEs: 39, 39 -> 
			// srcs: (1968, 49)(3) 1, (3592) 94 --> (4376) 94:NM0, NI0, *, 
			10'd50 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 39, 39 -> 39
			// srcs: (1971, 64)(1240) 0, (4376) 94 --> (5160) -94:NW5, ALU, -, NW5
			10'd51 : rdata = 48'b000100100000010100111111111000000101010000000000;
			// PEs: 32, 39 -> 39
			// srcs: (2046, 33)(3140) 47, (536) 1 --> (3673) 47:PEGB0, ND12, *, NI0
			10'd52 : rdata = 48'b000111110000000001100001100100000000000000000000;
			// PEs: 32, 39 -> 39
			// srcs: (2047, 34)(3140) 47, (537) -3 --> (3674) -141:PEGB0, ND6, *, NI1
			10'd53 : rdata = 48'b000111110000000001100000110100001000000000000000;
			// PEs: 39, 38 -> 38
			// srcs: (2048, 50)(3) 1, (3672) 94 --> (4456) 94:NM0, PENB, *, PEGB6
			10'd54 : rdata = 48'b000111000000000011011111110000000000000011100000;
			// PEs: 39, 39 -> 39
			// srcs: (2049, 51)(3) 1, (3673) 47 --> (4457) 47:NM0, NI0, *, NI2
			10'd55 : rdata = 48'b000111000000000010100000000100010000000000000000;
			// PEs: 39, 39 -> 39
			// srcs: (2050, 52)(3) 1, (3674) -141 --> (4458) -141:NM0, NI1, *, NI0
			10'd56 : rdata = 48'b000111000000000010100000001100000000000000000000;
			// PEs: 39, 39 -> 39
			// srcs: (2052, 65)(1321) -1, (4457) 47 --> (5241) -48:NW12, NI2, -, NW12
			10'd57 : rdata = 48'b000100100000110010100000010000000111000000000000;
			// PEs: 39, 39 -> 39
			// srcs: (2053, 66)(1322) 2, (4458) -141 --> (5242) 143:NW6, NI0, -, NW6
			10'd58 : rdata = 48'b000100100000011010100000000000000101100000000000;
			// PEs: 32, 39 -> 
			// srcs: (2127, 35)(3140) 47, (617) -1 --> (3754) -47:PEGB0, ND7, *, 
			10'd59 : rdata = 48'b000111110000000001100000111000000000000000000000;
			// PEs: 39, 39 -> 
			// srcs: (2130, 53)(3) 1, (3754) -47 --> (4538) -47:NM0, ALU, *, 
			10'd60 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 39, 39 -> 39
			// srcs: (2133, 67)(1402) -3, (4538) -47 --> (5322) 44:NW7, ALU, -, NW7
			10'd61 : rdata = 48'b000100100000011100111111111000000101110000000000;
			// PEs: 32, 39 -> 
			// srcs: (2207, 36)(3140) 47, (697) -3 --> (3834) -141:PEGB0, ND8, *, 
			10'd62 : rdata = 48'b000111110000000001100001000000000000000000000000;
			// PEs: 39, 39 -> 
			// srcs: (2210, 54)(3) 1, (3834) -141 --> (4618) -141:NM0, ALU, *, 
			10'd63 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 39, 39 -> 39
			// srcs: (2213, 68)(1482) 1, (4618) -141 --> (5402) 142:NW8, ALU, -, NW8
			10'd64 : rdata = 48'b000100100000100000111111111000000110000000000000;
			// PEs: 32, 39 -> 
			// srcs: (2230, 37)(3140) 47, (720) 0 --> (3857) 0:PEGB0, ND13, *, 
			10'd65 : rdata = 48'b000111110000000001100001101000000000000000000000;
			// PEs: 39, 39 -> 
			// srcs: (2233, 55)(3) 1, (3857) 0 --> (4641) 0:NM0, ALU, *, 
			10'd66 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 39, 39 -> 39
			// srcs: (2236, 69)(1505) -2, (4641) 0 --> (5425) -2:NW13, ALU, -, NW13
			10'd67 : rdata = 48'b000100100000110100111111111000000111010000000000;
			// PEs: 32, 39 -> 
			// srcs: (2289, 38)(3140) 47, (779) 1 --> (3916) 47:PEGB0, ND9, *, 
			10'd68 : rdata = 48'b000111110000000001100001001000000000000000000000;
			// PEs: 39, 39 -> 
			// srcs: (2292, 56)(3) 1, (3916) 47 --> (4700) 47:NM0, ALU, *, 
			10'd69 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 39, 39 -> 39
			// srcs: (2295, 70)(1564) -2, (4700) 47 --> (5484) -49:NW9, ALU, -, NW9
			10'd70 : rdata = 48'b000100100000100100111111111000000110010000000000;
			default : rdata = 48'b000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 40) begin
	always @(*) begin
		case(address)
			// PEs: 44 -> 16
			// srcs: (6, 0)(1626) 0 --> (1626) 0:PEGB4, pass, PUGB2
			10'd0 : rdata = 48'b110001110000100000000000000000000000000000001010;
			// PEs: 45 -> 16
			// srcs: (7, 1)(1627) 6 --> (1627) 6:PEGB5, pass, PUGB2
			10'd1 : rdata = 48'b110001110000101000000000000000000000000000001010;
			// PEs: 46 -> 16
			// srcs: (8, 2)(1629) 2 --> (1629) 2:PEGB6, pass, PUGB2
			10'd2 : rdata = 48'b110001110000110000000000000000000000000000001010;
			// PEs: 47 -> 16
			// srcs: (9, 3)(1630) -2 --> (1630) -2:PENB, pass, PUGB2
			10'd3 : rdata = 48'b110001101111111000000000000000000000000000001010;
			// PEs: 41 -> 48
			// srcs: (10, 16)(1703) 3 --> (1703) 3:PEGB1, pass, PUNB
			10'd4 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 42 -> 48
			// srcs: (11, 17)(1705) 6 --> (1705) 6:PEGB2, pass, PUNB
			10'd5 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 43 -> 48
			// srcs: (12, 18)(1706) 2 --> (1706) 2:PEGB3, pass, PUNB
			10'd6 : rdata = 48'b110001110000011000000000000000000000001000000000;
			// PEs: 44 -> 48
			// srcs: (13, 19)(1708) 0 --> (1708) 0:PEGB4, pass, PUNB
			10'd7 : rdata = 48'b110001110000100000000000000000000000001000000000;
			// PEs: 32 -> 40
			// srcs: (14, 7)(1693) 0 --> (1693) 0:PUNB, pass, NI0
			10'd8 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 32 -> 42
			// srcs: (15, 8)(1694) -6 --> (1694) -6:PUNB, pass, PEGB2
			10'd9 : rdata = 48'b110001101111111100000000000000000000000010100000;
			// PEs: 32 -> 40
			// srcs: (16, 10)(1696) 2 --> (1696) 2:PUNB, pass, NI1
			10'd10 : rdata = 48'b110001101111111100000000000100001000000000000000;
			// PEs: 32 -> 43
			// srcs: (17, 11)(1697) 2 --> (1697) 2:PUNB, pass, PEGB3
			10'd11 : rdata = 48'b110001101111111100000000000000000000000010110000;
			// PEs: 32 -> 40
			// srcs: (18, 13)(1699) 0 --> (1699) 0:PUNB, pass, NI2
			10'd12 : rdata = 48'b110001101111111100000000000100010000000000000000;
			// PEs: 32 -> 44
			// srcs: (19, 14)(1700) -2 --> (1700) -2:PUNB, pass, PEGB4
			10'd13 : rdata = 48'b110001101111111100000000000000000000000011000000;
			// PEs: 45 -> 48
			// srcs: (20, 20)(1709) 0 --> (1709) 0:PEGB5, pass, PUNB
			10'd14 : rdata = 48'b110001110000101000000000000000000000001000000000;
			// PEs: 46 -> 48
			// srcs: (21, 21)(1711) 0 --> (1711) 0:PEGB6, pass, PUNB
			10'd15 : rdata = 48'b110001110000110000000000000000000000001000000000;
			// PEs: 47 -> 48
			// srcs: (22, 22)(1712) -6 --> (1712) -6:PENB, pass, PUNB
			10'd16 : rdata = 48'b110001101111111000000000000000000000001000000000;
			// PEs: 32 -> 40
			// srcs: (23, 23)(1773) 0 --> (1773) 0:PUNB, pass, NI3
			10'd17 : rdata = 48'b110001101111111100000000000100011000000000000000;
			// PEs: 40 -> 42
			// srcs: (24, 9)(1693) 0 --> (1693) 0:NI0, pass, PEGB2
			10'd18 : rdata = 48'b110001010000000000000000000000000000000010100000;
			// PEs: 32 -> 45
			// srcs: (25, 24)(1774) 1 --> (1774) 1:PUNB, pass, PEGB5
			10'd19 : rdata = 48'b110001101111111100000000000000000000000011010000;
			// PEs: 40 -> 43
			// srcs: (26, 12)(1696) 2 --> (1696) 2:NI1, pass, PEGB3
			10'd20 : rdata = 48'b110001010000000100000000000000000000000010110000;
			// PEs: 32 -> 40
			// srcs: (27, 26)(1776) 9 --> (1776) 9:PUNB, pass, NI0
			10'd21 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 40 -> 44
			// srcs: (28, 15)(1699) 0 --> (1699) 0:NI2, pass, PEGB4
			10'd22 : rdata = 48'b110001010000001000000000000000000000000011000000;
			// PEs: 32 -> 46
			// srcs: (29, 27)(1777) 2 --> (1777) 2:PUNB, pass, PEGB6
			10'd23 : rdata = 48'b110001101111111100000000000000000000000011100000;
			// PEs: 32 -> 40
			// srcs: (30, 29)(1779) 0 --> (1779) 0:PUNB, pass, NI1
			10'd24 : rdata = 48'b110001101111111100000000000100001000000000000000;
			// PEs: 32 -> 47
			// srcs: (31, 30)(1780) -6 --> (1780) -6:PUNB, pass, PEGB7
			10'd25 : rdata = 48'b110001101111111100000000000000000000000011110000;
			// PEs: 41 -> 48
			// srcs: (32, 32)(1783) 2 --> (1783) 2:PEGB1, pass, PUNB
			10'd26 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 42 -> 48
			// srcs: (33, 33)(1785) 2 --> (1785) 2:PEGB2, pass, PUNB
			10'd27 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 40 -> 45
			// srcs: (34, 25)(1773) 0 --> (1773) 0:NI3, pass, PEGB5
			10'd28 : rdata = 48'b110001010000001100000000000000000000000011010000;
			// PEs: 8 -> 40
			// srcs: (35, 4)(1665) -1 --> (1665) -1:PUGB1, pass, NI2
			10'd29 : rdata = 48'b110001110000001100000000000100010000000000000000;
			// PEs: 43 -> 48
			// srcs: (36, 34)(1786) 2 --> (1786) 2:PEGB3, pass, PUNB
			10'd30 : rdata = 48'b110001110000011000000000000000000000001000000000;
			// PEs: 8 -> 41
			// srcs: (37, 5)(1666) 0 --> (1666) 0:PUGB1, pass, PENB
			10'd31 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 40 -> 46
			// srcs: (38, 28)(1776) 9 --> (1776) 9:NI0, pass, PEGB6
			10'd32 : rdata = 48'b110001010000000000000000000000000000000011100000;
			// PEs: 44 -> 16
			// srcs: (39, 35)(1788) 3 --> (1788) 3:PEGB4, pass, PUGB2
			10'd33 : rdata = 48'b110001110000100000000000000000000000000000001010;
			// PEs: 40 -> 47
			// srcs: (40, 31)(1779) 0 --> (1779) 0:NI1, pass, PEGB7
			10'd34 : rdata = 48'b110001010000000100000000000000000000000011110000;
			// PEs: 45 -> 16
			// srcs: (41, 36)(1789) 4 --> (1789) 4:PEGB5, pass, PUGB2
			10'd35 : rdata = 48'b110001110000101000000000000000000000000000001010;
			// PEs: 46 -> 24
			// srcs: (42, 37)(1791) 0 --> (1791) 0:PEGB6, pass, PUGB3
			10'd36 : rdata = 48'b110001110000110000000000000000000000000000001011;
			// PEs: 40 -> 41
			// srcs: (43, 6)(1665) -1 --> (1665) -1:NI2, pass, PENB
			10'd37 : rdata = 48'b110001010000001000000000000000000000000100000000;
			// PEs: 47 -> 24
			// srcs: (44, 38)(1792) 0 --> (1792) 0:PENB, pass, PUGB3
			10'd38 : rdata = 48'b110001101111111000000000000000000000000000001011;
			// PEs: 32 -> 40
			// srcs: (45, 39)(1855) 4 --> (1855) 4:PUNB, pass, NI0
			10'd39 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 32 -> 42
			// srcs: (46, 40)(1856) 0 --> (1856) 0:PUNB, pass, PEGB2
			10'd40 : rdata = 48'b110001101111111100000000000000000000000010100000;
			// PEs: 32 -> 40
			// srcs: (47, 42)(1858) 2 --> (1858) 2:PUNB, pass, NI1
			10'd41 : rdata = 48'b110001101111111100000000000100001000000000000000;
			// PEs: 32 -> 43
			// srcs: (48, 43)(1859) -4 --> (1859) -4:PUNB, pass, PEGB3
			10'd42 : rdata = 48'b110001101111111100000000000000000000000010110000;
			// PEs: 32 -> 40
			// srcs: (49, 45)(1861) 1 --> (1861) 1:PUNB, pass, NI2
			10'd43 : rdata = 48'b110001101111111100000000000100010000000000000000;
			// PEs: 32 -> 44
			// srcs: (50, 46)(1862) 0 --> (1862) 0:PUNB, pass, PEGB4
			10'd44 : rdata = 48'b110001101111111100000000000000000000000011000000;
			// PEs: 41 -> 48
			// srcs: (51, 48)(1865) -3 --> (1865) -3:PEGB1, pass, PUNB
			10'd45 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 46 -> 48
			// srcs: (52, 49)(1871) 0 --> (1871) 0:PEGB6, pass, PUNB
			10'd46 : rdata = 48'b110001110000110000000000000000000000001000000000;
			// PEs: 47 -> 48
			// srcs: (53, 50)(1872) 3 --> (1872) 3:PENB, pass, PUNB
			10'd47 : rdata = 48'b110001101111111000000000000000000000001000000000;
			// PEs: 48 -> 40
			// srcs: (54, 51)(1877) 0 --> (1877) 0:PUGB6, pass, NI3
			10'd48 : rdata = 48'b110001110000110100000000000100011000000000000000;
			// PEs: 40 -> 42
			// srcs: (55, 41)(1855) 4 --> (1855) 4:NI0, pass, PEGB2
			10'd49 : rdata = 48'b110001010000000000000000000000000000000010100000;
			// PEs: 48 -> 41
			// srcs: (56, 52)(1878) -2 --> (1878) -2:PUGB6, pass, PENB
			10'd50 : rdata = 48'b110001110000110100000000000000000000000100000000;
			// PEs: 40 -> 43
			// srcs: (57, 44)(1858) 2 --> (1858) 2:NI1, pass, PEGB3
			10'd51 : rdata = 48'b110001010000000100000000000000000000000010110000;
			// PEs: 42 -> 48
			// srcs: (58, 64)(1947) 1 --> (1947) 1:PEGB2, pass, PUNB
			10'd52 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 40 -> 44
			// srcs: (59, 47)(1861) 1 --> (1861) 1:NI2, pass, PEGB4
			10'd53 : rdata = 48'b110001010000001000000000000000000000000011000000;
			// PEs: 43 -> 48
			// srcs: (60, 65)(1948) -2 --> (1948) -2:PEGB3, pass, PUNB
			10'd54 : rdata = 48'b110001110000011000000000000000000000001000000000;
			// PEs: 44 -> 48
			// srcs: (61, 66)(1950) 9 --> (1950) 9:PEGB4, pass, PUNB
			10'd55 : rdata = 48'b110001110000100000000000000000000000001000000000;
			// PEs: 40 -> 41
			// srcs: (62, 53)(1877) 0 --> (1877) 0:NI3, pass, PENB
			10'd56 : rdata = 48'b110001010000001100000000000000000000000100000000;
			// PEs: 32 -> 40
			// srcs: (63, 54)(1935) 4 --> (1935) 4:PUNB, pass, NI0
			10'd57 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 32 -> 41
			// srcs: (64, 55)(1936) -3 --> (1936) -3:PUNB, pass, PENB
			10'd58 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 45 -> 48
			// srcs: (65, 67)(1951) 6 --> (1951) 6:PEGB5, pass, PUNB
			10'd59 : rdata = 48'b110001110000101000000000000000000000001000000000;
			// PEs: 46 -> 48
			// srcs: (66, 68)(1953) -3 --> (1953) -3:PEGB6, pass, PUNB
			10'd60 : rdata = 48'b110001110000110000000000000000000000001000000000;
			// PEs: 47 -> 48
			// srcs: (67, 69)(1954) 3 --> (1954) 3:PENB, pass, PUNB
			10'd61 : rdata = 48'b110001101111111000000000000000000000001000000000;
			// PEs: 42 -> 48
			// srcs: (68, 77)(2027) -6 --> (2027) -6:PEGB2, pass, PUNB
			10'd62 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 43 -> 48
			// srcs: (69, 78)(2028) 0 --> (2028) 0:PEGB3, pass, PUNB
			10'd63 : rdata = 48'b110001110000011000000000000000000000001000000000;
			// PEs: 40 -> 41
			// srcs: (70, 56)(1935) 4 --> (1935) 4:NI0, pass, PENB
			10'd64 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 32 -> 40
			// srcs: (71, 57)(1938) -2 --> (1938) -2:PUNB, pass, NI0
			10'd65 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 32 -> 41
			// srcs: (72, 58)(1939) -1 --> (1939) -1:PUNB, pass, PENB
			10'd66 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 44 -> 48
			// srcs: (73, 79)(2030) -1 --> (2030) -1:PEGB4, pass, PUNB
			10'd67 : rdata = 48'b110001110000100000000000000000000000001000000000;
			// PEs: 45 -> 48
			// srcs: (74, 80)(2031) -2 --> (2031) -2:PEGB5, pass, PUNB
			10'd68 : rdata = 48'b110001110000101000000000000000000000001000000000;
			// PEs: 46 -> 48
			// srcs: (75, 81)(2033) 9 --> (2033) 9:PEGB6, pass, PUNB
			10'd69 : rdata = 48'b110001110000110000000000000000000000001000000000;
			// PEs: 47 -> 48
			// srcs: (76, 82)(2034) 1 --> (2034) 1:PENB, pass, PUNB
			10'd70 : rdata = 48'b110001101111111000000000000000000000001000000000;
			// PEs: 42 -> 48
			// srcs: (77, 93)(2109) 6 --> (2109) 6:PEGB2, pass, PUNB
			10'd71 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 40 -> 41
			// srcs: (78, 59)(1938) -2 --> (1938) -2:NI0, pass, PENB
			10'd72 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 32 -> 40
			// srcs: (79, 60)(1941) 0 --> (1941) 0:PUNB, pass, NI0
			10'd73 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 32 -> 41
			// srcs: (80, 61)(1942) 2 --> (1942) 2:PUNB, pass, PENB
			10'd74 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 32 -> 45
			// srcs: (81, 63)(1944) 4 --> (1944) 4:PUNB, pass, PEGB5
			10'd75 : rdata = 48'b110001101111111100000000000000000000000011010000;
			// PEs: 43 -> 48
			// srcs: (82, 94)(2110) 6 --> (2110) 6:PEGB3, pass, PUNB
			10'd76 : rdata = 48'b110001110000011000000000000000000000001000000000;
			// PEs: 42 -> 48
			// srcs: (83, 105)(2189) -2 --> (2189) -2:PEGB2, pass, PUNB
			10'd77 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 43 -> 48
			// srcs: (84, 106)(2190) -2 --> (2190) -2:PEGB3, pass, PUNB
			10'd78 : rdata = 48'b110001110000011000000000000000000000001000000000;
			// PEs: 44 -> 48
			// srcs: (85, 107)(2192) -3 --> (2192) -3:PEGB4, pass, PUNB
			10'd79 : rdata = 48'b110001110000100000000000000000000000001000000000;
			// PEs: 40 -> 41
			// srcs: (86, 62)(1941) 0 --> (1941) 0:NI0, pass, PENB
			10'd80 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 32 -> 40
			// srcs: (87, 70)(2018) -2 --> (2018) -2:PUNB, pass, NI0
			10'd81 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 32 -> 41
			// srcs: (88, 71)(2019) 0 --> (2019) 0:PUNB, pass, PENB
			10'd82 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 45 -> 48
			// srcs: (89, 108)(2193) -6 --> (2193) -6:PEGB5, pass, PUNB
			10'd83 : rdata = 48'b110001110000101000000000000000000000001000000000;
			// PEs: 46 -> 48
			// srcs: (90, 109)(2195) -2 --> (2195) -2:PEGB6, pass, PUNB
			10'd84 : rdata = 48'b110001110000110000000000000000000000001000000000;
			// PEs: 47 -> 48
			// srcs: (91, 110)(2196) 2 --> (2196) 2:PENB, pass, PUNB
			10'd85 : rdata = 48'b110001101111111000000000000000000000001000000000;
			// PEs: 46 -> 0
			// srcs: (92, 127)(1579) -6 --> (1579) -6:PEGB6, pass, PUGB0
			10'd86 : rdata = 48'b110001110000110000000000000000000000000000001000;
			// PEs: 47 -> 0
			// srcs: (93, 128)(1582) -6 --> (1582) -6:PENB, pass, PUGB0
			10'd87 : rdata = 48'b110001101111111000000000000000000000000000001000;
			// PEs: 40 -> 41
			// srcs: (94, 72)(2018) -2 --> (2018) -2:NI0, pass, PENB
			10'd88 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 32 -> 40
			// srcs: (95, 73)(2021) 2 --> (2021) 2:PUNB, pass, NI0
			10'd89 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 32 -> 41
			// srcs: (96, 74)(2022) 0 --> (2022) 0:PUNB, pass, PENB
			10'd90 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 32 -> 46
			// srcs: (97, 76)(2024) 0 --> (2024) 0:PUNB, pass, PEGB6
			10'd91 : rdata = 48'b110001101111111100000000000000000000000011100000;
			// PEs: 43 -> 32
			// srcs: (98, 137)(2478) 4 --> (2478) 4:PEGB3, pass, PUGB4
			10'd92 : rdata = 48'b110001110000011000000000000000000000000000001100;
			// PEs: 41 -> 56
			// srcs: (99, 113)(1623) 0 --> (1623) 0:PEGB1, pass, PUGB7
			10'd93 : rdata = 48'b110001110000001000000000000000000000000000001111;
			// PEs: 42 -> 8
			// srcs: (100, 114)(1624) 0 --> (1624) 0:PEGB2, pass, PUGB1
			10'd94 : rdata = 48'b110001110000010000000000000000000000000000001001;
			// PEs: 42 -> 48
			// srcs: (101, 116)(1867) 6 --> (1867) 6:PEGB2, pass, PUNB
			10'd95 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 40 -> 41
			// srcs: (102, 75)(2021) 2 --> (2021) 2:NI0, pass, PENB
			10'd96 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 32 -> 40
			// srcs: (103, 83)(2097) 6 --> (2097) 6:PUNB, pass, NI0
			10'd97 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 32 -> 41
			// srcs: (104, 84)(2098) 0 --> (2098) 0:PUNB, pass, PENB
			10'd98 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 46 -> 16
			// srcs: (105, 150)(1759) 2 --> (1759) 2:PEGB6, pass, PUGB2
			10'd99 : rdata = 48'b110001110000110000000000000000000000000000001010;
			// PEs: 41 -> 0
			// srcs: (106, 181)(2799) -2 --> (2799) -2:PEGB1, pass, PUGB0
			10'd100 : rdata = 48'b110001110000001000000000000000000000000000001000;
			// PEs: 43 -> 8
			// srcs: (108, 115)(1625) 4 --> (1625) 4:PEGB3, pass, PUGB1
			10'd101 : rdata = 48'b110001110000011000000000000000000000000000001001;
			// PEs: 44 -> 8
			// srcs: (109, 148)(1753) -4 --> (1753) -4:PEGB4, pass, PUGB1
			10'd102 : rdata = 48'b110001110000100000000000000000000000000000001001;
			// PEs: 40 -> 41
			// srcs: (110, 85)(2097) 6 --> (2097) 6:NI0, pass, PENB
			10'd103 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 32 -> 40
			// srcs: (111, 86)(2100) -3 --> (2100) -3:PUNB, pass, NI0
			10'd104 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 32 -> 41
			// srcs: (112, 87)(2101) 6 --> (2101) 6:PUNB, pass, PENB
			10'd105 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 43 -> 48
			// srcs: (113, 117)(1868) -1 --> (1868) -1:PEGB3, pass, PUNB
			10'd106 : rdata = 48'b110001110000011000000000000000000000001000000000;
			// PEs: 41 -> 56
			// srcs: (114, 135)(2445) -1 --> (2445) -1:PEGB1, pass, PUGB7
			10'd107 : rdata = 48'b110001110000001000000000000000000000000000001111;
			// PEs: 42 -> 24
			// srcs: (115, 146)(1747) 0 --> (1747) 0:PEGB2, pass, PUGB3
			10'd108 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 43 -> 32
			// srcs: (116, 147)(1750) 0 --> (1750) 0:PEGB3, pass, PUGB4
			10'd109 : rdata = 48'b110001110000011000000000000000000000000000001100;
			// PEs: 47 -> 24
			// srcs: (117, 151)(1762) 0 --> (1762) 0:PENB, pass, PUGB3
			10'd110 : rdata = 48'b110001101111111000000000000000000000000000001011;
			// PEs: 40 -> 41
			// srcs: (118, 88)(2100) -3 --> (2100) -3:NI0, pass, PENB
			10'd111 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 32 -> 40
			// srcs: (119, 89)(2103) 0 --> (2103) 0:PUNB, pass, NI0
			10'd112 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 32 -> 41
			// srcs: (120, 90)(2104) 0 --> (2104) 0:PUNB, pass, PENB
			10'd113 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 32 -> 47
			// srcs: (121, 92)(2106) -6 --> (2106) -6:PUNB, pass, PEGB7
			10'd114 : rdata = 48'b110001101111111100000000000000000000000011110000;
			// PEs: 44 -> 48
			// srcs: (122, 118)(1869) 0 --> (1869) 0:PEGB4, pass, PUNB
			10'd115 : rdata = 48'b110001110000100000000000000000000000001000000000;
			// PEs: 41 -> 56
			// srcs: (123, 145)(1744) 1 --> (1744) 1:PEGB1, pass, PUGB7
			10'd116 : rdata = 48'b110001110000001000000000000000000000000000001111;
			// PEs: 45 -> 8
			// srcs: (124, 190)(2124) -3 --> (2124) -3:PEGB5, pass, PUGB1
			10'd117 : rdata = 48'b110001110000101000000000000000000000000000001001;
			// PEs: 47 -> 8
			// srcs: (125, 192)(2130) -4 --> (2130) -4:PENB, pass, PUGB1
			10'd118 : rdata = 48'b110001101111111000000000000000000000000000001001;
			// PEs: 40 -> 41
			// srcs: (126, 91)(2103) 0 --> (2103) 0:NI0, pass, PENB
			10'd119 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 32 -> 40
			// srcs: (127, 95)(2177) 0 --> (2177) 0:PUNB, pass, NI0
			10'd120 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 32 -> 41
			// srcs: (128, 96)(2178) 3 --> (2178) 3:PUNB, pass, PENB
			10'd121 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 45 -> 48
			// srcs: (130, 119)(1870) 0 --> (1870) 0:PEGB5, pass, PUNB
			10'd122 : rdata = 48'b110001110000101000000000000000000000001000000000;
			// PEs: 44 -> 24
			// srcs: (131, 163)(2640) 1 --> (2640) 1:PEGB4, pass, PUGB3
			10'd123 : rdata = 48'b110001110000100000000000000000000000000000001011;
			// PEs: 41 -> 16
			// srcs: (132, 182)(2802) 2 --> (2802) 2:PEGB1, pass, PUGB2
			10'd124 : rdata = 48'b110001110000001000000000000000000000000000001010;
			// PEs: 43 -> 56
			// srcs: (133, 188)(2118) -2 --> (2118) -2:PEGB3, pass, PUGB7
			10'd125 : rdata = 48'b110001110000011000000000000000000000000000001111;
			// PEs: 40 -> 41
			// srcs: (134, 97)(2177) 0 --> (2177) 0:NI0, pass, PENB
			10'd126 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 32 -> 40
			// srcs: (135, 98)(2180) 0 --> (2180) 0:PUNB, pass, NI0
			10'd127 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 32 -> 41
			// srcs: (136, 99)(2181) 2 --> (2181) 2:PUNB, pass, PENB
			10'd128 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 42 -> 8
			// srcs: (137, 214)(2295) 1 --> (2295) 1:PEGB2, pass, PUGB1
			10'd129 : rdata = 48'b110001110000010000000000000000000000000000001001;
			// PEs: 44 -> 48
			// srcs: (138, 123)(2112) 9 --> (2112) 9:PEGB4, pass, PUNB
			10'd130 : rdata = 48'b110001110000100000000000000000000000001000000000;
			// PEs: 44 -> 0
			// srcs: (139, 216)(2301) 0 --> (2301) 0:PEGB4, pass, PUGB0
			10'd131 : rdata = 48'b110001110000100000000000000000000000000000001000;
			// PEs: 47 -> 8
			// srcs: (140, 219)(2314) 4 --> (2314) 4:PENB, pass, PUGB1
			10'd132 : rdata = 48'b110001101111111000000000000000000000000000001001;
			// PEs: 40 -> 41
			// srcs: (142, 100)(2180) 0 --> (2180) 0:NI0, pass, PENB
			10'd133 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 32 -> 40
			// srcs: (143, 101)(2183) -2 --> (2183) -2:PUNB, pass, NI0
			10'd134 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 32 -> 41
			// srcs: (144, 102)(2184) -3 --> (2184) -3:PUNB, pass, PENB
			10'd135 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 44 -> 56
			// srcs: (145, 189)(2121) 0 --> (2121) 0:PEGB4, pass, PUGB7
			10'd136 : rdata = 48'b110001110000100000000000000000000000000000001111;
			// PEs: 45 -> 48
			// srcs: (146, 124)(2113) -1 --> (2113) -1:PEGB5, pass, PUNB
			10'd137 : rdata = 48'b110001110000101000000000000000000000001000000000;
			// PEs: 46 -> 56
			// srcs: (147, 191)(2127) -2 --> (2127) -2:PEGB6, pass, PUGB7
			10'd138 : rdata = 48'b110001110000110000000000000000000000000000001111;
			// PEs: 45 -> 24
			// srcs: (148, 217)(2304) 1 --> (2304) 1:PEGB5, pass, PUGB3
			10'd139 : rdata = 48'b110001110000101000000000000000000000000000001011;
			// PEs: 41 -> 32
			// srcs: (149, 203)(2960) 2 --> (2960) 2:PEGB1, pass, PUGB4
			10'd140 : rdata = 48'b110001110000001000000000000000000000000000001100;
			// PEs: 40 -> 41
			// srcs: (150, 103)(2183) -2 --> (2183) -2:NI0, pass, PENB
			10'd141 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 32 -> 41
			// srcs: (151, 104)(2186) 3 --> (2186) 3:PUNB, pass, PENB
			10'd142 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 32 -> 41
			// srcs: (152, 111)(2266) -3 --> (2266) -3:PUNB, pass, PENB
			10'd143 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 32 -> 41
			// srcs: (153, 112)(2348) -2 --> (2348) -2:PUNB, pass, PENB
			10'd144 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 46 -> 48
			// srcs: (154, 125)(2114) 2 --> (2114) 2:PEGB6, pass, PUNB
			10'd145 : rdata = 48'b110001110000110000000000000000000000001000000000;
			// PEs: 45 -> 8
			// srcs: (155, 224)(3128) 8 --> (3128) 8:PEGB5, pass, PUGB1
			10'd146 : rdata = 48'b110001110000101000000000000000000000000000001001;
			// PEs: 41 -> 56
			// srcs: (157, 204)(2962) -5 --> (2962) -5:PEGB1, pass, PUGB7
			10'd147 : rdata = 48'b110001110000001000000000000000000000000000001111;
			// PEs: 41 -> 56
			// srcs: (158, 205)(2967) 5 --> (2967) 5:PEGB1, pass, PUGB7
			10'd148 : rdata = 48'b110001110000001000000000000000000000000000001111;
			// PEs: 47 -> 48
			// srcs: (159, 126)(2115) 3 --> (2115) 3:PENB, pass, PUNB
			10'd149 : rdata = 48'b110001101111111000000000000000000000001000000000;
			// PEs: 43 -> 32
			// srcs: (162, 215)(2298) 0 --> (2298) 0:PEGB3, pass, PUGB4
			10'd150 : rdata = 48'b110001110000011000000000000000000000000000001100;
			// PEs: 41 -> 32
			// srcs: (163, 223)(3125) -2 --> (3125) -2:PEGB1, pass, PUGB4
			10'd151 : rdata = 48'b110001110000001000000000000000000000000000001100;
			// PEs: 42 -> 48
			// srcs: (167, 136)(2473) -6 --> (2473) -6:PEGB2, pass, PUNB
			10'd152 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 45 -> 48
			// srcs: (175, 149)(1756) -2 --> (1756) -2:PEGB5, pass, PUNB
			10'd153 : rdata = 48'b110001110000101000000000000000000000001000000000;
			// PEs: 45 -> 48
			// srcs: (183, 152)(2555) 1 --> (2555) 1:PEGB5, pass, PUNB
			10'd154 : rdata = 48'b110001110000101000000000000000000000001000000000;
			// PEs: 46 -> 48
			// srcs: (191, 153)(2558) 11 --> (2558) 11:PEGB6, pass, PUNB
			10'd155 : rdata = 48'b110001110000110000000000000000000000001000000000;
			// PEs: 47 -> 48
			// srcs: (196, 154)(2560) -6 --> (2560) -6:PENB, pass, PUNB
			10'd156 : rdata = 48'b110001101111111000000000000000000000001000000000;
			// PEs: 43 -> 48
			// srcs: (204, 162)(2637) -2 --> (2637) -2:PEGB3, pass, PUNB
			10'd157 : rdata = 48'b110001110000011000000000000000000000001000000000;
			// PEs: 41 -> 48
			// srcs: (212, 164)(2657) -2 --> (2657) -2:PEGB1, pass, PUNB
			10'd158 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 46 -> 48
			// srcs: (220, 183)(2804) 0 --> (2804) 0:PEGB6, pass, PUNB
			10'd159 : rdata = 48'b110001110000110000000000000000000000001000000000;
			// PEs: 32 -> 40
			// srcs: (221, 120)(2016) 1 --> (2016) 1:PUNB, pass, NI0
			10'd160 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 42 -> 48
			// srcs: (229, 187)(2111) 0 --> (2111) 0:PEGB2, pass, PUNB
			10'd161 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 32 -> 41
			// srcs: (237, 121)(2017) 0 --> (2017) 0:PUNB, pass, PENB
			10'd162 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 41 -> 48
			// srcs: (238, 202)(2957) 3 --> (2957) 3:PEGB1, pass, PUNB
			10'd163 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 40 -> 41
			// srcs: (243, 122)(2016) 1 --> (2016) 1:NI0, pass, PENB
			10'd164 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 16 -> 40
			// srcs: (244, 129)(2411) 0 --> (2411) 0:PUGB2, pass, NI0
			10'd165 : rdata = 48'b110001110000010100000000000100000000000000000000;
			// PEs: 0 -> 41
			// srcs: (245, 130)(1631) 0 --> (1631) 0:PUGB0, pass, PENB
			10'd166 : rdata = 48'b110001110000000100000000000000000000000100000000;
			// PEs: 41 -> 48
			// srcs: (246, 209)(3046) 1 --> (3046) 1:PEGB1, pass, PUNB
			10'd167 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 40 -> 41
			// srcs: (251, 131)(2411) 0 --> (2411) 0:NI0, pass, PENB
			10'd168 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 24 -> 40
			// srcs: (252, 132)(2436) 1 --> (2436) 1:PUGB3, pass, NI0
			10'd169 : rdata = 48'b110001110000011100000000000100000000000000000000;
			// PEs: 8 -> 41
			// srcs: (253, 133)(1658) 4 --> (1658) 4:PUGB1, pass, PENB
			10'd170 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 41 -> 48
			// srcs: (254, 213)(2292) -2 --> (2292) -2:PEGB1, pass, PUNB
			10'd171 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 40 -> 41
			// srcs: (259, 134)(2436) 1 --> (2436) 1:NI0, pass, PENB
			10'd172 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 24 -> 41
			// srcs: (260, 138)(1701) -1 --> (1701) -1:PUGB3, pass, PENB
			10'd173 : rdata = 48'b110001110000011100000000000000000000000100000000;
			// PEs: 48 -> 40
			// srcs: (261, 139)(2489) 0 --> (2489) 0:PUGB6, pass, NI0
			10'd174 : rdata = 48'b110001110000110100000000000100000000000000000000;
			// PEs: 24 -> 41
			// srcs: (262, 140)(1710) 2 --> (1710) 2:PUGB3, pass, PENB
			10'd175 : rdata = 48'b110001110000011100000000000000000000000100000000;
			// PEs: 46 -> 48
			// srcs: (263, 218)(2307) 2 --> (2307) 2:PEGB6, pass, PUNB
			10'd176 : rdata = 48'b110001110000110000000000000000000000001000000000;
			// PEs: 41 -> 48
			// srcs: (264, 229)(2412) 0 --> (2412) 0:PEGB1, pass, PUNB
			10'd177 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 41 -> 32
			// srcs: (266, 230)(2437) 5 --> (2437) 5:PEGB1, pass, PUGB4
			10'd178 : rdata = 48'b110001110000001000000000000000000000000000001100;
			// PEs: 40 -> 41
			// srcs: (268, 141)(2489) 0 --> (2489) 0:NI0, pass, PENB
			10'd179 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 8 -> 40
			// srcs: (269, 142)(2516) -2 --> (2516) -2:PUGB1, pass, NI0
			10'd180 : rdata = 48'b110001110000001100000000000100000000000000000000;
			// PEs: 32 -> 41
			// srcs: (270, 143)(1738) 0 --> (1738) 0:PUNB, pass, PENB
			10'd181 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 41 -> 24
			// srcs: (275, 235)(2490) 2 --> (2490) 2:PEGB1, pass, PUGB3
			10'd182 : rdata = 48'b110001110000001000000000000000000000000000001011;
			// PEs: 40 -> 41
			// srcs: (276, 144)(2516) -2 --> (2516) -2:NI0, pass, PENB
			10'd183 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 24 -> 40
			// srcs: (277, 155)(2571) 0 --> (2571) 0:PUGB3, pass, NI0
			10'd184 : rdata = 48'b110001110000011100000000000100000000000000000000;
			// PEs: 56 -> 41
			// srcs: (278, 156)(1793) -1 --> (1793) -1:PUGB7, pass, PENB
			10'd185 : rdata = 48'b110001110000111100000000000000000000000100000000;
			// PEs: 40 -> 41
			// srcs: (284, 157)(2571) 0 --> (2571) 0:NI0, pass, PENB
			10'd186 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 24 -> 40
			// srcs: (285, 158)(2614) -2 --> (2614) -2:PUGB3, pass, NI0
			10'd187 : rdata = 48'b110001110000011100000000000100000000000000000000;
			// PEs: 8 -> 41
			// srcs: (286, 159)(1836) 6 --> (1836) 6:PUGB1, pass, PENB
			10'd188 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 41 -> 56
			// srcs: (291, 240)(2572) -1 --> (2572) -1:PEGB1, pass, PUGB7
			10'd189 : rdata = 48'b110001110000001000000000000000000000000000001111;
			// PEs: 40 -> 41
			// srcs: (292, 160)(2614) -2 --> (2614) -2:NI0, pass, PENB
			10'd190 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 41 -> 56
			// srcs: (299, 241)(2615) 4 --> (2615) 4:PEGB1, pass, PUGB7
			10'd191 : rdata = 48'b110001110000001000000000000000000000000000001111;
			// PEs: 16 -> 41
			// srcs: (369, 161)(1857) -2 --> (1857) -2:PUGB2, pass, PENB
			10'd192 : rdata = 48'b110001110000010100000000000000000000000100000000;
			// PEs: 48 -> 40
			// srcs: (370, 165)(2666) -8 --> (2666) -8:PUGB6, pass, NI0
			10'd193 : rdata = 48'b110001110000110100000000000100000000000000000000;
			// PEs: 24 -> 41
			// srcs: (371, 166)(1888) -2 --> (1888) -2:PUGB3, pass, PENB
			10'd194 : rdata = 48'b110001110000011100000000000000000000000100000000;
			// PEs: 41 -> 48
			// srcs: (376, 242)(2636) 2 --> (2636) 2:PEGB1, pass, PUNB
			10'd195 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 40 -> 41
			// srcs: (377, 167)(2666) -8 --> (2666) -8:NI0, pass, PENB
			10'd196 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 16 -> 40
			// srcs: (378, 168)(2689) -2 --> (2689) -2:PUGB2, pass, NI0
			10'd197 : rdata = 48'b110001110000010100000000000100000000000000000000;
			// PEs: 32 -> 41
			// srcs: (379, 169)(1912) 3 --> (1912) 3:PUNB, pass, PENB
			10'd198 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 41 -> 48
			// srcs: (384, 246)(2667) -10 --> (2667) -10:PEGB1, pass, PUNB
			10'd199 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 40 -> 41
			// srcs: (385, 170)(2689) -2 --> (2689) -2:NI0, pass, PENB
			10'd200 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 32 -> 41
			// srcs: (386, 171)(2705) -4 --> (2705) -4:PUNB, pass, PENB
			10'd201 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 32 -> 41
			// srcs: (387, 172)(2709) -1 --> (2709) -1:PUNB, pass, PENB
			10'd202 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 32 -> 41
			// srcs: (388, 173)(2711) -4 --> (2711) -4:PUNB, pass, PENB
			10'd203 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 32 -> 40
			// srcs: (389, 174)(2788) -3 --> (2788) -3:PUNB, pass, NI0
			10'd204 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 0 -> 41
			// srcs: (390, 175)(2010) -2 --> (2010) -2:PUGB0, pass, PENB
			10'd205 : rdata = 48'b110001110000000100000000000000000000000100000000;
			// PEs: 41 -> 48
			// srcs: (392, 247)(2690) 1 --> (2690) 1:PEGB1, pass, PUNB
			10'd206 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 42 -> 48
			// srcs: (400, 254)(2886) -9 --> (2886) -9:PEGB2, pass, PUNB
			10'd207 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 40 -> 41
			// srcs: (401, 176)(2788) -3 --> (2788) -3:NI0, pass, PENB
			10'd208 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 32 -> 40
			// srcs: (402, 177)(2790) -10 --> (2790) -10:PUNB, pass, NI0
			10'd209 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 0 -> 41
			// srcs: (403, 178)(2013) 2 --> (2013) 2:PUGB0, pass, PENB
			10'd210 : rdata = 48'b110001110000000100000000000000000000000100000000;
			// PEs: 40 -> 41
			// srcs: (409, 179)(2790) -10 --> (2790) -10:NI0, pass, PENB
			10'd211 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 32 -> 41
			// srcs: (410, 180)(2796) 4 --> (2796) 4:PUNB, pass, PENB
			10'd212 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 41 -> 16
			// srcs: (417, 249)(2798) 5 --> (2798) 5:PEGB1, pass, PUGB2
			10'd213 : rdata = 48'b110001110000001000000000000000000000000000001010;
			// PEs: 42 -> 32
			// srcs: (425, 279)(2792) -13 --> (2792) -13:PEGB2, pass, PUGB4
			10'd214 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 32 -> 44
			// srcs: (607, 184)(2099) 0 --> (2099) 0:PUNB, pass, PEGB4
			10'd215 : rdata = 48'b110001101111111100000000000000000000000011000000;
			// PEs: 32 -> 47
			// srcs: (608, 185)(2102) 0 --> (2102) 0:PUNB, pass, PEGB7
			10'd216 : rdata = 48'b110001101111111100000000000000000000000011110000;
			// PEs: 32 -> 41
			// srcs: (625, 186)(2105) -1 --> (2105) -1:PUNB, pass, PENB
			10'd217 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 8 -> 40
			// srcs: (626, 193)(2919) 0 --> (2919) 0:PUGB1, pass, NI0
			10'd218 : rdata = 48'b110001110000001100000000000100000000000000000000;
			// PEs: 48 -> 41
			// srcs: (627, 194)(2142) -2 --> (2142) -2:PUGB6, pass, PENB
			10'd219 : rdata = 48'b110001110000110100000000000000000000000100000000;
			// PEs: 40 -> 41
			// srcs: (633, 195)(2919) 0 --> (2919) 0:NI0, pass, PENB
			10'd220 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 16 -> 40
			// srcs: (634, 196)(2933) 4 --> (2933) 4:PUGB2, pass, NI0
			10'd221 : rdata = 48'b110001110000010100000000000100000000000000000000;
			// PEs: 56 -> 41
			// srcs: (635, 197)(2157) 4 --> (2157) 4:PUGB7, pass, PENB
			10'd222 : rdata = 48'b110001110000111100000000000000000000000100000000;
			// PEs: 41 -> 48
			// srcs: (640, 255)(2920) -2 --> (2920) -2:PEGB1, pass, PUNB
			10'd223 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 40 -> 41
			// srcs: (641, 198)(2933) 4 --> (2933) 4:NI0, pass, PENB
			10'd224 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 32 -> 40
			// srcs: (642, 199)(2949) -2 --> (2949) -2:PUNB, pass, NI0
			10'd225 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 56 -> 41
			// srcs: (643, 200)(2170) -6 --> (2170) -6:PUGB7, pass, PENB
			10'd226 : rdata = 48'b110001110000111100000000000000000000000100000000;
			// PEs: 41 -> 48
			// srcs: (648, 256)(2934) 8 --> (2934) 8:PEGB1, pass, PUNB
			10'd227 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 40 -> 41
			// srcs: (649, 201)(2949) -2 --> (2949) -2:NI0, pass, PENB
			10'd228 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 56 -> 40
			// srcs: (650, 206)(2980) 4 --> (2980) 4:PUGB7, pass, NI0
			10'd229 : rdata = 48'b110001110000111100000000000100000000000000000000;
			// PEs: 8 -> 41
			// srcs: (651, 207)(2203) 1 --> (2203) 1:PUGB1, pass, PENB
			10'd230 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 41 -> 0
			// srcs: (656, 257)(2950) -8 --> (2950) -8:PEGB1, pass, PUGB0
			10'd231 : rdata = 48'b110001110000001000000000000000000000000000001000;
			// PEs: 40 -> 41
			// srcs: (657, 208)(2980) 4 --> (2980) 4:NI0, pass, PENB
			10'd232 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 32 -> 41
			// srcs: (658, 210)(2271) 4 --> (2271) 4:PUNB, pass, PENB
			10'd233 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 41 -> 48
			// srcs: (672, 259)(3049) -2 --> (3049) -2:PEGB1, pass, PUNB
			10'd234 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 32 -> 41
			// srcs: (674, 211)(2274) 4 --> (2274) 4:PUNB, pass, PENB
			10'd235 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 32 -> 41
			// srcs: (692, 212)(2277) 0 --> (2277) 0:PUNB, pass, PENB
			10'd236 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 32 -> 40
			// srcs: (693, 220)(3117) -1 --> (3117) -1:PUNB, pass, NI0
			10'd237 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 56 -> 41
			// srcs: (694, 221)(2341) -4 --> (2341) -4:PUGB7, pass, PENB
			10'd238 : rdata = 48'b110001110000111100000000000000000000000100000000;
			// PEs: 40 -> 41
			// srcs: (705, 222)(3117) -1 --> (3117) -1:NI0, pass, PENB
			10'd239 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 56 -> 41
			// srcs: (706, 225)(2356) 0 --> (2356) 0:PUGB7, pass, PENB
			10'd240 : rdata = 48'b110001110000111100000000000000000000000100000000;
			// PEs: 16 -> 40
			// srcs: (707, 226)(2398) -10 --> (2398) -10:PUGB2, pass, NI0
			10'd241 : rdata = 48'b110001110000010100000000000100000000000000000000;
			// PEs: 48 -> 41
			// srcs: (708, 227)(2400) 2 --> (2400) 2:PUGB6, pass, PENB
			10'd242 : rdata = 48'b110001110000110100000000000000000000000100000000;
			// PEs: 41 -> 8
			// srcs: (712, 263)(3118) -5 --> (3118) -5:PEGB1, pass, PUGB1
			10'd243 : rdata = 48'b110001110000001000000000000000000000000000001001;
			// PEs: 41 -> 24
			// srcs: (713, 264)(3131) -2 --> (3131) -2:PEGB1, pass, PUGB3
			10'd244 : rdata = 48'b110001110000001000000000000000000000000000001011;
			// PEs: 40 -> 41
			// srcs: (714, 228)(2398) -10 --> (2398) -10:NI0, pass, PENB
			10'd245 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 48 -> 40
			// srcs: (715, 231)(2441) 2 --> (2441) 2:PUGB6, pass, NI0
			10'd246 : rdata = 48'b110001110000110100000000000100000000000000000000;
			// PEs: 8 -> 41
			// srcs: (716, 232)(2443) 0 --> (2443) 0:PUGB1, pass, PENB
			10'd247 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 42 -> 24
			// srcs: (717, 287)(3056) -4 --> (3056) -4:PEGB2, pass, PUGB3
			10'd248 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 41 -> 16
			// srcs: (721, 268)(2401) -8 --> (2401) -8:PEGB1, pass, PUGB2
			10'd249 : rdata = 48'b110001110000001000000000000000000000000000001010;
			// PEs: 40 -> 41
			// srcs: (722, 233)(2441) 2 --> (2441) 2:NI0, pass, PENB
			10'd250 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 32 -> 41
			// srcs: (723, 234)(2479) 0 --> (2479) 0:PUNB, pass, PENB
			10'd251 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 32 -> 41
			// srcs: (724, 236)(2515) 1 --> (2515) 1:PUNB, pass, PENB
			10'd252 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 32 -> 40
			// srcs: (725, 237)(2543) 0 --> (2543) 0:PUNB, pass, NI0
			10'd253 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 48 -> 41
			// srcs: (726, 238)(2545) -5 --> (2545) -5:PUGB6, pass, PENB
			10'd254 : rdata = 48'b110001110000110100000000000000000000000100000000;
			// PEs: 32 -> 46
			// srcs: (727, 248)(2704) -6 --> (2704) -6:PUNB, pass, PEGB6
			10'd255 : rdata = 48'b110001101111111100000000000000000000000011100000;
			// PEs: 41 -> 8
			// srcs: (729, 269)(2444) 2 --> (2444) 2:PEGB1, pass, PUGB1
			10'd256 : rdata = 48'b110001110000001000000000000000000000000000001001;
			// PEs: 40 -> 41
			// srcs: (732, 239)(2543) 0 --> (2543) 0:NI0, pass, PENB
			10'd257 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 24 -> 40
			// srcs: (733, 243)(2641) 7 --> (2641) 7:PUGB3, pass, NI0
			10'd258 : rdata = 48'b110001110000011100000000000100000000000000000000;
			// PEs: 56 -> 41
			// srcs: (734, 244)(2643) -5 --> (2643) -5:PUGB7, pass, PENB
			10'd259 : rdata = 48'b110001110000111100000000000000000000000100000000;
			// PEs: 41 -> 48
			// srcs: (739, 272)(2546) -5 --> (2546) -5:PEGB1, pass, PUNB
			10'd260 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 40 -> 41
			// srcs: (740, 245)(2641) 7 --> (2641) 7:NI0, pass, PENB
			10'd261 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 0 -> 40
			// srcs: (741, 250)(2809) -6 --> (2809) -6:PUGB0, pass, NI0
			10'd262 : rdata = 48'b110001110000000100000000000100000000000000000000;
			// PEs: 16 -> 41
			// srcs: (742, 251)(2811) -3 --> (2811) -3:PUGB2, pass, PENB
			10'd263 : rdata = 48'b110001110000010100000000000000000000000100000000;
			// PEs: 41 -> 48
			// srcs: (747, 273)(2644) 2 --> (2644) 2:PEGB1, pass, PUNB
			10'd264 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 40 -> 41
			// srcs: (748, 252)(2809) -6 --> (2809) -6:NI0, pass, PENB
			10'd265 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 32 -> 41
			// srcs: (749, 253)(2875) 8 --> (2875) 8:PUNB, pass, PENB
			10'd266 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 8 -> 41
			// srcs: (750, 258)(2979) -7 --> (2979) -7:PUGB1, pass, PENB
			10'd267 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 24 -> 40
			// srcs: (751, 260)(3081) 1 --> (3081) 1:PUGB3, pass, NI0
			10'd268 : rdata = 48'b110001110000011100000000000100000000000000000000;
			// PEs: 48 -> 41
			// srcs: (752, 261)(3083) -2 --> (3083) -2:PUGB6, pass, PENB
			10'd269 : rdata = 48'b110001110000110100000000000000000000000100000000;
			// PEs: 47 -> 48
			// srcs: (757, 278)(2725) 4 --> (2725) 4:PENB, pass, PUNB
			10'd270 : rdata = 48'b110001101111111000000000000000000000001000000000;
			// PEs: 41 -> 48
			// srcs: (758, 280)(2812) -9 --> (2812) -9:PEGB1, pass, PUNB
			10'd271 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 43 -> 48
			// srcs: (759, 285)(2884) 2 --> (2884) 2:PEGB3, pass, PUNB
			10'd272 : rdata = 48'b110001110000011000000000000000000000001000000000;
			// PEs: 40 -> 41
			// srcs: (763, 262)(3081) 1 --> (3081) 1:NI0, pass, PENB
			10'd273 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 16 -> 40
			// srcs: (764, 265)(2362) -7 --> (2362) -7:PUGB2, pass, NI0
			10'd274 : rdata = 48'b110001110000010100000000000100000000000000000000;
			// PEs: 48 -> 41
			// srcs: (765, 266)(2367) -22 --> (2367) -22:PUGB6, pass, PENB
			10'd275 : rdata = 48'b110001110000110100000000000000000000000100000000;
			// PEs: 41 -> 0
			// srcs: (766, 286)(2982) -2 --> (2982) -2:PEGB1, pass, PUGB0
			10'd276 : rdata = 48'b110001110000001000000000000000000000000000001000;
			// PEs: 40 -> 41
			// srcs: (771, 267)(2362) -7 --> (2362) -7:NI0, pass, PENB
			10'd277 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 8 -> 41
			// srcs: (772, 270)(2487) 14 --> (2487) 14:PUGB1, pass, PENB
			10'd278 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 0 -> 41
			// srcs: (773, 271)(2523) 4 --> (2523) 4:PUGB0, pass, PENB
			10'd279 : rdata = 48'b110001110000000100000000000000000000000100000000;
			// PEs: 16 -> 40
			// srcs: (774, 274)(2654) 10 --> (2654) 10:PUGB2, pass, NI0
			10'd280 : rdata = 48'b110001110000010100000000000100000000000000000000;
			// PEs: 32 -> 41
			// srcs: (775, 275)(2659) -2 --> (2659) -2:PUNB, pass, PENB
			10'd281 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 32 -> 45
			// srcs: (776, 277)(2702) 13 --> (2702) 13:PUNB, pass, PEGB5
			10'd282 : rdata = 48'b110001101111111100000000000000000000000011010000;
			// PEs: 41 -> 16
			// srcs: (778, 289)(2368) -29 --> (2368) -29:PEGB1, pass, PUGB2
			10'd283 : rdata = 48'b110001110000001000000000000000000000000000001010;
			// PEs: 41 -> 0
			// srcs: (779, 293)(2488) 11 --> (2488) 11:PEGB1, pass, PUGB0
			10'd284 : rdata = 48'b110001110000001000000000000000000000000000001000;
			// PEs: 41 -> 24
			// srcs: (780, 294)(2524) 3 --> (2524) 3:PEGB1, pass, PUGB3
			10'd285 : rdata = 48'b110001110000001000000000000000000000000000001011;
			// PEs: 40 -> 41
			// srcs: (781, 276)(2654) 10 --> (2654) 10:NI0, pass, PENB
			10'd286 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 32 -> 40
			// srcs: (782, 281)(2824) 10 --> (2824) 10:PUNB, pass, NI0
			10'd287 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 56 -> 41
			// srcs: (783, 282)(2829) -9 --> (2829) -9:PUGB7, pass, PENB
			10'd288 : rdata = 48'b110001110000111100000000000000000000000100000000;
			// PEs: 40 -> 41
			// srcs: (789, 283)(2824) 10 --> (2824) 10:NI0, pass, PENB
			10'd289 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 46 -> 56
			// srcs: (791, 307)(2720) -2 --> (2720) -2:PEGB6, pass, PUGB7
			10'd290 : rdata = 48'b110001110000110000000000000000000000000000001111;
			// PEs: 41 -> 24
			// srcs: (796, 296)(2830) 1 --> (2830) 1:PEGB1, pass, PUGB3
			10'd291 : rdata = 48'b110001110000001000000000000000000000000000001011;
			// PEs: 32 -> 41
			// srcs: (1115, 284)(2873) -2 --> (2873) -2:PUNB, pass, PENB
			10'd292 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 24 -> 41
			// srcs: (1116, 288)(3079) 2 --> (3079) 2:PUGB3, pass, PENB
			10'd293 : rdata = 48'b110001110000011100000000000000000000000100000000;
			// PEs: 32 -> 40
			// srcs: (1117, 290)(2416) 3 --> (2416) 3:PUNB, pass, NI0
			10'd294 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 56 -> 41
			// srcs: (1118, 291)(2427) -7 --> (2427) -7:PUGB7, pass, PENB
			10'd295 : rdata = 48'b110001110000111100000000000000000000000100000000;
			// PEs: 41 -> 48
			// srcs: (1122, 300)(2879) 12 --> (2879) 12:PEGB1, pass, PUNB
			10'd296 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 40 -> 41
			// srcs: (1125, 292)(2416) 3 --> (2416) 3:NI0, pass, PENB
			10'd297 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 0 -> 41
			// srcs: (1126, 295)(2671) -14 --> (2671) -14:PUGB0, pass, PENB
			10'd298 : rdata = 48'b110001110000000100000000000000000000000100000000;
			// PEs: 0 -> 40
			// srcs: (1127, 297)(2856) 9 --> (2856) 9:PUGB0, pass, NI0
			10'd299 : rdata = 48'b110001110000000100000000000100000000000000000000;
			// PEs: 32 -> 41
			// srcs: (1128, 298)(2867) 2 --> (2867) 2:PUNB, pass, PENB
			10'd300 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 41 -> 48
			// srcs: (1132, 302)(2428) -4 --> (2428) -4:PEGB1, pass, PUNB
			10'd301 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 41 -> 48
			// srcs: (1133, 306)(2672) -6 --> (2672) -6:PEGB1, pass, PUNB
			10'd302 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 40 -> 41
			// srcs: (1136, 299)(2856) 9 --> (2856) 9:NI0, pass, PENB
			10'd303 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 32 -> 41
			// srcs: (1137, 301)(3074) -1 --> (3074) -1:PUNB, pass, PENB
			10'd304 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 41 -> 48
			// srcs: (1143, 308)(2868) 11 --> (2868) 11:PEGB1, pass, PUNB
			10'd305 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 41 -> 0
			// srcs: (1144, 309)(3086) 0 --> (3086) 0:PEGB1, pass, PUGB0
			10'd306 : rdata = 48'b110001110000001000000000000000000000000000001000;
			// PEs: 16 -> 40
			// srcs: (1177, 303)(2623) 27 --> (2623) 27:PUGB2, pass, NI0
			10'd307 : rdata = 48'b110001110000010100000000000100000000000000000000;
			// PEs: 32 -> 41
			// srcs: (1178, 304)(2646) 21 --> (2646) 21:PUNB, pass, PENB
			10'd308 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 40 -> 41
			// srcs: (1184, 305)(2623) 27 --> (2623) 27:NI0, pass, PENB
			10'd309 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 0 -> 40
			// srcs: (1186, 310)(2501) 26 --> (2501) 26:PUGB0, pass, NI0
			10'd310 : rdata = 48'b110001110000000100000000000100000000000000000000;
			// PEs: 32 -> 41
			// srcs: (1187, 311)(2549) -2 --> (2549) -2:PUNB, pass, PENB
			10'd311 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 41 -> 48
			// srcs: (1191, 313)(2647) 48 --> (2647) 48:PEGB1, pass, PUNB
			10'd312 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 40 -> 41
			// srcs: (1193, 312)(2501) 26 --> (2501) 26:NI0, pass, PENB
			10'd313 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 41 -> 0
			// srcs: (1200, 314)(2550) 24 --> (2550) 24:PEGB1, pass, PUGB0
			10'd314 : rdata = 48'b110001110000001000000000000000000000000000001000;
			// PEs: 32 -> 40
			// srcs: (1444, 315)(3039) -38 --> (3039) -38:PUNB, pass, NI0
			10'd315 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 8 -> 41
			// srcs: (1447, 316)(3136) -25 --> (3136) -25:PUGB1, pass, PENB
			10'd316 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 40 -> 41
			// srcs: (1454, 317)(3039) -38 --> (3039) -38:NI0, pass, PENB
			10'd317 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 41 -> 48
			// srcs: (1461, 318)(3137) -63 --> (3137) -63:PEGB1, pass, PUNB
			10'd318 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 8 -> 46
			// srcs: (1516, 319)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd319 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 47
			// srcs: (1519, 320)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd320 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 41
			// srcs: (1559, 321)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd321 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 42
			// srcs: (1560, 322)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd322 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 43
			// srcs: (1561, 323)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd323 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 44
			// srcs: (1562, 324)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd324 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 45
			// srcs: (1563, 325)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd325 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 46
			// srcs: (1565, 326)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd326 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 47
			// srcs: (1566, 327)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd327 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 41
			// srcs: (1639, 328)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd328 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 42
			// srcs: (1641, 329)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd329 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 43
			// srcs: (1642, 330)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd330 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 44
			// srcs: (1644, 331)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd331 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 45
			// srcs: (1645, 332)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd332 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 46
			// srcs: (1647, 333)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd333 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 47
			// srcs: (1648, 334)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd334 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 41
			// srcs: (1680, 335)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd335 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 42
			// srcs: (1683, 336)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd336 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 43
			// srcs: (1686, 337)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd337 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 44
			// srcs: (1689, 338)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd338 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 45
			// srcs: (1692, 339)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd339 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 46
			// srcs: (1695, 340)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd340 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 47
			// srcs: (1698, 341)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd341 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 41
			// srcs: (1719, 342)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd342 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 42
			// srcs: (1721, 343)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd343 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 43
			// srcs: (1722, 344)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd344 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 44
			// srcs: (1724, 345)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd345 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 45
			// srcs: (1725, 346)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd346 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 46
			// srcs: (1727, 347)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd347 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 47
			// srcs: (1728, 348)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd348 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 41
			// srcs: (1801, 349)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd349 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 42
			// srcs: (1803, 350)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd350 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 43
			// srcs: (1804, 351)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd351 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 44
			// srcs: (1805, 352)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd352 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 45
			// srcs: (1806, 353)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd353 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 46
			// srcs: (1807, 354)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd354 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 47
			// srcs: (1808, 355)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd355 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 41
			// srcs: (1864, 356)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd356 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 42
			// srcs: (1867, 357)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd357 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 43
			// srcs: (1870, 358)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd358 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 44
			// srcs: (1873, 359)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd359 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 45
			// srcs: (1876, 360)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd360 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 46
			// srcs: (1879, 361)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd361 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 41
			// srcs: (1881, 362)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd362 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 47
			// srcs: (1882, 363)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd363 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 42
			// srcs: (1883, 364)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd364 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 43
			// srcs: (1884, 365)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd365 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 44
			// srcs: (1886, 366)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd366 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 45
			// srcs: (1887, 367)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd367 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 46
			// srcs: (1889, 368)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd368 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 47
			// srcs: (1890, 369)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd369 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 41
			// srcs: (1961, 370)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd370 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 42
			// srcs: (1963, 371)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd371 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 43
			// srcs: (1964, 372)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd372 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 44
			// srcs: (1966, 373)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd373 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 45
			// srcs: (1967, 374)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd374 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 46
			// srcs: (1969, 375)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd375 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 47
			// srcs: (1970, 376)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd376 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 41
			// srcs: (2043, 377)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd377 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 41
			// srcs: (2044, 378)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd378 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 42
			// srcs: (2045, 379)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd379 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 43
			// srcs: (2046, 380)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd380 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 42
			// srcs: (2047, 381)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd381 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 44
			// srcs: (2048, 382)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd382 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 45
			// srcs: (2049, 383)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd383 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 46
			// srcs: (2050, 384)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd384 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 47
			// srcs: (2051, 385)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd385 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 43
			// srcs: (2054, 386)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd386 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 44
			// srcs: (2057, 387)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd387 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 45
			// srcs: (2060, 388)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd388 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 46
			// srcs: (2063, 389)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd389 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 47
			// srcs: (2066, 390)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd390 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 41
			// srcs: (2123, 391)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd391 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 42
			// srcs: (2125, 392)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd392 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 43
			// srcs: (2126, 393)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd393 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 44
			// srcs: (2128, 394)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd394 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 45
			// srcs: (2129, 395)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd395 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 46
			// srcs: (2131, 396)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd396 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 47
			// srcs: (2132, 397)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd397 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 41
			// srcs: (2203, 398)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd398 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 42
			// srcs: (2205, 399)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd399 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 43
			// srcs: (2206, 400)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd400 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 44
			// srcs: (2208, 401)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd401 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 45
			// srcs: (2209, 402)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd402 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 46
			// srcs: (2211, 403)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd403 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 47
			// srcs: (2212, 404)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd404 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 41
			// srcs: (2228, 405)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd405 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 42
			// srcs: (2231, 406)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd406 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 43
			// srcs: (2234, 407)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd407 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 44
			// srcs: (2237, 408)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd408 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 45
			// srcs: (2240, 409)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd409 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 46
			// srcs: (2243, 410)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd410 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 47
			// srcs: (2250, 411)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd411 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 41
			// srcs: (2285, 412)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd412 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 42
			// srcs: (2287, 413)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd413 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 43
			// srcs: (2288, 414)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd414 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 44
			// srcs: (2290, 415)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd415 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 45
			// srcs: (2291, 416)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd416 : rdata = 48'b110001110000001100000000000000000000000011010000;
			default : rdata = 48'b000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 41) begin
	always @(*) begin
		case(address)
			// PEs: 41, 41 -> 41
			// srcs: (1, 0)(54) 0, (839) -2 --> (1623) 0:ND0, NW0, *, NI0
			10'd0 : rdata = 48'b000110110000000001000000000100000000000000000000;
			// PEs: 41, 41 -> 40
			// srcs: (2, 1)(134) -3, (919) -1 --> (1703) 3:ND1, NW1, *, PEGB0
			10'd1 : rdata = 48'b000110110000000101000000001000000000000010000000;
			// PEs: 41, 41 -> 40
			// srcs: (3, 2)(214) 1, (999) 2 --> (1783) 2:ND2, NW2, *, PEGB0
			10'd2 : rdata = 48'b000110110000001001000000010000000000000010000000;
			// PEs: 41, 41 -> 40
			// srcs: (4, 3)(296) 1, (1081) -3 --> (1865) -3:ND3, NW3, *, PEGB0
			10'd3 : rdata = 48'b000110110000001101000000011000000000000010000000;
			// PEs: 41, 41 -> 45
			// srcs: (5, 4)(376) -2, (1161) 1 --> (1945) -2:ND4, NW4, *, PEGB5
			10'd4 : rdata = 48'b000110110000010001000000100000000000000011010000;
			// PEs: 41, 41 -> 46
			// srcs: (6, 5)(456) 0, (1241) -1 --> (2025) 0:ND5, NW5, *, PEGB6
			10'd5 : rdata = 48'b000110110000010101000000101000000000000011100000;
			// PEs: 41, 41 -> 47
			// srcs: (7, 6)(538) -3, (1323) -1 --> (2107) 3:ND6, NW6, *, PEGB7
			10'd6 : rdata = 48'b000110110000011001000000110000000000000011110000;
			// PEs: 41, 41 -> 41
			// srcs: (8, 7)(618) 1, (1403) 2 --> (2187) 2:ND7, NW7, *, NI1
			10'd7 : rdata = 48'b000110110000011101000000111100001000000000000000;
			// PEs: 41, 41 -> 41
			// srcs: (9, 8)(698) 2, (1483) 2 --> (2267) 4:ND8, NW8, *, NI2
			10'd8 : rdata = 48'b000110110000100001000001000100010000000000000000;
			// PEs: 41, 41 -> 41
			// srcs: (10, 9)(780) 0, (1565) -1 --> (2349) 0:ND9, NW9, *, NI3
			10'd9 : rdata = 48'b000110110000100101000001001100011000000000000000;
			// PEs: 41, 41 -> 41
			// srcs: (11, 10)(175) 1, (960) 1 --> (1744) 1:ND10, NW10, *, NI4
			10'd10 : rdata = 48'b000110110000101001000001010100100000000000000000;
			// PEs: 41, 41 -> 41
			// srcs: (12, 11)(359) 1, (1144) -1 --> (1928) -1:ND11, NW11, *, NI5
			10'd11 : rdata = 48'b000110110000101101000001011100101000000000000000;
			// PEs: 41, 41 -> 42
			// srcs: (13, 12)(539) -3, (1324) 2 --> (2108) -6:ND12, NW12, *, PENB
			10'd12 : rdata = 48'b000110110000110001000001100000000000000100000000;
			// PEs: 41, 41 -> 41
			// srcs: (14, 13)(723) -2, (1508) 1 --> (2292) -2:ND13, NW13, *, NI6
			10'd13 : rdata = 48'b000110110000110101000001101100110000000000000000;
			// PEs: 40 -> 
			// srcs: (39, 14)(1666) 0 --> (1666) 0:PENB, pass, 
			10'd14 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 40, 41 -> 41
			// srcs: (45, 15)(1665) -1, (1666) 0 --> (2445) -1:PENB, ALU, +, NI7
			10'd15 : rdata = 48'b000011101111111000111111111100111000000000000000;
			// PEs: 40 -> 
			// srcs: (58, 16)(1878) -2 --> (1878) -2:PENB, pass, 
			10'd16 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 40, 41 -> 41
			// srcs: (64, 17)(1877) 0, (1878) -2 --> (2657) -2:PENB, ALU, +, NI8
			10'd17 : rdata = 48'b000011101111111000111111111101000000000000000000;
			// PEs: 40 -> 
			// srcs: (66, 18)(1936) -3 --> (1936) -3:PENB, pass, 
			10'd18 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 40, 41 -> 47
			// srcs: (72, 19)(1935) 4, (1936) -3 --> (2714) 1:PENB, ALU, +, PEGB7
			10'd19 : rdata = 48'b000011101111111000111111111000000000000011110000;
			// PEs: 40 -> 
			// srcs: (74, 20)(1939) -1 --> (1939) -1:PENB, pass, 
			10'd20 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 40, 41 -> 46
			// srcs: (80, 21)(1938) -2, (1939) -1 --> (2716) -3:PENB, ALU, +, PEGB6
			10'd21 : rdata = 48'b000011101111111000111111111000000000000011100000;
			// PEs: 40 -> 
			// srcs: (82, 22)(1942) 2 --> (1942) 2:PENB, pass, 
			10'd22 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 40, 41 -> 46
			// srcs: (88, 23)(1941) 0, (1942) 2 --> (2721) 2:PENB, ALU, +, PEGB6
			10'd23 : rdata = 48'b000011101111111000111111111000000000000011100000;
			// PEs: 40 -> 41
			// srcs: (90, 24)(2019) 0 --> (2019) 0:PENB, pass, NI9
			10'd24 : rdata = 48'b110001101111111000000000000101001000000000000000;
			// PEs: 41 -> 40
			// srcs: (94, 43)(1623) 0 --> (1623) 0:NI0, pass, PEGB0
			10'd25 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 40, 41 -> 40
			// srcs: (96, 25)(2018) -2, (2019) 0 --> (2799) -2:PENB, NI9, +, PEGB0
			10'd26 : rdata = 48'b000011101111111010100001001000000000000010000000;
			// PEs: 40 -> 
			// srcs: (98, 26)(2022) 0 --> (2022) 0:PENB, pass, 
			10'd27 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 40, 41 -> 41
			// srcs: (104, 27)(2021) 2, (2022) 0 --> (2802) 2:PENB, ALU, +, NI0
			10'd28 : rdata = 48'b000011101111111000111111111100000000000000000000;
			// PEs: 40 -> 41
			// srcs: (106, 28)(2098) 0 --> (2098) 0:PENB, pass, NI9
			10'd29 : rdata = 48'b110001101111111000000000000101001000000000000000;
			// PEs: 41 -> 40
			// srcs: (107, 50)(2445) -1 --> (2445) -1:NI7, pass, PEGB0
			10'd30 : rdata = 48'b110001010000011100000000000000000000000010000000;
			// PEs: 40, 41 -> 44
			// srcs: (112, 29)(2097) 6, (2098) 0 --> (2876) 6:PENB, NI9, +, PEGB4
			10'd31 : rdata = 48'b000011101111111010100001001000000000000011000000;
			// PEs: 40 -> 41
			// srcs: (114, 30)(2101) 6 --> (2101) 6:PENB, pass, NI7
			10'd32 : rdata = 48'b110001101111111000000000000100111000000000000000;
			// PEs: 41 -> 40
			// srcs: (117, 56)(1744) 1 --> (1744) 1:NI4, pass, PEGB0
			10'd33 : rdata = 48'b110001010000010000000000000000000000000010000000;
			// PEs: 40, 41 -> 47
			// srcs: (120, 31)(2100) -3, (2101) 6 --> (2880) 3:PENB, NI7, +, PEGB7
			10'd34 : rdata = 48'b000011101111111010100000111000000000000011110000;
			// PEs: 40 -> 41
			// srcs: (122, 32)(2104) 0 --> (2104) 0:PENB, pass, NI4
			10'd35 : rdata = 48'b110001101111111000000000000100100000000000000000;
			// PEs: 41 -> 40
			// srcs: (126, 75)(2802) 2 --> (2802) 2:NI0, pass, PEGB0
			10'd36 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 40, 41 -> 41
			// srcs: (128, 33)(2103) 0, (2104) 0 --> (2882) 0:PENB, NI4, +, NI0
			10'd37 : rdata = 48'b000011101111111010100000100100000000000000000000;
			// PEs: 40 -> 
			// srcs: (130, 34)(2178) 3 --> (2178) 3:PENB, pass, 
			10'd38 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 40, 41 -> 41
			// srcs: (136, 35)(2177) 0, (2178) 3 --> (2957) 3:PENB, ALU, +, NI4
			10'd39 : rdata = 48'b000011101111111000111111111100100000000000000000;
			// PEs: 40 -> 
			// srcs: (138, 36)(2181) 2 --> (2181) 2:PENB, pass, 
			10'd40 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 40, 41 -> 40
			// srcs: (144, 37)(2180) 0, (2181) 2 --> (2960) 2:PENB, ALU, +, PEGB0
			10'd41 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 40 -> 
			// srcs: (146, 38)(2184) -3 --> (2184) -3:PENB, pass, 
			10'd42 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 40, 41 -> 40
			// srcs: (152, 39)(2183) -2, (2184) -3 --> (2962) -5:PENB, ALU, +, PEGB0
			10'd43 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 40, 41 -> 40
			// srcs: (153, 40)(2186) 3, (2187) 2 --> (2967) 5:PENB, NI1, +, PEGB0
			10'd44 : rdata = 48'b000011101111111010100000001000000000000010000000;
			// PEs: 40, 41 -> 41
			// srcs: (154, 41)(2266) -3, (2267) 4 --> (3046) 1:PENB, NI2, +, NI1
			10'd45 : rdata = 48'b000011101111111010100000010100001000000000000000;
			// PEs: 40, 41 -> 40
			// srcs: (155, 42)(2348) -2, (2349) 0 --> (3125) -2:PENB, NI3, +, PEGB0
			10'd46 : rdata = 48'b000011101111111010100000011000000000000010000000;
			// PEs: 41 -> 40
			// srcs: (207, 62)(2657) -2 --> (2657) -2:NI8, pass, PEGB0
			10'd47 : rdata = 48'b110001010000100000000000000000000000000010000000;
			// PEs: 41 -> 40
			// srcs: (232, 83)(2957) 3 --> (2957) 3:NI4, pass, PEGB0
			10'd48 : rdata = 48'b110001010000010000000000000000000000000010000000;
			// PEs: 40 -> 41
			// srcs: (239, 44)(2017) 0 --> (2017) 0:PENB, pass, NI2
			10'd49 : rdata = 48'b110001101111111000000000000100010000000000000000;
			// PEs: 41 -> 40
			// srcs: (241, 86)(3046) 1 --> (3046) 1:NI1, pass, PEGB0
			10'd50 : rdata = 48'b110001010000000100000000000000000000000010000000;
			// PEs: 40, 41 -> 41
			// srcs: (245, 45)(2016) 1, (2017) 0 --> (2797) 1:PENB, NI2, +, NI1
			10'd51 : rdata = 48'b000011101111111010100000010100001000000000000000;
			// PEs: 40 -> 41
			// srcs: (247, 46)(1631) 0 --> (1631) 0:PENB, pass, NI2
			10'd52 : rdata = 48'b110001101111111000000000000100010000000000000000;
			// PEs: 41 -> 40
			// srcs: (249, 90)(2292) -2 --> (2292) -2:NI6, pass, PEGB0
			10'd53 : rdata = 48'b110001010000011000000000000000000000000010000000;
			// PEs: 40, 41 -> 40
			// srcs: (253, 47)(2411) 0, (1631) 0 --> (2412) 0:PENB, NI2, +, PEGB0
			10'd54 : rdata = 48'b000011101111111010100000010000000000000010000000;
			// PEs: 40 -> 
			// srcs: (255, 48)(1658) 4 --> (1658) 4:PENB, pass, 
			10'd55 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 40, 41 -> 40
			// srcs: (261, 49)(2436) 1, (1658) 4 --> (2437) 5:PENB, ALU, +, PEGB0
			10'd56 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 44, 40 -> 41
			// srcs: (262, 51)(2480) -2, (1701) -1 --> (2481) -3:PEGB4, PENB, +, NI2
			10'd57 : rdata = 48'b000011110000100011011111110100010000000000000000;
			// PEs: 40 -> 
			// srcs: (264, 52)(1710) 2 --> (1710) 2:PENB, pass, 
			10'd58 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 40, 41 -> 40
			// srcs: (270, 53)(2489) 0, (1710) 2 --> (2490) 2:PENB, ALU, +, PEGB0
			10'd59 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 40 -> 
			// srcs: (272, 54)(1738) 0 --> (1738) 0:PENB, pass, 
			10'd60 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 40, 41 -> 41
			// srcs: (278, 55)(2516) -2, (1738) 0 --> (2517) -2:PENB, ALU, +, NI3
			10'd61 : rdata = 48'b000011101111111000111111111100011000000000000000;
			// PEs: 40 -> 
			// srcs: (280, 57)(1793) -1 --> (1793) -1:PENB, pass, 
			10'd62 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 40, 41 -> 40
			// srcs: (286, 58)(2571) 0, (1793) -1 --> (2572) -1:PENB, ALU, +, PEGB0
			10'd63 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 40 -> 
			// srcs: (288, 59)(1836) 6 --> (1836) 6:PENB, pass, 
			10'd64 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 40, 41 -> 40
			// srcs: (294, 60)(2614) -2, (1836) 6 --> (2615) 4:PENB, ALU, +, PEGB0
			10'd65 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 42, 40 -> 40
			// srcs: (371, 61)(2635) 4, (1857) -2 --> (2636) 2:PEGB2, PENB, +, PEGB0
			10'd66 : rdata = 48'b000011110000010011011111110000000000000010000000;
			// PEs: 40 -> 
			// srcs: (373, 63)(1888) -2 --> (1888) -2:PENB, pass, 
			10'd67 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 40, 41 -> 40
			// srcs: (379, 64)(2666) -8, (1888) -2 --> (2667) -10:PENB, ALU, +, PEGB0
			10'd68 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 40 -> 
			// srcs: (381, 65)(1912) 3 --> (1912) 3:PENB, pass, 
			10'd69 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 40, 41 -> 40
			// srcs: (387, 66)(2689) -2, (1912) 3 --> (2690) 1:PENB, ALU, +, PEGB0
			10'd70 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 40, 41 -> 46
			// srcs: (388, 67)(2705) -4, (1928) -1 --> (2706) -5:PENB, NI5, +, PEGB6
			10'd71 : rdata = 48'b000011101111111010100000101000000000000011100000;
			// PEs: 40, 42 -> 41
			// srcs: (396, 68)(2709) -1, (1931) 0 --> (2710) -1:PENB, PEGB2, +, NI4
			10'd72 : rdata = 48'b000011101111111011100000100100100000000000000000;
			// PEs: 40, 43 -> 42
			// srcs: (397, 69)(2711) -4, (1934) -2 --> (2712) -6:PENB, PEGB3, +, PENB
			10'd73 : rdata = 48'b000011101111111011100000110000000000000100000000;
			// PEs: 40 -> 
			// srcs: (398, 70)(2010) -2 --> (2010) -2:PENB, pass, 
			10'd74 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 40, 41 -> 41
			// srcs: (403, 71)(2788) -3, (2010) -2 --> (2789) -5:PENB, ALU, +, NI5
			10'd75 : rdata = 48'b000011101111111000111111111100101000000000000000;
			// PEs: 41 -> 42
			// srcs: (404, 104)(2710) -1 --> (2710) -1:NI4, pass, PENB
			10'd76 : rdata = 48'b110001010000010000000000000000000000000100000000;
			// PEs: 40 -> 
			// srcs: (405, 72)(2013) 2 --> (2013) 2:PENB, pass, 
			10'd77 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 40, 41 -> 42
			// srcs: (411, 73)(2790) -10, (2013) 2 --> (2791) -8:PENB, ALU, +, PENB
			10'd78 : rdata = 48'b000011101111111000111111111000000000000100000000;
			// PEs: 40, 41 -> 40
			// srcs: (412, 74)(2796) 4, (2797) 1 --> (2798) 5:PENB, NI1, +, PEGB0
			10'd79 : rdata = 48'b000011101111111010100000001000000000000010000000;
			// PEs: 41 -> 42
			// srcs: (418, 105)(2789) -5 --> (2789) -5:NI5, pass, PENB
			10'd80 : rdata = 48'b110001010000010100000000000000000000000100000000;
			// PEs: 41, 40 -> 43
			// srcs: (627, 76)(2882) 0, (2105) -1 --> (2883) -1:NI0, PENB, +, PEGB3
			10'd81 : rdata = 48'b000011010000000011011111110000000000000010110000;
			// PEs: 40 -> 
			// srcs: (629, 77)(2142) -2 --> (2142) -2:PENB, pass, 
			10'd82 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 40, 41 -> 40
			// srcs: (635, 78)(2919) 0, (2142) -2 --> (2920) -2:PENB, ALU, +, PEGB0
			10'd83 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 40 -> 
			// srcs: (637, 79)(2157) 4 --> (2157) 4:PENB, pass, 
			10'd84 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 40, 41 -> 40
			// srcs: (643, 80)(2933) 4, (2157) 4 --> (2934) 8:PENB, ALU, +, PEGB0
			10'd85 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 40 -> 
			// srcs: (645, 81)(2170) -6 --> (2170) -6:PENB, pass, 
			10'd86 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 40, 41 -> 40
			// srcs: (651, 82)(2949) -2, (2170) -6 --> (2950) -8:PENB, ALU, +, PEGB0
			10'd87 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 40 -> 
			// srcs: (653, 84)(2203) 1 --> (2203) 1:PENB, pass, 
			10'd88 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 40, 41 -> 41
			// srcs: (659, 85)(2980) 4, (2203) 1 --> (2981) 5:PENB, ALU, +, NI0
			10'd89 : rdata = 48'b000011101111111000111111111100000000000000000000;
			// PEs: 42, 40 -> 40
			// srcs: (667, 87)(3048) -6, (2271) 4 --> (3049) -2:PEGB2, PENB, +, PEGB0
			10'd90 : rdata = 48'b000011110000010011011111110000000000000010000000;
			// PEs: 43, 40 -> 41
			// srcs: (676, 88)(3052) -6, (2274) 4 --> (3053) -2:PEGB3, PENB, +, NI1
			10'd91 : rdata = 48'b000011110000011011011111110100001000000000000000;
			// PEs: 44, 40 -> 42
			// srcs: (701, 89)(3054) -2, (2277) 0 --> (3055) -2:PEGB4, PENB, +, PENB
			10'd92 : rdata = 48'b000011110000100011011111110000000000000100000000;
			// PEs: 40 -> 
			// srcs: (702, 91)(2341) -4 --> (2341) -4:PENB, pass, 
			10'd93 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 40, 41 -> 40
			// srcs: (707, 92)(3117) -1, (2341) -4 --> (3118) -5:PENB, ALU, +, PEGB0
			10'd94 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 46, 40 -> 40
			// srcs: (708, 93)(3130) -2, (2356) 0 --> (3131) -2:PEGB6, PENB, +, PEGB0
			10'd95 : rdata = 48'b000011110000110011011111110000000000000010000000;
			// PEs: 41 -> 42
			// srcs: (709, 110)(3053) -2 --> (3053) -2:NI1, pass, PENB
			10'd96 : rdata = 48'b110001010000000100000000000000000000000100000000;
			// PEs: 40 -> 
			// srcs: (710, 94)(2400) 2 --> (2400) 2:PENB, pass, 
			10'd97 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 40, 41 -> 40
			// srcs: (716, 95)(2398) -10, (2400) 2 --> (2401) -8:PENB, ALU, +, PEGB0
			10'd98 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 40 -> 
			// srcs: (718, 96)(2443) 0 --> (2443) 0:PENB, pass, 
			10'd99 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 40, 41 -> 40
			// srcs: (724, 97)(2441) 2, (2443) 0 --> (2444) 2:PENB, ALU, +, PEGB0
			10'd100 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 40, 41 -> 41
			// srcs: (725, 98)(2479) 0, (2481) -3 --> (2482) -3:PENB, NI2, +, NI1
			10'd101 : rdata = 48'b000011101111111010100000010100001000000000000000;
			// PEs: 40, 41 -> 41
			// srcs: (726, 99)(2515) 1, (2517) -2 --> (2518) -1:PENB, NI3, +, NI2
			10'd102 : rdata = 48'b000011101111111010100000011100010000000000000000;
			// PEs: 40 -> 
			// srcs: (728, 100)(2545) -5 --> (2545) -5:PENB, pass, 
			10'd103 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 40, 41 -> 40
			// srcs: (734, 101)(2543) 0, (2545) -5 --> (2546) -5:PENB, ALU, +, PEGB0
			10'd104 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 40 -> 
			// srcs: (736, 102)(2643) -5 --> (2643) -5:PENB, pass, 
			10'd105 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 40, 41 -> 40
			// srcs: (742, 103)(2641) 7, (2643) -5 --> (2644) 2:PENB, ALU, +, PEGB0
			10'd106 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 40 -> 
			// srcs: (744, 106)(2811) -3 --> (2811) -3:PENB, pass, 
			10'd107 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 40, 41 -> 40
			// srcs: (750, 107)(2809) -6, (2811) -3 --> (2812) -9:PENB, ALU, +, PEGB0
			10'd108 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 40, 44 -> 41
			// srcs: (758, 108)(2875) 8, (2877) 6 --> (2878) 14:PENB, PEGB4, +, NI3
			10'd109 : rdata = 48'b000011101111111011100001000100011000000000000000;
			// PEs: 40, 41 -> 40
			// srcs: (759, 109)(2979) -7, (2981) 5 --> (2982) -2:PENB, NI0, +, PEGB0
			10'd110 : rdata = 48'b000011101111111010100000000000000000000010000000;
			// PEs: 40 -> 
			// srcs: (760, 111)(3083) -2 --> (3083) -2:PENB, pass, 
			10'd111 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 40, 41 -> 41
			// srcs: (765, 112)(3081) 1, (3083) -2 --> (3084) -1:PENB, ALU, +, NI0
			10'd112 : rdata = 48'b000011101111111000111111111100000000000000000000;
			// PEs: 40 -> 
			// srcs: (767, 113)(2367) -22 --> (2367) -22:PENB, pass, 
			10'd113 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 40, 41 -> 40
			// srcs: (773, 114)(2362) -7, (2367) -22 --> (2368) -29:PENB, ALU, +, PEGB0
			10'd114 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 41, 40 -> 40
			// srcs: (774, 115)(2482) -3, (2487) 14 --> (2488) 11:NI1, PENB, +, PEGB0
			10'd115 : rdata = 48'b000011010000000111011111110000000000000010000000;
			// PEs: 41, 40 -> 40
			// srcs: (775, 116)(2518) -1, (2523) 4 --> (2524) 3:NI2, PENB, +, PEGB0
			10'd116 : rdata = 48'b000011010000001011011111110000000000000010000000;
			// PEs: 40 -> 
			// srcs: (777, 117)(2659) -2 --> (2659) -2:PENB, pass, 
			10'd117 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 40, 41 -> 41
			// srcs: (783, 118)(2654) 10, (2659) -2 --> (2660) 8:PENB, ALU, +, NI1
			10'd118 : rdata = 48'b000011101111111000111111111100001000000000000000;
			// PEs: 40 -> 
			// srcs: (785, 119)(2829) -9 --> (2829) -9:PENB, pass, 
			10'd119 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 40, 41 -> 40
			// srcs: (791, 120)(2824) 10, (2829) -9 --> (2830) 1:PENB, ALU, +, PEGB0
			10'd120 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 40, 41 -> 40
			// srcs: (1117, 121)(2873) -2, (2878) 14 --> (2879) 12:PENB, NI3, +, PEGB0
			10'd121 : rdata = 48'b000011101111111010100000011000000000000010000000;
			// PEs: 40, 41 -> 41
			// srcs: (1118, 122)(3079) 2, (3084) -1 --> (3085) 1:PENB, NI0, +, NI2
			10'd122 : rdata = 48'b000011101111111010100000000100010000000000000000;
			// PEs: 40 -> 
			// srcs: (1120, 123)(2427) -7 --> (2427) -7:PENB, pass, 
			10'd123 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 40, 41 -> 40
			// srcs: (1127, 124)(2416) 3, (2427) -7 --> (2428) -4:PENB, ALU, +, PEGB0
			10'd124 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 41, 40 -> 40
			// srcs: (1128, 125)(2660) 8, (2671) -14 --> (2672) -6:NI1, PENB, +, PEGB0
			10'd125 : rdata = 48'b000011010000000111011111110000000000000010000000;
			// PEs: 40 -> 
			// srcs: (1130, 126)(2867) 2 --> (2867) 2:PENB, pass, 
			10'd126 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 40, 41 -> 40
			// srcs: (1138, 127)(2856) 9, (2867) 2 --> (2868) 11:PENB, ALU, +, PEGB0
			10'd127 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 40, 41 -> 40
			// srcs: (1139, 128)(3074) -1, (3085) 1 --> (3086) 0:PENB, NI2, +, PEGB0
			10'd128 : rdata = 48'b000011101111111010100000010000000000000010000000;
			// PEs: 40 -> 
			// srcs: (1180, 129)(2646) 21 --> (2646) 21:PENB, pass, 
			10'd129 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 40, 41 -> 40
			// srcs: (1186, 130)(2623) 27, (2646) 21 --> (2647) 48:PENB, ALU, +, PEGB0
			10'd130 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 40 -> 
			// srcs: (1189, 131)(2549) -2 --> (2549) -2:PENB, pass, 
			10'd131 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 40, 41 -> 40
			// srcs: (1195, 132)(2501) 26, (2549) -2 --> (2550) 24:PENB, ALU, +, PEGB0
			10'd132 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 40 -> 
			// srcs: (1449, 133)(3136) -25 --> (3136) -25:PENB, pass, 
			10'd133 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 40, 41 -> 40
			// srcs: (1456, 134)(3039) -38, (3136) -25 --> (3137) -63:PENB, ALU, +, PEGB0
			10'd134 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 40, 41 -> 42
			// srcs: (1561, 135)(3140) 47, (54) 0 --> (3191) 0:PENB, ND0, *, PENB
			10'd135 : rdata = 48'b000111101111111001100000000000000000000100000000;
			// PEs: 41, 42 -> 41
			// srcs: (1570, 149)(839) -2, (3975) 0 --> (4759) -2:NW0, PEGB2, -, NW0
			10'd136 : rdata = 48'b000100100000000011100000100000000100000000000000;
			// PEs: 40, 41 -> 42
			// srcs: (1641, 136)(3140) 47, (134) -3 --> (3271) -141:PENB, ND1, *, PENB
			10'd137 : rdata = 48'b000111101111111001100000001000000000000100000000;
			// PEs: 41, 42 -> 41
			// srcs: (1650, 150)(919) -1, (4055) -141 --> (4839) 140:NW1, PEGB2, -, NW1
			10'd138 : rdata = 48'b000100100000000111100000100000000100010000000000;
			// PEs: 40, 41 -> 42
			// srcs: (1682, 137)(3140) 47, (175) 1 --> (3312) 47:PENB, ND10, *, PENB
			10'd139 : rdata = 48'b000111101111111001100001010000000000000100000000;
			// PEs: 41, 42 -> 41
			// srcs: (1691, 151)(960) 1, (4096) 47 --> (4880) -46:NW10, PEGB2, -, NW10
			10'd140 : rdata = 48'b000100100000101011100000100000000110100000000000;
			// PEs: 40, 41 -> 42
			// srcs: (1721, 138)(3140) 47, (214) 1 --> (3351) 47:PENB, ND2, *, PENB
			10'd141 : rdata = 48'b000111101111111001100000010000000000000100000000;
			// PEs: 41, 42 -> 41
			// srcs: (1730, 152)(999) 2, (4135) 47 --> (4919) -45:NW2, PEGB2, -, NW2
			10'd142 : rdata = 48'b000100100000001011100000100000000100100000000000;
			// PEs: 40, 41 -> 42
			// srcs: (1803, 139)(3140) 47, (296) 1 --> (3433) 47:PENB, ND3, *, PENB
			10'd143 : rdata = 48'b000111101111111001100000011000000000000100000000;
			// PEs: 41, 42 -> 41
			// srcs: (1812, 153)(1081) -3, (4217) 47 --> (5001) -50:NW3, PEGB2, -, NW3
			10'd144 : rdata = 48'b000100100000001111100000100000000100110000000000;
			// PEs: 40, 41 -> 42
			// srcs: (1866, 140)(3140) 47, (359) 1 --> (3496) 47:PENB, ND11, *, PENB
			10'd145 : rdata = 48'b000111101111111001100001011000000000000100000000;
			// PEs: 41, 42 -> 41
			// srcs: (1875, 154)(1144) -1, (4280) 47 --> (5064) -48:NW11, PEGB2, -, NW11
			10'd146 : rdata = 48'b000100100000101111100000100000000110110000000000;
			// PEs: 40, 41 -> 42
			// srcs: (1883, 141)(3140) 47, (376) -2 --> (3513) -94:PENB, ND4, *, PENB
			10'd147 : rdata = 48'b000111101111111001100000100000000000000100000000;
			// PEs: 41, 42 -> 41
			// srcs: (1892, 155)(1161) 1, (4297) -94 --> (5081) 95:NW4, PEGB2, -, NW4
			10'd148 : rdata = 48'b000100100000010011100000100000000101000000000000;
			// PEs: 40, 41 -> 42
			// srcs: (1963, 142)(3140) 47, (456) 0 --> (3593) 0:PENB, ND5, *, PENB
			10'd149 : rdata = 48'b000111101111111001100000101000000000000100000000;
			// PEs: 41, 42 -> 41
			// srcs: (1972, 156)(1241) -1, (4377) 0 --> (5161) -1:NW5, PEGB2, -, NW5
			10'd150 : rdata = 48'b000100100000010111100000100000000101010000000000;
			// PEs: 40, 41 -> 42
			// srcs: (2045, 143)(3140) 47, (538) -3 --> (3675) -141:PENB, ND6, *, PENB
			10'd151 : rdata = 48'b000111101111111001100000110000000000000100000000;
			// PEs: 40, 41 -> 42
			// srcs: (2046, 144)(3140) 47, (539) -3 --> (3676) -141:PENB, ND12, *, PENB
			10'd152 : rdata = 48'b000111101111111001100001100000000000000100000000;
			// PEs: 41, 42 -> 41
			// srcs: (2054, 157)(1323) -1, (4459) -141 --> (5243) 140:NW6, PEGB2, -, NW6
			10'd153 : rdata = 48'b000100100000011011100000100000000101100000000000;
			// PEs: 41, 42 -> 41
			// srcs: (2055, 158)(1324) 2, (4460) -141 --> (5244) 143:NW12, PEGB2, -, NW12
			10'd154 : rdata = 48'b000100100000110011100000100000000111000000000000;
			// PEs: 40, 41 -> 42
			// srcs: (2125, 145)(3140) 47, (618) 1 --> (3755) 47:PENB, ND7, *, PENB
			10'd155 : rdata = 48'b000111101111111001100000111000000000000100000000;
			// PEs: 41, 42 -> 41
			// srcs: (2134, 159)(1403) 2, (4539) 47 --> (5323) -45:NW7, PEGB2, -, NW7
			10'd156 : rdata = 48'b000100100000011111100000100000000101110000000000;
			// PEs: 40, 41 -> 42
			// srcs: (2205, 146)(3140) 47, (698) 2 --> (3835) 94:PENB, ND8, *, PENB
			10'd157 : rdata = 48'b000111101111111001100001000000000000000100000000;
			// PEs: 41, 42 -> 41
			// srcs: (2214, 160)(1483) 2, (4619) 94 --> (5403) -92:NW8, PEGB2, -, NW8
			10'd158 : rdata = 48'b000100100000100011100000100000000110000000000000;
			// PEs: 40, 41 -> 42
			// srcs: (2230, 147)(3140) 47, (723) -2 --> (3860) -94:PENB, ND13, *, PENB
			10'd159 : rdata = 48'b000111101111111001100001101000000000000100000000;
			// PEs: 41, 42 -> 41
			// srcs: (2239, 161)(1508) 1, (4644) -94 --> (5428) 95:NW13, PEGB2, -, NW13
			10'd160 : rdata = 48'b000100100000110111100000100000000111010000000000;
			// PEs: 40, 41 -> 42
			// srcs: (2287, 148)(3140) 47, (780) 0 --> (3917) 0:PENB, ND9, *, PENB
			10'd161 : rdata = 48'b000111101111111001100001001000000000000100000000;
			// PEs: 41, 42 -> 41
			// srcs: (2296, 162)(1565) -1, (4701) 0 --> (5485) -1:NW9, PEGB2, -, NW9
			10'd162 : rdata = 48'b000100100000100111100000100000000110010000000000;
			default : rdata = 48'b000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 42) begin
	always @(*) begin
		case(address)
			// PEs: 42, 42 -> 42
			// srcs: (1, 0)(55) 2, (840) 0 --> (1624) 0:ND0, NW0, *, NI0
			10'd0 : rdata = 48'b000110110000000001000000000100000000000000000000;
			// PEs: 42, 42 -> 40
			// srcs: (2, 1)(136) -3, (921) -2 --> (1705) 6:ND1, NW1, *, PEGB0
			10'd1 : rdata = 48'b000110110000000101000000001000000000000010000000;
			// PEs: 42, 42 -> 40
			// srcs: (3, 2)(216) 1, (1001) 2 --> (1785) 2:ND2, NW2, *, PEGB0
			10'd2 : rdata = 48'b000110110000001001000000010000000000000010000000;
			// PEs: 42, 42 -> 42
			// srcs: (4, 3)(298) -3, (1083) -2 --> (1867) 6:ND3, NW3, *, NI1
			10'd3 : rdata = 48'b000110110000001101000000011100001000000000000000;
			// PEs: 42, 42 -> 40
			// srcs: (5, 4)(378) 1, (1163) 1 --> (1947) 1:ND4, NW4, *, PEGB0
			10'd4 : rdata = 48'b000110110000010001000000100000000000000010000000;
			// PEs: 42, 42 -> 40
			// srcs: (6, 5)(458) -3, (1243) 2 --> (2027) -6:ND5, NW5, *, PEGB0
			10'd5 : rdata = 48'b000110110000010101000000101000000000000010000000;
			// PEs: 42, 42 -> 40
			// srcs: (7, 6)(540) -2, (1325) -3 --> (2109) 6:ND6, NW6, *, PEGB0
			10'd6 : rdata = 48'b000110110000011001000000110000000000000010000000;
			// PEs: 42, 42 -> 40
			// srcs: (8, 7)(620) -1, (1405) 2 --> (2189) -2:ND7, NW7, *, PEGB0
			10'd7 : rdata = 48'b000110110000011101000000111000000000000010000000;
			// PEs: 42, 42 -> 42
			// srcs: (9, 8)(700) -3, (1485) 2 --> (2269) -6:ND8, NW8, *, NI2
			10'd8 : rdata = 48'b000110110000100001000001000100010000000000000000;
			// PEs: 42, 42 -> 45
			// srcs: (10, 9)(782) 1, (1567) -1 --> (2351) -1:ND9, NW9, *, PEGB5
			10'd9 : rdata = 48'b000110110000100101000001001000000000000011010000;
			// PEs: 42, 42 -> 42
			// srcs: (11, 10)(178) 1, (963) 0 --> (1747) 0:ND10, NW10, *, NI3
			10'd10 : rdata = 48'b000110110000101001000001010100011000000000000000;
			// PEs: 42, 42 -> 42
			// srcs: (12, 11)(362) -1, (1147) 0 --> (1931) 0:ND11, NW11, *, NI4
			10'd11 : rdata = 48'b000110110000101101000001011100100000000000000000;
			// PEs: 42, 42 -> 42
			// srcs: (13, 12)(542) 0, (1327) 1 --> (2111) 0:ND12, NW12, *, NI5
			10'd12 : rdata = 48'b000110110000110001000001100100101000000000000000;
			// PEs: 42, 42 -> 42
			// srcs: (14, 13)(726) 1, (1511) 1 --> (2295) 1:ND13, NW13, *, NI6
			10'd13 : rdata = 48'b000110110000110101000001101100110000000000000000;
			// PEs: 42, 43 -> 42
			// srcs: (15, 18)(2269) -6, (2270) 0 --> (3048) -6:NI2, PEGB3, +, NI7
			10'd14 : rdata = 48'b000011010000001011100000110100111000000000000000;
			// PEs: 40 -> 
			// srcs: (20, 14)(1694) -6 --> (1694) -6:PEGB0, pass, 
			10'd15 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 40, 42 -> 42
			// srcs: (29, 15)(1693) 0, (1694) -6 --> (2473) -6:PEGB0, ALU, +, NI2
			10'd16 : rdata = 48'b000011110000000000111111111100010000000000000000;
			// PEs: 40 -> 
			// srcs: (51, 16)(1856) 0 --> (1856) 0:PEGB0, pass, 
			10'd17 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 40, 42 -> 41
			// srcs: (60, 17)(1855) 4, (1856) 0 --> (2635) 4:PEGB0, ALU, +, PEGB1
			10'd18 : rdata = 48'b000011110000000000111111111000000000000010010000;
			// PEs: 42 -> 40
			// srcs: (94, 19)(1624) 0 --> (1624) 0:NI0, pass, PEGB0
			10'd19 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 42 -> 40
			// srcs: (95, 20)(1867) 6 --> (1867) 6:NI1, pass, PEGB0
			10'd20 : rdata = 48'b110001010000000100000000000000000000000010000000;
			// PEs: 42 -> 40
			// srcs: (107, 22)(1747) 0 --> (1747) 0:NI3, pass, PEGB0
			10'd21 : rdata = 48'b110001010000001100000000000000000000000010000000;
			// PEs: 42 -> 40
			// srcs: (131, 27)(2295) 1 --> (2295) 1:NI6, pass, PEGB0
			10'd22 : rdata = 48'b110001010000011000000000000000000000000010000000;
			// PEs: 47, 41 -> 42
			// srcs: (134, 24)(2885) -3, (2108) -6 --> (2886) -9:PEGB7, PENB, +, NI0
			10'd23 : rdata = 48'b000011110000111011011111110100000000000000000000;
			// PEs: 42 -> 40
			// srcs: (162, 21)(2473) -6 --> (2473) -6:NI2, pass, PEGB0
			10'd24 : rdata = 48'b110001010000001000000000000000000000000010000000;
			// PEs: 42 -> 40
			// srcs: (224, 25)(2111) 0 --> (2111) 0:NI5, pass, PEGB0
			10'd25 : rdata = 48'b110001010000010100000000000000000000000010000000;
			// PEs: 42 -> 41
			// srcs: (391, 23)(1931) 0 --> (1931) 0:NI4, pass, PEGB1
			10'd26 : rdata = 48'b110001010000010000000000000000000000000010010000;
			// PEs: 42 -> 40
			// srcs: (395, 32)(2886) -9 --> (2886) -9:NI0, pass, PEGB0
			10'd27 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 41 -> 
			// srcs: (399, 28)(2712) -6 --> (2712) -6:PENB, pass, 
			10'd28 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 41, 42 -> 46
			// srcs: (406, 29)(2710) -1, (2712) -6 --> (2713) -7:PENB, ALU, +, PEGB6
			10'd29 : rdata = 48'b000011101111111000111111111000000000000011100000;
			// PEs: 41 -> 
			// srcs: (413, 30)(2791) -8 --> (2791) -8:PENB, pass, 
			10'd30 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 41, 42 -> 40
			// srcs: (420, 31)(2789) -5, (2791) -8 --> (2792) -13:PENB, ALU, +, PEGB0
			10'd31 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 42 -> 41
			// srcs: (662, 26)(3048) -6 --> (3048) -6:NI7, pass, PEGB1
			10'd32 : rdata = 48'b110001010000011100000000000000000000000010010000;
			// PEs: 41 -> 
			// srcs: (703, 33)(3055) -2 --> (3055) -2:PENB, pass, 
			10'd33 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 41, 42 -> 40
			// srcs: (711, 34)(3053) -2, (3055) -2 --> (3056) -4:PENB, ALU, +, PEGB0
			10'd34 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 42, 41 -> 41
			// srcs: (1564, 49)(3) 1, (3191) 0 --> (3975) 0:NM0, PENB, *, PEGB1
			10'd35 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 40, 42 -> 43
			// srcs: (1565, 35)(3140) 47, (55) 2 --> (3192) 94:PEGB0, ND0, *, PENB
			10'd36 : rdata = 48'b000111110000000001100000000000000000000100000000;
			// PEs: 42, 43 -> 42
			// srcs: (1574, 66)(840) 0, (3976) 94 --> (4760) -94:NW0, PEGB3, -, NW0
			10'd37 : rdata = 48'b000100100000000011100000110000000100000000000000;
			// PEs: 42, 41 -> 41
			// srcs: (1644, 50)(3) 1, (3271) -141 --> (4055) -141:NM0, PENB, *, PEGB1
			10'd38 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 40, 42 -> 43
			// srcs: (1646, 36)(3140) 47, (136) -3 --> (3273) -141:PEGB0, ND1, *, PENB
			10'd39 : rdata = 48'b000111110000000001100000001000000000000100000000;
			// PEs: 42, 43 -> 42
			// srcs: (1655, 67)(921) -2, (4057) -141 --> (4841) 139:NW1, PEGB3, -, NW1
			10'd40 : rdata = 48'b000100100000000111100000110000000100010000000000;
			// PEs: 42, 41 -> 41
			// srcs: (1685, 51)(3) 1, (3312) 47 --> (4096) 47:NM0, PENB, *, PEGB1
			10'd41 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 40, 42 -> 
			// srcs: (1688, 37)(3140) 47, (178) 1 --> (3315) 47:PEGB0, ND10, *, 
			10'd42 : rdata = 48'b000111110000000001100001010000000000000000000000;
			// PEs: 42, 42 -> 
			// srcs: (1691, 52)(3) 1, (3315) 47 --> (4099) 47:NM0, ALU, *, 
			10'd43 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 42, 42 -> 42
			// srcs: (1694, 68)(963) 0, (4099) 47 --> (4883) -47:NW10, ALU, -, NW10
			10'd44 : rdata = 48'b000100100000101000111111111000000110100000000000;
			// PEs: 42, 41 -> 41
			// srcs: (1724, 53)(3) 1, (3351) 47 --> (4135) 47:NM0, PENB, *, PEGB1
			10'd45 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 40, 42 -> 43
			// srcs: (1726, 38)(3140) 47, (216) 1 --> (3353) 47:PEGB0, ND2, *, PENB
			10'd46 : rdata = 48'b000111110000000001100000010000000000000100000000;
			// PEs: 42, 43 -> 42
			// srcs: (1735, 69)(1001) 2, (4137) 47 --> (4921) -45:NW2, PEGB3, -, NW2
			10'd47 : rdata = 48'b000100100000001011100000110000000100100000000000;
			// PEs: 42, 41 -> 41
			// srcs: (1806, 54)(3) 1, (3433) 47 --> (4217) 47:NM0, PENB, *, PEGB1
			10'd48 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 40, 42 -> 43
			// srcs: (1808, 39)(3140) 47, (298) -3 --> (3435) -141:PEGB0, ND3, *, PENB
			10'd49 : rdata = 48'b000111110000000001100000011000000000000100000000;
			// PEs: 42, 43 -> 42
			// srcs: (1817, 70)(1083) -2, (4219) -141 --> (5003) 139:NW3, PEGB3, -, NW3
			10'd50 : rdata = 48'b000100100000001111100000110000000100110000000000;
			// PEs: 42, 41 -> 41
			// srcs: (1869, 55)(3) 1, (3496) 47 --> (4280) 47:NM0, PENB, *, PEGB1
			10'd51 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 40, 42 -> 
			// srcs: (1872, 40)(3140) 47, (362) -1 --> (3499) -47:PEGB0, ND11, *, 
			10'd52 : rdata = 48'b000111110000000001100001011000000000000000000000;
			// PEs: 42, 42 -> 
			// srcs: (1875, 56)(3) 1, (3499) -47 --> (4283) -47:NM0, ALU, *, 
			10'd53 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 42, 42 -> 42
			// srcs: (1878, 71)(1147) 0, (4283) -47 --> (5067) 47:NW11, ALU, -, NW11
			10'd54 : rdata = 48'b000100100000101100111111111000000110110000000000;
			// PEs: 42, 41 -> 41
			// srcs: (1886, 57)(3) 1, (3513) -94 --> (4297) -94:NM0, PENB, *, PEGB1
			10'd55 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 40, 42 -> 43
			// srcs: (1888, 41)(3140) 47, (378) 1 --> (3515) 47:PEGB0, ND4, *, PENB
			10'd56 : rdata = 48'b000111110000000001100000100000000000000100000000;
			// PEs: 42, 43 -> 42
			// srcs: (1897, 72)(1163) 1, (4299) 47 --> (5083) -46:NW4, PEGB3, -, NW4
			10'd57 : rdata = 48'b000100100000010011100000110000000101000000000000;
			// PEs: 42, 41 -> 41
			// srcs: (1966, 58)(3) 1, (3593) 0 --> (4377) 0:NM0, PENB, *, PEGB1
			10'd58 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 40, 42 -> 43
			// srcs: (1968, 42)(3140) 47, (458) -3 --> (3595) -141:PEGB0, ND5, *, PENB
			10'd59 : rdata = 48'b000111110000000001100000101000000000000100000000;
			// PEs: 42, 43 -> 42
			// srcs: (1977, 73)(1243) 2, (4379) -141 --> (5163) 143:NW5, PEGB3, -, NW5
			10'd60 : rdata = 48'b000100100000010111100000110000000101010000000000;
			// PEs: 42, 41 -> 41
			// srcs: (2048, 59)(3) 1, (3675) -141 --> (4459) -141:NM0, PENB, *, PEGB1
			10'd61 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 42, 41 -> 41
			// srcs: (2049, 60)(3) 1, (3676) -141 --> (4460) -141:NM0, PENB, *, PEGB1
			10'd62 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 40, 42 -> 43
			// srcs: (2050, 43)(3140) 47, (540) -2 --> (3677) -94:PEGB0, ND6, *, PENB
			10'd63 : rdata = 48'b000111110000000001100000110000000000000100000000;
			// PEs: 40, 42 -> 43
			// srcs: (2052, 44)(3140) 47, (542) 0 --> (3679) 0:PEGB0, ND12, *, PENB
			10'd64 : rdata = 48'b000111110000000001100001100000000000000100000000;
			// PEs: 42, 43 -> 42
			// srcs: (2059, 74)(1325) -3, (4461) -94 --> (5245) 91:NW6, PEGB3, -, NW6
			10'd65 : rdata = 48'b000100100000011011100000110000000101100000000000;
			// PEs: 42, 43 -> 42
			// srcs: (2061, 75)(1327) 1, (4463) 0 --> (5247) 1:NW12, PEGB3, -, NW12
			10'd66 : rdata = 48'b000100100000110011100000110000000111000000000000;
			// PEs: 42, 41 -> 41
			// srcs: (2128, 61)(3) 1, (3755) 47 --> (4539) 47:NM0, PENB, *, PEGB1
			10'd67 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 40, 42 -> 43
			// srcs: (2130, 45)(3140) 47, (620) -1 --> (3757) -47:PEGB0, ND7, *, PENB
			10'd68 : rdata = 48'b000111110000000001100000111000000000000100000000;
			// PEs: 42, 43 -> 42
			// srcs: (2139, 76)(1405) 2, (4541) -47 --> (5325) 49:NW7, PEGB3, -, NW7
			10'd69 : rdata = 48'b000100100000011111100000110000000101110000000000;
			// PEs: 42, 41 -> 41
			// srcs: (2208, 62)(3) 1, (3835) 94 --> (4619) 94:NM0, PENB, *, PEGB1
			10'd70 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 40, 42 -> 43
			// srcs: (2210, 46)(3140) 47, (700) -3 --> (3837) -141:PEGB0, ND8, *, PENB
			10'd71 : rdata = 48'b000111110000000001100001000000000000000100000000;
			// PEs: 42, 43 -> 42
			// srcs: (2219, 77)(1485) 2, (4621) -141 --> (5405) 143:NW8, PEGB3, -, NW8
			10'd72 : rdata = 48'b000100100000100011100000110000000110000000000000;
			// PEs: 42, 41 -> 41
			// srcs: (2233, 63)(3) 1, (3860) -94 --> (4644) -94:NM0, PENB, *, PEGB1
			10'd73 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 40, 42 -> 
			// srcs: (2236, 47)(3140) 47, (726) 1 --> (3863) 47:PEGB0, ND13, *, 
			10'd74 : rdata = 48'b000111110000000001100001101000000000000000000000;
			// PEs: 42, 42 -> 
			// srcs: (2239, 64)(3) 1, (3863) 47 --> (4647) 47:NM0, ALU, *, 
			10'd75 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 42, 42 -> 42
			// srcs: (2242, 78)(1511) 1, (4647) 47 --> (5431) -46:NW13, ALU, -, NW13
			10'd76 : rdata = 48'b000100100000110100111111111000000111010000000000;
			// PEs: 42, 41 -> 41
			// srcs: (2290, 65)(3) 1, (3917) 0 --> (4701) 0:NM0, PENB, *, PEGB1
			10'd77 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 40, 42 -> 43
			// srcs: (2292, 48)(3140) 47, (782) 1 --> (3919) 47:PEGB0, ND9, *, PENB
			10'd78 : rdata = 48'b000111110000000001100001001000000000000100000000;
			// PEs: 42, 43 -> 42
			// srcs: (2301, 79)(1567) -1, (4703) 47 --> (5487) -48:NW9, PEGB3, -, NW9
			10'd79 : rdata = 48'b000100100000100111100000110000000110010000000000;
			default : rdata = 48'b000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 43) begin
	always @(*) begin
		case(address)
			// PEs: 43, 43 -> 43
			// srcs: (1, 0)(56) -2, (841) -2 --> (1625) 4:ND0, NW0, *, NI0
			10'd0 : rdata = 48'b000110110000000001000000000100000000000000000000;
			// PEs: 43, 43 -> 40
			// srcs: (2, 1)(137) 2, (922) 1 --> (1706) 2:ND1, NW1, *, PEGB0
			10'd1 : rdata = 48'b000110110000000101000000001000000000000010000000;
			// PEs: 43, 43 -> 40
			// srcs: (3, 2)(217) 1, (1002) 2 --> (1786) 2:ND2, NW2, *, PEGB0
			10'd2 : rdata = 48'b000110110000001001000000010000000000000010000000;
			// PEs: 43, 43 -> 43
			// srcs: (4, 3)(299) 1, (1084) -1 --> (1868) -1:ND3, NW3, *, NI1
			10'd3 : rdata = 48'b000110110000001101000000011100001000000000000000;
			// PEs: 43, 43 -> 40
			// srcs: (5, 4)(379) 2, (1164) -1 --> (1948) -2:ND4, NW4, *, PEGB0
			10'd4 : rdata = 48'b000110110000010001000000100000000000000010000000;
			// PEs: 43, 43 -> 40
			// srcs: (6, 5)(459) 2, (1244) 0 --> (2028) 0:ND5, NW5, *, PEGB0
			10'd5 : rdata = 48'b000110110000010101000000101000000000000010000000;
			// PEs: 43, 43 -> 40
			// srcs: (7, 6)(541) -2, (1326) -3 --> (2110) 6:ND6, NW6, *, PEGB0
			10'd6 : rdata = 48'b000110110000011001000000110000000000000010000000;
			// PEs: 43, 43 -> 40
			// srcs: (8, 7)(621) -1, (1406) 2 --> (2190) -2:ND7, NW7, *, PEGB0
			10'd7 : rdata = 48'b000110110000011101000000111000000000000010000000;
			// PEs: 43, 43 -> 42
			// srcs: (9, 8)(701) -3, (1486) 0 --> (2270) 0:ND8, NW8, *, PEGB2
			10'd8 : rdata = 48'b000110110000100001000001000000000000000010100000;
			// PEs: 43, 43 -> 45
			// srcs: (10, 9)(783) -3, (1568) -3 --> (2352) 9:ND9, NW9, *, PEGB5
			10'd9 : rdata = 48'b000110110000100101000001001000000000000011010000;
			// PEs: 43, 43 -> 43
			// srcs: (11, 10)(181) 0, (966) 2 --> (1750) 0:ND10, NW10, *, NI2
			10'd10 : rdata = 48'b000110110000101001000001010100010000000000000000;
			// PEs: 43, 43 -> 41
			// srcs: (12, 11)(365) 1, (1150) -2 --> (1934) -2:ND11, NW11, *, PEGB1
			10'd11 : rdata = 48'b000110110000101101000001011000000000000010010000;
			// PEs: 43, 43 -> 43
			// srcs: (13, 12)(549) 2, (1334) -1 --> (2118) -2:ND12, NW12, *, NI3
			10'd12 : rdata = 48'b000110110000110001000001100100011000000000000000;
			// PEs: 43, 43 -> 43
			// srcs: (14, 13)(729) 0, (1514) -2 --> (2298) 0:ND13, NW13, *, NI4
			10'd13 : rdata = 48'b000110110000110101000001101100100000000000000000;
			// PEs: 45 -> 
			// srcs: (15, 18)(2273) -2 --> (2273) -2:PEGB5, pass, 
			10'd14 : rdata = 48'b110001110000101000000000000000000000000000000000;
			// PEs: 44, 43 -> 41
			// srcs: (17, 19)(2272) -4, (2273) -2 --> (3052) -6:PEGB4, ALU, +, PEGB1
			10'd15 : rdata = 48'b000011110000100000111111111000000000000010010000;
			// PEs: 40 -> 
			// srcs: (22, 14)(1697) 2 --> (1697) 2:PEGB0, pass, 
			10'd16 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 40, 43 -> 40
			// srcs: (31, 15)(1696) 2, (1697) 2 --> (2478) 4:PEGB0, ALU, +, PEGB0
			10'd17 : rdata = 48'b000011110000000000111111111000000000000010000000;
			// PEs: 40 -> 
			// srcs: (53, 16)(1859) -4 --> (1859) -4:PEGB0, pass, 
			10'd18 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 40, 43 -> 43
			// srcs: (62, 17)(1858) 2, (1859) -4 --> (2637) -2:PEGB0, ALU, +, NI5
			10'd19 : rdata = 48'b000011110000000000111111111100101000000000000000;
			// PEs: 43 -> 40
			// srcs: (103, 20)(1625) 4 --> (1625) 4:NI0, pass, PEGB0
			10'd20 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 43 -> 40
			// srcs: (107, 21)(1868) -1 --> (1868) -1:NI1, pass, PEGB0
			10'd21 : rdata = 48'b110001010000000100000000000000000000000010000000;
			// PEs: 43 -> 40
			// srcs: (108, 22)(1750) 0 --> (1750) 0:NI2, pass, PEGB0
			10'd22 : rdata = 48'b110001010000001000000000000000000000000010000000;
			// PEs: 43 -> 40
			// srcs: (126, 24)(2118) -2 --> (2118) -2:NI3, pass, PEGB0
			10'd23 : rdata = 48'b110001010000001100000000000000000000000010000000;
			// PEs: 43 -> 40
			// srcs: (157, 25)(2298) 0 --> (2298) 0:NI4, pass, PEGB0
			10'd24 : rdata = 48'b110001010000010000000000000000000000000010000000;
			// PEs: 43 -> 40
			// srcs: (199, 23)(2637) -2 --> (2637) -2:NI5, pass, PEGB0
			10'd25 : rdata = 48'b110001010000010100000000000000000000000010000000;
			// PEs: 41 -> 
			// srcs: (632, 26)(2883) -1 --> (2883) -1:PEGB1, pass, 
			10'd26 : rdata = 48'b110001110000001000000000000000000000000000000000;
			// PEs: 47, 43 -> 40
			// srcs: (635, 27)(2881) 3, (2883) -1 --> (2884) 2:PEGB7, ALU, +, PEGB0
			10'd27 : rdata = 48'b000011110000111000111111111000000000000010000000;
			// PEs: 40, 43 -> 43
			// srcs: (1566, 28)(3140) 47, (56) -2 --> (3193) -94:PEGB0, ND0, *, NI0
			10'd28 : rdata = 48'b000111110000000001100000000100000000000000000000;
			// PEs: 43, 42 -> 42
			// srcs: (1568, 42)(3) 1, (3192) 94 --> (3976) 94:NM0, PENB, *, PEGB2
			10'd29 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 43, 43 -> 
			// srcs: (1569, 43)(3) 1, (3193) -94 --> (3977) -94:NM0, NI0, *, 
			10'd30 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 43, 43 -> 43
			// srcs: (1572, 59)(841) -2, (3977) -94 --> (4761) 92:NW0, ALU, -, NW0
			10'd31 : rdata = 48'b000100100000000000111111111000000100000000000000;
			// PEs: 40, 43 -> 44
			// srcs: (1647, 29)(3140) 47, (137) 2 --> (3274) 94:PEGB0, ND1, *, PENB
			10'd32 : rdata = 48'b000111110000000001100000001000000000000100000000;
			// PEs: 43, 42 -> 42
			// srcs: (1649, 44)(3) 1, (3273) -141 --> (4057) -141:NM0, PENB, *, PEGB2
			10'd33 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 43, 44 -> 43
			// srcs: (1656, 60)(922) 1, (4058) 94 --> (4842) -93:NW1, PEGB4, -, NW1
			10'd34 : rdata = 48'b000100100000000111100001000000000100010000000000;
			// PEs: 40, 43 -> 
			// srcs: (1691, 30)(3140) 47, (181) 0 --> (3318) 0:PEGB0, ND10, *, 
			10'd35 : rdata = 48'b000111110000000001100001010000000000000000000000;
			// PEs: 43, 43 -> 
			// srcs: (1694, 45)(3) 1, (3318) 0 --> (4102) 0:NM0, ALU, *, 
			10'd36 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 43, 43 -> 43
			// srcs: (1697, 61)(966) 2, (4102) 0 --> (4886) 2:NW10, ALU, -, NW10
			10'd37 : rdata = 48'b000100100000101000111111111000000110100000000000;
			// PEs: 40, 43 -> 44
			// srcs: (1727, 31)(3140) 47, (217) 1 --> (3354) 47:PEGB0, ND2, *, PENB
			10'd38 : rdata = 48'b000111110000000001100000010000000000000100000000;
			// PEs: 43, 42 -> 42
			// srcs: (1729, 46)(3) 1, (3353) 47 --> (4137) 47:NM0, PENB, *, PEGB2
			10'd39 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 43, 44 -> 43
			// srcs: (1736, 62)(1002) 2, (4138) 47 --> (4922) -45:NW2, PEGB4, -, NW2
			10'd40 : rdata = 48'b000100100000001011100001000000000100100000000000;
			// PEs: 40, 43 -> 44
			// srcs: (1809, 32)(3140) 47, (299) 1 --> (3436) 47:PEGB0, ND3, *, PENB
			10'd41 : rdata = 48'b000111110000000001100000011000000000000100000000;
			// PEs: 43, 42 -> 42
			// srcs: (1811, 47)(3) 1, (3435) -141 --> (4219) -141:NM0, PENB, *, PEGB2
			10'd42 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 43, 44 -> 43
			// srcs: (1818, 63)(1084) -1, (4220) 47 --> (5004) -48:NW3, PEGB4, -, NW3
			10'd43 : rdata = 48'b000100100000001111100001000000000100110000000000;
			// PEs: 40, 43 -> 
			// srcs: (1875, 33)(3140) 47, (365) 1 --> (3502) 47:PEGB0, ND11, *, 
			10'd44 : rdata = 48'b000111110000000001100001011000000000000000000000;
			// PEs: 43, 43 -> 
			// srcs: (1878, 48)(3) 1, (3502) 47 --> (4286) 47:NM0, ALU, *, 
			10'd45 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 43, 43 -> 43
			// srcs: (1881, 64)(1150) -2, (4286) 47 --> (5070) -49:NW11, ALU, -, NW11
			10'd46 : rdata = 48'b000100100000101100111111111000000110110000000000;
			// PEs: 40, 43 -> 43
			// srcs: (1889, 34)(3140) 47, (379) 2 --> (3516) 94:PEGB0, ND4, *, NI0
			10'd47 : rdata = 48'b000111110000000001100000100100000000000000000000;
			// PEs: 43, 42 -> 42
			// srcs: (1891, 49)(3) 1, (3515) 47 --> (4299) 47:NM0, PENB, *, PEGB2
			10'd48 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 43, 43 -> 
			// srcs: (1892, 50)(3) 1, (3516) 94 --> (4300) 94:NM0, NI0, *, 
			10'd49 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 43, 43 -> 43
			// srcs: (1895, 65)(1164) -1, (4300) 94 --> (5084) -95:NW4, ALU, -, NW4
			10'd50 : rdata = 48'b000100100000010000111111111000000101000000000000;
			// PEs: 40, 43 -> 44
			// srcs: (1969, 35)(3140) 47, (459) 2 --> (3596) 94:PEGB0, ND5, *, PENB
			10'd51 : rdata = 48'b000111110000000001100000101000000000000100000000;
			// PEs: 43, 42 -> 42
			// srcs: (1971, 51)(3) 1, (3595) -141 --> (4379) -141:NM0, PENB, *, PEGB2
			10'd52 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 43, 44 -> 43
			// srcs: (1978, 66)(1244) 0, (4380) 94 --> (5164) -94:NW5, PEGB4, -, NW5
			10'd53 : rdata = 48'b000100100000010111100001000000000101010000000000;
			// PEs: 40, 43 -> 44
			// srcs: (2051, 36)(3140) 47, (541) -2 --> (3678) -94:PEGB0, ND6, *, PENB
			10'd54 : rdata = 48'b000111110000000001100000110000000000000100000000;
			// PEs: 43, 42 -> 42
			// srcs: (2053, 52)(3) 1, (3677) -94 --> (4461) -94:NM0, PENB, *, PEGB2
			10'd55 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 43, 42 -> 42
			// srcs: (2055, 53)(3) 1, (3679) 0 --> (4463) 0:NM0, PENB, *, PEGB2
			10'd56 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 40, 43 -> 43
			// srcs: (2059, 37)(3140) 47, (549) 2 --> (3686) 94:PEGB0, ND12, *, NI0
			10'd57 : rdata = 48'b000111110000000001100001100100000000000000000000;
			// PEs: 43, 44 -> 43
			// srcs: (2060, 67)(1326) -3, (4462) -94 --> (5246) 91:NW6, PEGB4, -, NW6
			10'd58 : rdata = 48'b000100100000011011100001000000000101100000000000;
			// PEs: 43, 43 -> 
			// srcs: (2062, 54)(3) 1, (3686) 94 --> (4470) 94:NM0, NI0, *, 
			10'd59 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 43, 43 -> 43
			// srcs: (2065, 68)(1334) -1, (4470) 94 --> (5254) -95:NW12, ALU, -, NW12
			10'd60 : rdata = 48'b000100100000110000111111111000000111000000000000;
			// PEs: 40, 43 -> 44
			// srcs: (2131, 38)(3140) 47, (621) -1 --> (3758) -47:PEGB0, ND7, *, PENB
			10'd61 : rdata = 48'b000111110000000001100000111000000000000100000000;
			// PEs: 43, 42 -> 42
			// srcs: (2133, 55)(3) 1, (3757) -47 --> (4541) -47:NM0, PENB, *, PEGB2
			10'd62 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 43, 44 -> 43
			// srcs: (2140, 69)(1406) 2, (4542) -47 --> (5326) 49:NW7, PEGB4, -, NW7
			10'd63 : rdata = 48'b000100100000011111100001000000000101110000000000;
			// PEs: 40, 43 -> 44
			// srcs: (2211, 39)(3140) 47, (701) -3 --> (3838) -141:PEGB0, ND8, *, PENB
			10'd64 : rdata = 48'b000111110000000001100001000000000000000100000000;
			// PEs: 43, 42 -> 42
			// srcs: (2213, 56)(3) 1, (3837) -141 --> (4621) -141:NM0, PENB, *, PEGB2
			10'd65 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 43, 44 -> 43
			// srcs: (2220, 70)(1486) 0, (4622) -141 --> (5406) 141:NW8, PEGB4, -, NW8
			10'd66 : rdata = 48'b000100100000100011100001000000000110000000000000;
			// PEs: 40, 43 -> 
			// srcs: (2239, 40)(3140) 47, (729) 0 --> (3866) 0:PEGB0, ND13, *, 
			10'd67 : rdata = 48'b000111110000000001100001101000000000000000000000;
			// PEs: 43, 43 -> 
			// srcs: (2242, 57)(3) 1, (3866) 0 --> (4650) 0:NM0, ALU, *, 
			10'd68 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 43, 43 -> 43
			// srcs: (2245, 71)(1514) -2, (4650) 0 --> (5434) -2:NW13, ALU, -, NW13
			10'd69 : rdata = 48'b000100100000110100111111111000000111010000000000;
			// PEs: 40, 43 -> 44
			// srcs: (2293, 41)(3140) 47, (783) -3 --> (3920) -141:PEGB0, ND9, *, PENB
			10'd70 : rdata = 48'b000111110000000001100001001000000000000100000000;
			// PEs: 43, 42 -> 42
			// srcs: (2295, 58)(3) 1, (3919) 47 --> (4703) 47:NM0, PENB, *, PEGB2
			10'd71 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 43, 44 -> 43
			// srcs: (2302, 72)(1568) -3, (4704) -141 --> (5488) 138:NW9, PEGB4, -, NW9
			10'd72 : rdata = 48'b000100100000100111100001000000000110010000000000;
			default : rdata = 48'b000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 44) begin
	always @(*) begin
		case(address)
			// PEs: 44, 44 -> 40
			// srcs: (1, 0)(57) 0, (842) -2 --> (1626) 0:ND0, NW0, *, PEGB0
			10'd0 : rdata = 48'b000110110000000001000000000000000000000010000000;
			// PEs: 44, 44 -> 40
			// srcs: (2, 1)(139) 0, (924) 1 --> (1708) 0:ND1, NW1, *, PEGB0
			10'd1 : rdata = 48'b000110110000000101000000001000000000000010000000;
			// PEs: 44, 44 -> 40
			// srcs: (3, 2)(219) -1, (1004) -3 --> (1788) 3:ND2, NW2, *, PEGB0
			10'd2 : rdata = 48'b000110110000001001000000010000000000000010000000;
			// PEs: 44, 44 -> 44
			// srcs: (4, 3)(300) 0, (1085) -3 --> (1869) 0:ND3, NW3, *, NI0
			10'd3 : rdata = 48'b000110110000001101000000011100000000000000000000;
			// PEs: 44, 44 -> 40
			// srcs: (5, 4)(381) -3, (1166) -3 --> (1950) 9:ND4, NW4, *, PEGB0
			10'd4 : rdata = 48'b000110110000010001000000100000000000000010000000;
			// PEs: 44, 44 -> 40
			// srcs: (6, 5)(461) 1, (1246) -1 --> (2030) -1:ND5, NW5, *, PEGB0
			10'd5 : rdata = 48'b000110110000010101000000101000000000000010000000;
			// PEs: 44, 44 -> 44
			// srcs: (7, 6)(543) -3, (1328) -3 --> (2112) 9:ND6, NW6, *, NI1
			10'd6 : rdata = 48'b000110110000011001000000110100001000000000000000;
			// PEs: 44, 44 -> 40
			// srcs: (8, 7)(623) 1, (1408) -3 --> (2192) -3:ND7, NW7, *, PEGB0
			10'd7 : rdata = 48'b000110110000011101000000111000000000000010000000;
			// PEs: 44, 44 -> 43
			// srcs: (9, 8)(703) -2, (1488) 2 --> (2272) -4:ND8, NW8, *, PEGB3
			10'd8 : rdata = 48'b000110110000100001000001000000000000000010110000;
			// PEs: 44, 44 -> 46
			// srcs: (10, 9)(785) -2, (1570) 1 --> (2354) -2:ND9, NW9, *, PEGB6
			10'd9 : rdata = 48'b000110110000100101000001001000000000000011100000;
			// PEs: 44, 44 -> 40
			// srcs: (11, 10)(184) -2, (969) 2 --> (1753) -4:ND10, NW10, *, PEGB0
			10'd10 : rdata = 48'b000110110000101001000001010000000000000010000000;
			// PEs: 44, 44 -> 47
			// srcs: (12, 11)(368) -3, (1153) -2 --> (1937) 6:ND11, NW11, *, PEGB7
			10'd11 : rdata = 48'b000110110000101101000001011000000000000011110000;
			// PEs: 44, 44 -> 44
			// srcs: (13, 12)(552) -1, (1337) 0 --> (2121) 0:ND12, NW12, *, NI2
			10'd12 : rdata = 48'b000110110000110001000001100100010000000000000000;
			// PEs: 44, 44 -> 44
			// srcs: (14, 13)(732) -1, (1517) 0 --> (2301) 0:ND13, NW13, *, NI3
			10'd13 : rdata = 48'b000110110000110101000001101100011000000000000000;
			// PEs: 47 -> 
			// srcs: (15, 18)(2276) -1 --> (2276) -1:PEGB7, pass, 
			10'd14 : rdata = 48'b110001110000111000000000000000000000000000000000;
			// PEs: 46, 44 -> 44
			// srcs: (17, 19)(2275) -1, (2276) -1 --> (3054) -2:PEGB6, ALU, +, NI4
			10'd15 : rdata = 48'b000011110000110000111111111100100000000000000000;
			// PEs: 40 -> 
			// srcs: (24, 14)(1700) -2 --> (1700) -2:PEGB0, pass, 
			10'd16 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 40, 44 -> 41
			// srcs: (33, 15)(1699) 0, (1700) -2 --> (2480) -2:PEGB0, ALU, +, PEGB1
			10'd17 : rdata = 48'b000011110000000000111111111000000000000010010000;
			// PEs: 40 -> 
			// srcs: (55, 16)(1862) 0 --> (1862) 0:PEGB0, pass, 
			10'd18 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 40, 44 -> 44
			// srcs: (64, 17)(1861) 1, (1862) 0 --> (2640) 1:PEGB0, ALU, +, NI5
			10'd19 : rdata = 48'b000011110000000000111111111100101000000000000000;
			// PEs: 44 -> 40
			// srcs: (116, 20)(1869) 0 --> (1869) 0:NI0, pass, PEGB0
			10'd20 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 44 -> 40
			// srcs: (126, 22)(2640) 1 --> (2640) 1:NI5, pass, PEGB0
			10'd21 : rdata = 48'b110001010000010100000000000000000000000010000000;
			// PEs: 44 -> 40
			// srcs: (133, 21)(2112) 9 --> (2112) 9:NI1, pass, PEGB0
			10'd22 : rdata = 48'b110001010000000100000000000000000000000010000000;
			// PEs: 44 -> 40
			// srcs: (134, 27)(2301) 0 --> (2301) 0:NI3, pass, PEGB0
			10'd23 : rdata = 48'b110001010000001100000000000000000000000010000000;
			// PEs: 44 -> 40
			// srcs: (139, 25)(2121) 0 --> (2121) 0:NI2, pass, PEGB0
			10'd24 : rdata = 48'b110001010000001000000000000000000000000010000000;
			// PEs: 40 -> 
			// srcs: (612, 23)(2099) 0 --> (2099) 0:PEGB0, pass, 
			10'd25 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 41, 44 -> 44
			// srcs: (614, 24)(2876) 6, (2099) 0 --> (2877) 6:PEGB1, ALU, +, NI0
			10'd26 : rdata = 48'b000011110000001000111111111100000000000000000000;
			// PEs: 44 -> 41
			// srcs: (696, 26)(3054) -2 --> (3054) -2:NI4, pass, PEGB1
			10'd27 : rdata = 48'b110001010000010000000000000000000000000010010000;
			// PEs: 44 -> 41
			// srcs: (753, 28)(2877) 6 --> (2877) 6:NI0, pass, PEGB1
			10'd28 : rdata = 48'b110001010000000000000000000000000000000010010000;
			// PEs: 40, 44 -> 45
			// srcs: (1567, 29)(3140) 47, (57) 0 --> (3194) 0:PEGB0, ND0, *, PENB
			10'd29 : rdata = 48'b000111110000000001100000000000000000000100000000;
			// PEs: 44, 45 -> 44
			// srcs: (1576, 59)(842) -2, (3978) 0 --> (4762) -2:NW0, PEGB5, -, NW0
			10'd30 : rdata = 48'b000100100000000011100001010000000100000000000000;
			// PEs: 40, 44 -> 44
			// srcs: (1649, 30)(3140) 47, (139) 0 --> (3276) 0:PEGB0, ND1, *, NI0
			10'd31 : rdata = 48'b000111110000000001100000001100000000000000000000;
			// PEs: 44, 43 -> 43
			// srcs: (1650, 43)(3) 1, (3274) 94 --> (4058) 94:NM0, PENB, *, PEGB3
			10'd32 : rdata = 48'b000111000000000011011111110000000000000010110000;
			// PEs: 44, 44 -> 
			// srcs: (1652, 44)(3) 1, (3276) 0 --> (4060) 0:NM0, NI0, *, 
			10'd33 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 44, 44 -> 44
			// srcs: (1655, 60)(924) 1, (4060) 0 --> (4844) 1:NW1, ALU, -, NW1
			10'd34 : rdata = 48'b000100100000000100111111111000000100010000000000;
			// PEs: 40, 44 -> 
			// srcs: (1694, 31)(3140) 47, (184) -2 --> (3321) -94:PEGB0, ND10, *, 
			10'd35 : rdata = 48'b000111110000000001100001010000000000000000000000;
			// PEs: 44, 44 -> 
			// srcs: (1697, 45)(3) 1, (3321) -94 --> (4105) -94:NM0, ALU, *, 
			10'd36 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 44, 44 -> 44
			// srcs: (1700, 61)(969) 2, (4105) -94 --> (4889) 96:NW10, ALU, -, NW10
			10'd37 : rdata = 48'b000100100000101000111111111000000110100000000000;
			// PEs: 40, 44 -> 45
			// srcs: (1729, 32)(3140) 47, (219) -1 --> (3356) -47:PEGB0, ND2, *, PENB
			10'd38 : rdata = 48'b000111110000000001100000010000000000000100000000;
			// PEs: 44, 43 -> 43
			// srcs: (1730, 46)(3) 1, (3354) 47 --> (4138) 47:NM0, PENB, *, PEGB3
			10'd39 : rdata = 48'b000111000000000011011111110000000000000010110000;
			// PEs: 44, 45 -> 44
			// srcs: (1738, 62)(1004) -3, (4140) -47 --> (4924) 44:NW2, PEGB5, -, NW2
			10'd40 : rdata = 48'b000100100000001011100001010000000100100000000000;
			// PEs: 40, 44 -> 44
			// srcs: (1810, 33)(3140) 47, (300) 0 --> (3437) 0:PEGB0, ND3, *, NI0
			10'd41 : rdata = 48'b000111110000000001100000011100000000000000000000;
			// PEs: 44, 43 -> 43
			// srcs: (1812, 47)(3) 1, (3436) 47 --> (4220) 47:NM0, PENB, *, PEGB3
			10'd42 : rdata = 48'b000111000000000011011111110000000000000010110000;
			// PEs: 44, 44 -> 
			// srcs: (1813, 48)(3) 1, (3437) 0 --> (4221) 0:NM0, NI0, *, 
			10'd43 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 44, 44 -> 44
			// srcs: (1816, 63)(1085) -3, (4221) 0 --> (5005) -3:NW3, ALU, -, NW3
			10'd44 : rdata = 48'b000100100000001100111111111000000100110000000000;
			// PEs: 40, 44 -> 
			// srcs: (1878, 34)(3140) 47, (368) -3 --> (3505) -141:PEGB0, ND11, *, 
			10'd45 : rdata = 48'b000111110000000001100001011000000000000000000000;
			// PEs: 44, 44 -> 
			// srcs: (1881, 49)(3) 1, (3505) -141 --> (4289) -141:NM0, ALU, *, 
			10'd46 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 44, 44 -> 44
			// srcs: (1884, 64)(1153) -2, (4289) -141 --> (5073) 139:NW11, ALU, -, NW11
			10'd47 : rdata = 48'b000100100000101100111111111000000110110000000000;
			// PEs: 40, 44 -> 
			// srcs: (1891, 35)(3140) 47, (381) -3 --> (3518) -141:PEGB0, ND4, *, 
			10'd48 : rdata = 48'b000111110000000001100000100000000000000000000000;
			// PEs: 44, 44 -> 
			// srcs: (1894, 50)(3) 1, (3518) -141 --> (4302) -141:NM0, ALU, *, 
			10'd49 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 44, 44 -> 44
			// srcs: (1897, 65)(1166) -3, (4302) -141 --> (5086) 138:NW4, ALU, -, NW4
			10'd50 : rdata = 48'b000100100000010000111111111000000101000000000000;
			// PEs: 40, 44 -> 45
			// srcs: (1971, 36)(3140) 47, (461) 1 --> (3598) 47:PEGB0, ND5, *, PENB
			10'd51 : rdata = 48'b000111110000000001100000101000000000000100000000;
			// PEs: 44, 43 -> 43
			// srcs: (1972, 51)(3) 1, (3596) 94 --> (4380) 94:NM0, PENB, *, PEGB3
			10'd52 : rdata = 48'b000111000000000011011111110000000000000010110000;
			// PEs: 44, 45 -> 44
			// srcs: (1980, 66)(1246) -1, (4382) 47 --> (5166) -48:NW5, PEGB5, -, NW5
			10'd53 : rdata = 48'b000100100000010111100001010000000101010000000000;
			// PEs: 40, 44 -> 45
			// srcs: (2053, 37)(3140) 47, (543) -3 --> (3680) -141:PEGB0, ND6, *, PENB
			10'd54 : rdata = 48'b000111110000000001100000110000000000000100000000;
			// PEs: 44, 43 -> 43
			// srcs: (2054, 52)(3) 1, (3678) -94 --> (4462) -94:NM0, PENB, *, PEGB3
			10'd55 : rdata = 48'b000111000000000011011111110000000000000010110000;
			// PEs: 40, 44 -> 44
			// srcs: (2062, 38)(3140) 47, (552) -1 --> (3689) -47:PEGB0, ND12, *, NI0
			10'd56 : rdata = 48'b000111110000000001100001100100000000000000000000;
			// PEs: 44, 45 -> 44
			// srcs: (2063, 67)(1328) -3, (4464) -141 --> (5248) 138:NW6, PEGB5, -, NW6
			10'd57 : rdata = 48'b000100100000011011100001010000000101100000000000;
			// PEs: 44, 44 -> 
			// srcs: (2065, 53)(3) 1, (3689) -47 --> (4473) -47:NM0, NI0, *, 
			10'd58 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 44, 44 -> 44
			// srcs: (2068, 68)(1337) 0, (4473) -47 --> (5257) 47:NW12, ALU, -, NW12
			10'd59 : rdata = 48'b000100100000110000111111111000000111000000000000;
			// PEs: 40, 44 -> 45
			// srcs: (2133, 39)(3140) 47, (623) 1 --> (3760) 47:PEGB0, ND7, *, PENB
			10'd60 : rdata = 48'b000111110000000001100000111000000000000100000000;
			// PEs: 44, 43 -> 43
			// srcs: (2134, 54)(3) 1, (3758) -47 --> (4542) -47:NM0, PENB, *, PEGB3
			10'd61 : rdata = 48'b000111000000000011011111110000000000000010110000;
			// PEs: 44, 45 -> 44
			// srcs: (2142, 69)(1408) -3, (4544) 47 --> (5328) -50:NW7, PEGB5, -, NW7
			10'd62 : rdata = 48'b000100100000011111100001010000000101110000000000;
			// PEs: 40, 44 -> 44
			// srcs: (2213, 40)(3140) 47, (703) -2 --> (3840) -94:PEGB0, ND8, *, NI0
			10'd63 : rdata = 48'b000111110000000001100001000100000000000000000000;
			// PEs: 44, 43 -> 43
			// srcs: (2214, 55)(3) 1, (3838) -141 --> (4622) -141:NM0, PENB, *, PEGB3
			10'd64 : rdata = 48'b000111000000000011011111110000000000000010110000;
			// PEs: 44, 44 -> 
			// srcs: (2216, 56)(3) 1, (3840) -94 --> (4624) -94:NM0, NI0, *, 
			10'd65 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 44, 44 -> 44
			// srcs: (2219, 70)(1488) 2, (4624) -94 --> (5408) 96:NW8, ALU, -, NW8
			10'd66 : rdata = 48'b000100100000100000111111111000000110000000000000;
			// PEs: 40, 44 -> 
			// srcs: (2242, 41)(3140) 47, (732) -1 --> (3869) -47:PEGB0, ND13, *, 
			10'd67 : rdata = 48'b000111110000000001100001101000000000000000000000;
			// PEs: 44, 44 -> 
			// srcs: (2245, 57)(3) 1, (3869) -47 --> (4653) -47:NM0, ALU, *, 
			10'd68 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 44, 44 -> 44
			// srcs: (2248, 71)(1517) 0, (4653) -47 --> (5437) 47:NW13, ALU, -, NW13
			10'd69 : rdata = 48'b000100100000110100111111111000000111010000000000;
			// PEs: 40, 44 -> 45
			// srcs: (2295, 42)(3140) 47, (785) -2 --> (3922) -94:PEGB0, ND9, *, PENB
			10'd70 : rdata = 48'b000111110000000001100001001000000000000100000000;
			// PEs: 44, 43 -> 43
			// srcs: (2296, 58)(3) 1, (3920) -141 --> (4704) -141:NM0, PENB, *, PEGB3
			10'd71 : rdata = 48'b000111000000000011011111110000000000000010110000;
			// PEs: 44, 45 -> 44
			// srcs: (2304, 72)(1570) 1, (4706) -94 --> (5490) 95:NW9, PEGB5, -, NW9
			10'd72 : rdata = 48'b000100100000100111100001010000000110010000000000;
			default : rdata = 48'b000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 45) begin
	always @(*) begin
		case(address)
			// PEs: 45, 45 -> 40
			// srcs: (1, 0)(58) -3, (843) -2 --> (1627) 6:ND0, NW0, *, PEGB0
			10'd0 : rdata = 48'b000110110000000001000000000000000000000010000000;
			// PEs: 45, 45 -> 40
			// srcs: (2, 1)(140) 0, (925) -3 --> (1709) 0:ND1, NW1, *, PEGB0
			10'd1 : rdata = 48'b000110110000000101000000001000000000000010000000;
			// PEs: 45, 45 -> 40
			// srcs: (3, 2)(220) 2, (1005) 2 --> (1789) 4:ND2, NW2, *, PEGB0
			10'd2 : rdata = 48'b000110110000001001000000010000000000000010000000;
			// PEs: 45, 45 -> 45
			// srcs: (4, 3)(301) 0, (1086) 0 --> (1870) 0:ND3, NW3, *, NI0
			10'd3 : rdata = 48'b000110110000001101000000011100000000000000000000;
			// PEs: 45, 45 -> 40
			// srcs: (5, 4)(382) -2, (1167) -3 --> (1951) 6:ND4, NW4, *, PEGB0
			10'd4 : rdata = 48'b000110110000010001000000100000000000000010000000;
			// PEs: 45, 45 -> 40
			// srcs: (6, 5)(462) -1, (1247) 2 --> (2031) -2:ND5, NW5, *, PEGB0
			10'd5 : rdata = 48'b000110110000010101000000101000000000000010000000;
			// PEs: 45, 45 -> 45
			// srcs: (7, 6)(544) 1, (1329) -1 --> (2113) -1:ND6, NW6, *, NI1
			10'd6 : rdata = 48'b000110110000011001000000110100001000000000000000;
			// PEs: 45, 45 -> 40
			// srcs: (8, 7)(624) 2, (1409) -3 --> (2193) -6:ND7, NW7, *, PEGB0
			10'd7 : rdata = 48'b000110110000011101000000111000000000000010000000;
			// PEs: 45, 45 -> 43
			// srcs: (9, 8)(704) -1, (1489) 2 --> (2273) -2:ND8, NW8, *, PEGB3
			10'd8 : rdata = 48'b000110110000100001000001000000000000000010110000;
			// PEs: 45, 45 -> 46
			// srcs: (10, 9)(786) 0, (1571) 1 --> (2355) 0:ND9, NW9, *, PENB
			10'd9 : rdata = 48'b000110110000100101000001001000000000000100000000;
			// PEs: 45, 45 -> 45
			// srcs: (11, 10)(187) 2, (972) -1 --> (1756) -2:ND10, NW10, *, NI2
			10'd10 : rdata = 48'b000110110000101001000001010100010000000000000000;
			// PEs: 45, 45 -> 46
			// srcs: (12, 11)(371) 1, (1156) -1 --> (1940) -1:ND11, NW11, *, PENB
			10'd11 : rdata = 48'b000110110000101101000001011000000000000100000000;
			// PEs: 45, 45 -> 40
			// srcs: (13, 12)(555) -3, (1340) 1 --> (2124) -3:ND12, NW12, *, PEGB0
			10'd12 : rdata = 48'b000110110000110001000001100000000000000010000000;
			// PEs: 45, 45 -> 45
			// srcs: (14, 13)(735) -1, (1520) -1 --> (2304) 1:ND13, NW13, *, NI3
			10'd13 : rdata = 48'b000110110000110101000001101100011000000000000000;
			// PEs: 43 -> 
			// srcs: (15, 18)(2352) 9 --> (2352) 9:PEGB3, pass, 
			10'd14 : rdata = 48'b110001110000011000000000000000000000000000000000;
			// PEs: 42, 45 -> 45
			// srcs: (18, 19)(2351) -1, (2352) 9 --> (3128) 8:PEGB2, ALU, +, NI4
			10'd15 : rdata = 48'b000011110000010000111111111100100000000000000000;
			// PEs: 40 -> 
			// srcs: (30, 14)(1774) 1 --> (1774) 1:PEGB0, pass, 
			10'd16 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 40, 45 -> 45
			// srcs: (39, 15)(1773) 0, (1774) 1 --> (2555) 1:PEGB0, ALU, +, NI5
			10'd17 : rdata = 48'b000011110000000000111111111100101000000000000000;
			// PEs: 40 -> 
			// srcs: (86, 16)(1944) 4 --> (1944) 4:PEGB0, pass, 
			10'd18 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 45, 41 -> 47
			// srcs: (88, 17)(1944) 4, (1945) -2 --> (2723) 2:ALU, PEGB1, +, PEGB7
			10'd19 : rdata = 48'b000010011111111111100000010000000000000011110000;
			// PEs: 45 -> 40
			// srcs: (125, 20)(1870) 0 --> (1870) 0:NI0, pass, PEGB0
			10'd20 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 45 -> 40
			// srcs: (141, 21)(2113) -1 --> (2113) -1:NI1, pass, PEGB0
			10'd21 : rdata = 48'b110001010000000100000000000000000000000010000000;
			// PEs: 45 -> 40
			// srcs: (142, 24)(2304) 1 --> (2304) 1:NI3, pass, PEGB0
			10'd22 : rdata = 48'b110001010000001100000000000000000000000010000000;
			// PEs: 45 -> 40
			// srcs: (143, 25)(3128) 8 --> (3128) 8:NI4, pass, PEGB0
			10'd23 : rdata = 48'b110001010000010000000000000000000000000010000000;
			// PEs: 45 -> 40
			// srcs: (170, 22)(1756) -2 --> (1756) -2:NI2, pass, PEGB0
			10'd24 : rdata = 48'b110001010000001000000000000000000000000010000000;
			// PEs: 45 -> 40
			// srcs: (178, 23)(2555) 1 --> (2555) 1:NI5, pass, PEGB0
			10'd25 : rdata = 48'b110001010000010100000000000000000000000010000000;
			// PEs: 40 -> 
			// srcs: (781, 26)(2702) 13 --> (2702) 13:PEGB0, pass, 
			10'd26 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 45, 46 -> 46
			// srcs: (783, 27)(2702) 13, (2707) -11 --> (2708) 2:ALU, PEGB6, +, PENB
			10'd27 : rdata = 48'b000010011111111111100001100000000000000100000000;
			// PEs: 40, 45 -> 45
			// srcs: (1568, 28)(3140) 47, (58) -3 --> (3195) -141:PEGB0, ND0, *, NI0
			10'd28 : rdata = 48'b000111110000000001100000000100000000000000000000;
			// PEs: 45, 44 -> 44
			// srcs: (1570, 42)(3) 1, (3194) 0 --> (3978) 0:NM0, PENB, *, PEGB4
			10'd29 : rdata = 48'b000111000000000011011111110000000000000011000000;
			// PEs: 45, 45 -> 
			// srcs: (1571, 43)(3) 1, (3195) -141 --> (3979) -141:NM0, NI0, *, 
			10'd30 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 45, 45 -> 45
			// srcs: (1574, 59)(843) -2, (3979) -141 --> (4763) 139:NW0, ALU, -, NW0
			10'd31 : rdata = 48'b000100100000000000111111111000000100000000000000;
			// PEs: 40, 45 -> 
			// srcs: (1650, 29)(3140) 47, (140) 0 --> (3277) 0:PEGB0, ND1, *, 
			10'd32 : rdata = 48'b000111110000000001100000001000000000000000000000;
			// PEs: 45, 45 -> 
			// srcs: (1653, 44)(3) 1, (3277) 0 --> (4061) 0:NM0, ALU, *, 
			10'd33 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 45, 45 -> 45
			// srcs: (1656, 60)(925) -3, (4061) 0 --> (4845) -3:NW1, ALU, -, NW1
			10'd34 : rdata = 48'b000100100000000100111111111000000100010000000000;
			// PEs: 40, 45 -> 
			// srcs: (1697, 30)(3140) 47, (187) 2 --> (3324) 94:PEGB0, ND10, *, 
			10'd35 : rdata = 48'b000111110000000001100001010000000000000000000000;
			// PEs: 45, 45 -> 
			// srcs: (1700, 45)(3) 1, (3324) 94 --> (4108) 94:NM0, ALU, *, 
			10'd36 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 45, 45 -> 45
			// srcs: (1703, 61)(972) -1, (4108) 94 --> (4892) -95:NW10, ALU, -, NW10
			10'd37 : rdata = 48'b000100100000101000111111111000000110100000000000;
			// PEs: 40, 45 -> 45
			// srcs: (1730, 31)(3140) 47, (220) 2 --> (3357) 94:PEGB0, ND2, *, NI0
			10'd38 : rdata = 48'b000111110000000001100000010100000000000000000000;
			// PEs: 45, 44 -> 44
			// srcs: (1732, 46)(3) 1, (3356) -47 --> (4140) -47:NM0, PENB, *, PEGB4
			10'd39 : rdata = 48'b000111000000000011011111110000000000000011000000;
			// PEs: 45, 45 -> 
			// srcs: (1733, 47)(3) 1, (3357) 94 --> (4141) 94:NM0, NI0, *, 
			10'd40 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 45, 45 -> 45
			// srcs: (1736, 62)(1005) 2, (4141) 94 --> (4925) -92:NW2, ALU, -, NW2
			10'd41 : rdata = 48'b000100100000001000111111111000000100100000000000;
			// PEs: 40, 45 -> 
			// srcs: (1811, 32)(3140) 47, (301) 0 --> (3438) 0:PEGB0, ND3, *, 
			10'd42 : rdata = 48'b000111110000000001100000011000000000000000000000;
			// PEs: 45, 45 -> 
			// srcs: (1814, 48)(3) 1, (3438) 0 --> (4222) 0:NM0, ALU, *, 
			10'd43 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 45, 45 -> 45
			// srcs: (1817, 63)(1086) 0, (4222) 0 --> (5006) 0:NW3, ALU, -, NW3
			10'd44 : rdata = 48'b000100100000001100111111111000000100110000000000;
			// PEs: 40, 45 -> 
			// srcs: (1881, 33)(3140) 47, (371) 1 --> (3508) 47:PEGB0, ND11, *, 
			10'd45 : rdata = 48'b000111110000000001100001011000000000000000000000;
			// PEs: 45, 45 -> 
			// srcs: (1884, 49)(3) 1, (3508) 47 --> (4292) 47:NM0, ALU, *, 
			10'd46 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 45, 45 -> 45
			// srcs: (1887, 64)(1156) -1, (4292) 47 --> (5076) -48:NW11, ALU, -, NW11
			10'd47 : rdata = 48'b000100100000101100111111111000000110110000000000;
			// PEs: 40, 45 -> 
			// srcs: (1892, 34)(3140) 47, (382) -2 --> (3519) -94:PEGB0, ND4, *, 
			10'd48 : rdata = 48'b000111110000000001100000100000000000000000000000;
			// PEs: 45, 45 -> 
			// srcs: (1895, 50)(3) 1, (3519) -94 --> (4303) -94:NM0, ALU, *, 
			10'd49 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 45, 45 -> 45
			// srcs: (1898, 65)(1167) -3, (4303) -94 --> (5087) 91:NW4, ALU, -, NW4
			10'd50 : rdata = 48'b000100100000010000111111111000000101000000000000;
			// PEs: 40, 45 -> 46
			// srcs: (1972, 35)(3140) 47, (462) -1 --> (3599) -47:PEGB0, ND5, *, PENB
			10'd51 : rdata = 48'b000111110000000001100000101000000000000100000000;
			// PEs: 45, 44 -> 44
			// srcs: (1974, 51)(3) 1, (3598) 47 --> (4382) 47:NM0, PENB, *, PEGB4
			10'd52 : rdata = 48'b000111000000000011011111110000000000000011000000;
			// PEs: 45, 46 -> 45
			// srcs: (1981, 66)(1247) 2, (4383) -47 --> (5167) 49:NW5, PEGB6, -, NW5
			10'd53 : rdata = 48'b000100100000010111100001100000000101010000000000;
			// PEs: 40, 45 -> 46
			// srcs: (2054, 36)(3140) 47, (544) 1 --> (3681) 47:PEGB0, ND6, *, PENB
			10'd54 : rdata = 48'b000111110000000001100000110000000000000100000000;
			// PEs: 45, 44 -> 44
			// srcs: (2056, 52)(3) 1, (3680) -141 --> (4464) -141:NM0, PENB, *, PEGB4
			10'd55 : rdata = 48'b000111000000000011011111110000000000000011000000;
			// PEs: 45, 46 -> 45
			// srcs: (2063, 67)(1329) -1, (4465) 47 --> (5249) -48:NW6, PEGB6, -, NW6
			10'd56 : rdata = 48'b000100100000011011100001100000000101100000000000;
			// PEs: 40, 45 -> 
			// srcs: (2065, 37)(3140) 47, (555) -3 --> (3692) -141:PEGB0, ND12, *, 
			10'd57 : rdata = 48'b000111110000000001100001100000000000000000000000;
			// PEs: 45, 45 -> 
			// srcs: (2068, 53)(3) 1, (3692) -141 --> (4476) -141:NM0, ALU, *, 
			10'd58 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 45, 45 -> 45
			// srcs: (2071, 68)(1340) 1, (4476) -141 --> (5260) 142:NW12, ALU, -, NW12
			10'd59 : rdata = 48'b000100100000110000111111111000000111000000000000;
			// PEs: 40, 45 -> 45
			// srcs: (2134, 38)(3140) 47, (624) 2 --> (3761) 94:PEGB0, ND7, *, NI0
			10'd60 : rdata = 48'b000111110000000001100000111100000000000000000000;
			// PEs: 45, 44 -> 44
			// srcs: (2136, 54)(3) 1, (3760) 47 --> (4544) 47:NM0, PENB, *, PEGB4
			10'd61 : rdata = 48'b000111000000000011011111110000000000000011000000;
			// PEs: 45, 45 -> 
			// srcs: (2137, 55)(3) 1, (3761) 94 --> (4545) 94:NM0, NI0, *, 
			10'd62 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 45, 45 -> 45
			// srcs: (2140, 69)(1409) -3, (4545) 94 --> (5329) -97:NW7, ALU, -, NW7
			10'd63 : rdata = 48'b000100100000011100111111111000000101110000000000;
			// PEs: 40, 45 -> 
			// srcs: (2214, 39)(3140) 47, (704) -1 --> (3841) -47:PEGB0, ND8, *, 
			10'd64 : rdata = 48'b000111110000000001100001000000000000000000000000;
			// PEs: 45, 45 -> 
			// srcs: (2217, 56)(3) 1, (3841) -47 --> (4625) -47:NM0, ALU, *, 
			10'd65 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 45, 45 -> 45
			// srcs: (2220, 70)(1489) 2, (4625) -47 --> (5409) 49:NW8, ALU, -, NW8
			10'd66 : rdata = 48'b000100100000100000111111111000000110000000000000;
			// PEs: 40, 45 -> 
			// srcs: (2245, 40)(3140) 47, (735) -1 --> (3872) -47:PEGB0, ND13, *, 
			10'd67 : rdata = 48'b000111110000000001100001101000000000000000000000;
			// PEs: 45, 45 -> 
			// srcs: (2248, 57)(3) 1, (3872) -47 --> (4656) -47:NM0, ALU, *, 
			10'd68 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 45, 45 -> 45
			// srcs: (2251, 71)(1520) -1, (4656) -47 --> (5440) 46:NW13, ALU, -, NW13
			10'd69 : rdata = 48'b000100100000110100111111111000000111010000000000;
			// PEs: 40, 45 -> 46
			// srcs: (2296, 41)(3140) 47, (786) 0 --> (3923) 0:PEGB0, ND9, *, PENB
			10'd70 : rdata = 48'b000111110000000001100001001000000000000100000000;
			// PEs: 45, 44 -> 44
			// srcs: (2298, 58)(3) 1, (3922) -94 --> (4706) -94:NM0, PENB, *, PEGB4
			10'd71 : rdata = 48'b000111000000000011011111110000000000000011000000;
			// PEs: 45, 46 -> 45
			// srcs: (2305, 72)(1571) 1, (4707) 0 --> (5491) 1:NW9, PEGB6, -, NW9
			10'd72 : rdata = 48'b000100100000100111100001100000000110010000000000;
			default : rdata = 48'b000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 46) begin
	always @(*) begin
		case(address)
			// PEs: 46, 46 -> 40
			// srcs: (1, 0)(60) -2, (845) -1 --> (1629) 2:ND0, NW0, *, PEGB0
			10'd0 : rdata = 48'b000110110000000001000000000000000000000010000000;
			// PEs: 46, 46 -> 40
			// srcs: (2, 1)(142) 1, (927) 0 --> (1711) 0:ND1, NW1, *, PEGB0
			10'd1 : rdata = 48'b000110110000000101000000001000000000000010000000;
			// PEs: 46, 46 -> 40
			// srcs: (3, 2)(222) -1, (1007) 0 --> (1791) 0:ND2, NW2, *, PEGB0
			10'd2 : rdata = 48'b000110110000001001000000010000000000000010000000;
			// PEs: 46, 46 -> 40
			// srcs: (4, 3)(302) -1, (1087) 0 --> (1871) 0:ND3, NW3, *, PEGB0
			10'd3 : rdata = 48'b000110110000001101000000011000000000000010000000;
			// PEs: 46, 46 -> 40
			// srcs: (5, 4)(384) -3, (1169) 1 --> (1953) -3:ND4, NW4, *, PEGB0
			10'd4 : rdata = 48'b000110110000010001000000100000000000000010000000;
			// PEs: 46, 46 -> 40
			// srcs: (6, 5)(464) -3, (1249) -3 --> (2033) 9:ND5, NW5, *, PEGB0
			10'd5 : rdata = 48'b000110110000010101000000101000000000000010000000;
			// PEs: 46, 46 -> 46
			// srcs: (7, 6)(545) -2, (1330) -1 --> (2114) 2:ND6, NW6, *, NI0
			10'd6 : rdata = 48'b000110110000011001000000110100000000000000000000;
			// PEs: 46, 46 -> 40
			// srcs: (8, 7)(626) 1, (1411) -2 --> (2195) -2:ND7, NW7, *, PEGB0
			10'd7 : rdata = 48'b000110110000011101000000111000000000000010000000;
			// PEs: 46, 46 -> 44
			// srcs: (9, 8)(706) 1, (1491) -1 --> (2275) -1:ND8, NW8, *, PEGB4
			10'd8 : rdata = 48'b000110110000100001000001000000000000000011000000;
			// PEs: 46, 46 -> 40
			// srcs: (10, 9)(10) -3, (795) 2 --> (1579) -6:ND9, NW9, *, PEGB0
			10'd9 : rdata = 48'b000110110000100101000001001000000000000010000000;
			// PEs: 46, 46 -> 40
			// srcs: (11, 10)(190) -2, (975) -1 --> (1759) 2:ND10, NW10, *, PEGB0
			10'd10 : rdata = 48'b000110110000101001000001010000000000000010000000;
			// PEs: 46, 46 -> 46
			// srcs: (12, 11)(374) 2, (1159) 2 --> (1943) 4:ND11, NW11, *, NI1
			10'd11 : rdata = 48'b000110110000101101000001011100001000000000000000;
			// PEs: 46, 46 -> 40
			// srcs: (13, 12)(558) 2, (1343) -1 --> (2127) -2:ND12, NW12, *, PEGB0
			10'd12 : rdata = 48'b000110110000110001000001100000000000000010000000;
			// PEs: 46, 46 -> 46
			// srcs: (14, 13)(738) 2, (1523) 1 --> (2307) 2:ND13, NW13, *, NI2
			10'd13 : rdata = 48'b000110110000110101000001101100010000000000000000;
			// PEs: 44, 45 -> 41
			// srcs: (16, 18)(2354) -2, (2355) 0 --> (3130) -2:PEGB4, PENB, +, PEGB1
			10'd14 : rdata = 48'b000011110000100011011111110000000000000010010000;
			// PEs: 40 -> 
			// srcs: (34, 14)(1777) 2 --> (1777) 2:PEGB0, pass, 
			10'd15 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 40, 46 -> 46
			// srcs: (43, 15)(1776) 9, (1777) 2 --> (2558) 11:PEGB0, ALU, +, NI3
			10'd16 : rdata = 48'b000011110000000000111111111100011000000000000000;
			// PEs: 40 -> 
			// srcs: (102, 16)(2024) 0 --> (2024) 0:PEGB0, pass, 
			10'd17 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 46, 41 -> 46
			// srcs: (104, 17)(2024) 0, (2025) 0 --> (2804) 0:ALU, PEGB1, +, NI4
			10'd18 : rdata = 48'b000010011111111111100000010100100000000000000000;
			// PEs: 41, 45 -> 47
			// srcs: (105, 21)(2716) -3, (1940) -1 --> (2717) -4:PEGB1, PENB, +, PENB
			10'd19 : rdata = 48'b000011110000001011011111110000000000000100000000;
			// PEs: 41, 46 -> 47
			// srcs: (106, 22)(2721) 2, (1943) 4 --> (2722) 6:PEGB1, NI1, +, PENB
			10'd20 : rdata = 48'b000011110000001010100000001000000000000100000000;
			// PEs: 46 -> 40
			// srcs: (149, 19)(2114) 2 --> (2114) 2:NI0, pass, PEGB0
			10'd21 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 46 -> 40
			// srcs: (186, 20)(2558) 11 --> (2558) 11:NI3, pass, PEGB0
			10'd22 : rdata = 48'b110001010000001100000000000000000000000010000000;
			// PEs: 46 -> 40
			// srcs: (215, 23)(2804) 0 --> (2804) 0:NI4, pass, PEGB0
			10'd23 : rdata = 48'b110001010000010000000000000000000000000010000000;
			// PEs: 46 -> 40
			// srcs: (257, 24)(2307) 2 --> (2307) 2:NI2, pass, PEGB0
			10'd24 : rdata = 48'b110001010000001000000000000000000000000010000000;
			// PEs: 42 -> 
			// srcs: (411, 27)(2713) -7 --> (2713) -7:PEGB2, pass, 
			10'd25 : rdata = 48'b110001110000010000000000000000000000000000000000;
			// PEs: 46, 47 -> 46
			// srcs: (414, 28)(2713) -7, (2718) 3 --> (2719) -4:ALU, PEGB7, +, NI0
			10'd26 : rdata = 48'b000010011111111111100001110100000000000000000000;
			// PEs: 40 -> 
			// srcs: (732, 25)(2704) -6 --> (2704) -6:PEGB0, pass, 
			10'd27 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 46, 41 -> 45
			// srcs: (734, 26)(2704) -6, (2706) -5 --> (2707) -11:ALU, PEGB1, +, PEGB5
			10'd28 : rdata = 48'b000010011111111111100000010000000000000011010000;
			// PEs: 45, 46 -> 40
			// srcs: (786, 29)(2708) 2, (2719) -4 --> (2720) -2:PENB, NI0, +, PEGB0
			10'd29 : rdata = 48'b000011101111111010100000000000000000000010000000;
			// PEs: 40, 46 -> 
			// srcs: (1521, 30)(3140) 47, (10) -3 --> (3147) -141:PEGB0, ND9, *, 
			10'd30 : rdata = 48'b000111110000000001100001001000000000000000000000;
			// PEs: 46, 46 -> 
			// srcs: (1524, 44)(3) 1, (3147) -141 --> (3931) -141:NM0, ALU, *, 
			10'd31 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 46, 46 -> 46
			// srcs: (1527, 59)(795) 2, (3931) -141 --> (4715) 143:NW9, ALU, -, NW9
			10'd32 : rdata = 48'b000100100000100100111111111000000110010000000000;
			// PEs: 40, 46 -> 47
			// srcs: (1570, 31)(3140) 47, (60) -2 --> (3197) -94:PEGB0, ND0, *, PENB
			10'd33 : rdata = 48'b000111110000000001100000000000000000000100000000;
			// PEs: 46, 47 -> 46
			// srcs: (1579, 60)(845) -1, (3981) -94 --> (4765) 93:NW0, PEGB7, -, NW0
			10'd34 : rdata = 48'b000100100000000011100001110000000100000000000000;
			// PEs: 40, 46 -> 
			// srcs: (1652, 32)(3140) 47, (142) 1 --> (3279) 47:PEGB0, ND1, *, 
			10'd35 : rdata = 48'b000111110000000001100000001000000000000000000000;
			// PEs: 46, 46 -> 
			// srcs: (1655, 45)(3) 1, (3279) 47 --> (4063) 47:NM0, ALU, *, 
			10'd36 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 46, 46 -> 46
			// srcs: (1658, 61)(927) 0, (4063) 47 --> (4847) -47:NW1, ALU, -, NW1
			10'd37 : rdata = 48'b000100100000000100111111111000000100010000000000;
			// PEs: 40, 46 -> 
			// srcs: (1700, 33)(3140) 47, (190) -2 --> (3327) -94:PEGB0, ND10, *, 
			10'd38 : rdata = 48'b000111110000000001100001010000000000000000000000;
			// PEs: 46, 46 -> 
			// srcs: (1703, 46)(3) 1, (3327) -94 --> (4111) -94:NM0, ALU, *, 
			10'd39 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 46, 46 -> 46
			// srcs: (1706, 62)(975) -1, (4111) -94 --> (4895) 93:NW10, ALU, -, NW10
			10'd40 : rdata = 48'b000100100000101000111111111000000110100000000000;
			// PEs: 40, 46 -> 
			// srcs: (1732, 34)(3140) 47, (222) -1 --> (3359) -47:PEGB0, ND2, *, 
			10'd41 : rdata = 48'b000111110000000001100000010000000000000000000000;
			// PEs: 46, 46 -> 
			// srcs: (1735, 47)(3) 1, (3359) -47 --> (4143) -47:NM0, ALU, *, 
			10'd42 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 46, 46 -> 46
			// srcs: (1738, 63)(1007) 0, (4143) -47 --> (4927) 47:NW2, ALU, -, NW2
			10'd43 : rdata = 48'b000100100000001000111111111000000100100000000000;
			// PEs: 40, 46 -> 
			// srcs: (1812, 35)(3140) 47, (302) -1 --> (3439) -47:PEGB0, ND3, *, 
			10'd44 : rdata = 48'b000111110000000001100000011000000000000000000000;
			// PEs: 46, 46 -> 
			// srcs: (1815, 48)(3) 1, (3439) -47 --> (4223) -47:NM0, ALU, *, 
			10'd45 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 46, 46 -> 46
			// srcs: (1818, 64)(1087) 0, (4223) -47 --> (5007) 47:NW3, ALU, -, NW3
			10'd46 : rdata = 48'b000100100000001100111111111000000100110000000000;
			// PEs: 40, 46 -> 
			// srcs: (1884, 36)(3140) 47, (374) 2 --> (3511) 94:PEGB0, ND11, *, 
			10'd47 : rdata = 48'b000111110000000001100001011000000000000000000000;
			// PEs: 46, 46 -> 
			// srcs: (1887, 49)(3) 1, (3511) 94 --> (4295) 94:NM0, ALU, *, 
			10'd48 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 46, 46 -> 46
			// srcs: (1890, 65)(1159) 2, (4295) 94 --> (5079) -92:NW11, ALU, -, NW11
			10'd49 : rdata = 48'b000100100000101100111111111000000110110000000000;
			// PEs: 40, 46 -> 
			// srcs: (1894, 37)(3140) 47, (384) -3 --> (3521) -141:PEGB0, ND4, *, 
			10'd50 : rdata = 48'b000111110000000001100000100000000000000000000000;
			// PEs: 46, 46 -> 
			// srcs: (1897, 50)(3) 1, (3521) -141 --> (4305) -141:NM0, ALU, *, 
			10'd51 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 46, 46 -> 46
			// srcs: (1900, 66)(1169) 1, (4305) -141 --> (5089) 142:NW4, ALU, -, NW4
			10'd52 : rdata = 48'b000100100000010000111111111000000101000000000000;
			// PEs: 40, 46 -> 47
			// srcs: (1974, 38)(3140) 47, (464) -3 --> (3601) -141:PEGB0, ND5, *, PENB
			10'd53 : rdata = 48'b000111110000000001100000101000000000000100000000;
			// PEs: 46, 45 -> 45
			// srcs: (1975, 51)(3) 1, (3599) -47 --> (4383) -47:NM0, PENB, *, PEGB5
			10'd54 : rdata = 48'b000111000000000011011111110000000000000011010000;
			// PEs: 46, 47 -> 46
			// srcs: (1983, 67)(1249) -3, (4385) -141 --> (5169) 138:NW5, PEGB7, -, NW5
			10'd55 : rdata = 48'b000100100000010111100001110000000101010000000000;
			// PEs: 40, 46 -> 46
			// srcs: (2055, 39)(3140) 47, (545) -2 --> (3682) -94:PEGB0, ND6, *, NI0
			10'd56 : rdata = 48'b000111110000000001100000110100000000000000000000;
			// PEs: 46, 45 -> 45
			// srcs: (2057, 52)(3) 1, (3681) 47 --> (4465) 47:NM0, PENB, *, PEGB5
			10'd57 : rdata = 48'b000111000000000011011111110000000000000011010000;
			// PEs: 46, 46 -> 
			// srcs: (2058, 53)(3) 1, (3682) -94 --> (4466) -94:NM0, NI0, *, 
			10'd58 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 46, 46 -> 46
			// srcs: (2061, 68)(1330) -1, (4466) -94 --> (5250) 93:NW6, ALU, -, NW6
			10'd59 : rdata = 48'b000100100000011000111111111000000101100000000000;
			// PEs: 40, 46 -> 
			// srcs: (2068, 40)(3140) 47, (558) 2 --> (3695) 94:PEGB0, ND12, *, 
			10'd60 : rdata = 48'b000111110000000001100001100000000000000000000000;
			// PEs: 46, 46 -> 
			// srcs: (2071, 54)(3) 1, (3695) 94 --> (4479) 94:NM0, ALU, *, 
			10'd61 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 46, 46 -> 46
			// srcs: (2074, 69)(1343) -1, (4479) 94 --> (5263) -95:NW12, ALU, -, NW12
			10'd62 : rdata = 48'b000100100000110000111111111000000111000000000000;
			// PEs: 40, 46 -> 
			// srcs: (2136, 41)(3140) 47, (626) 1 --> (3763) 47:PEGB0, ND7, *, 
			10'd63 : rdata = 48'b000111110000000001100000111000000000000000000000;
			// PEs: 46, 46 -> 
			// srcs: (2139, 55)(3) 1, (3763) 47 --> (4547) 47:NM0, ALU, *, 
			10'd64 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 46, 46 -> 46
			// srcs: (2142, 70)(1411) -2, (4547) 47 --> (5331) -49:NW7, ALU, -, NW7
			10'd65 : rdata = 48'b000100100000011100111111111000000101110000000000;
			// PEs: 40, 46 -> 
			// srcs: (2216, 42)(3140) 47, (706) 1 --> (3843) 47:PEGB0, ND8, *, 
			10'd66 : rdata = 48'b000111110000000001100001000000000000000000000000;
			// PEs: 46, 46 -> 
			// srcs: (2219, 56)(3) 1, (3843) 47 --> (4627) 47:NM0, ALU, *, 
			10'd67 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 46, 46 -> 46
			// srcs: (2222, 71)(1491) -1, (4627) 47 --> (5411) -48:NW8, ALU, -, NW8
			10'd68 : rdata = 48'b000100100000100000111111111000000110000000000000;
			// PEs: 40, 46 -> 
			// srcs: (2248, 43)(3140) 47, (738) 2 --> (3875) 94:PEGB0, ND13, *, 
			10'd69 : rdata = 48'b000111110000000001100001101000000000000000000000;
			// PEs: 46, 46 -> 
			// srcs: (2251, 57)(3) 1, (3875) 94 --> (4659) 94:NM0, ALU, *, 
			10'd70 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 46, 46 -> 46
			// srcs: (2254, 72)(1523) 1, (4659) 94 --> (5443) -93:NW13, ALU, -, NW13
			10'd71 : rdata = 48'b000100100000110100111111111000000111010000000000;
			// PEs: 46, 45 -> 45
			// srcs: (2299, 58)(3) 1, (3923) 0 --> (4707) 0:NM0, PENB, *, PEGB5
			10'd72 : rdata = 48'b000111000000000011011111110000000000000011010000;
			default : rdata = 48'b000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 47) begin
	always @(*) begin
		case(address)
			// PEs: 47, 47 -> 40
			// srcs: (1, 0)(61) -2, (846) 1 --> (1630) -2:ND0, NW0, *, PENB
			10'd0 : rdata = 48'b000110110000000001000000000000000000000100000000;
			// PEs: 47, 47 -> 40
			// srcs: (2, 1)(143) -3, (928) 2 --> (1712) -6:ND1, NW1, *, PENB
			10'd1 : rdata = 48'b000110110000000101000000001000000000000100000000;
			// PEs: 47, 47 -> 40
			// srcs: (3, 2)(223) 0, (1008) 2 --> (1792) 0:ND2, NW2, *, PENB
			10'd2 : rdata = 48'b000110110000001001000000010000000000000100000000;
			// PEs: 47, 47 -> 40
			// srcs: (4, 3)(303) -1, (1088) -3 --> (1872) 3:ND3, NW3, *, PENB
			10'd3 : rdata = 48'b000110110000001101000000011000000000000100000000;
			// PEs: 47, 47 -> 40
			// srcs: (5, 4)(385) -3, (1170) -1 --> (1954) 3:ND4, NW4, *, PENB
			10'd4 : rdata = 48'b000110110000010001000000100000000000000100000000;
			// PEs: 47, 47 -> 40
			// srcs: (6, 5)(465) 1, (1250) 1 --> (2034) 1:ND5, NW5, *, PENB
			10'd5 : rdata = 48'b000110110000010101000000101000000000000100000000;
			// PEs: 47, 47 -> 47
			// srcs: (7, 6)(546) -1, (1331) -3 --> (2115) 3:ND6, NW6, *, NI0
			10'd6 : rdata = 48'b000110110000011001000000110100000000000000000000;
			// PEs: 47, 47 -> 40
			// srcs: (8, 7)(627) 2, (1412) 1 --> (2196) 2:ND7, NW7, *, PENB
			10'd7 : rdata = 48'b000110110000011101000000111000000000000100000000;
			// PEs: 47, 47 -> 44
			// srcs: (9, 8)(707) 1, (1492) -1 --> (2276) -1:ND8, NW8, *, PEGB4
			10'd8 : rdata = 48'b000110110000100001000001000000000000000011000000;
			// PEs: 47, 47 -> 40
			// srcs: (10, 9)(13) -3, (798) 2 --> (1582) -6:ND9, NW9, *, PENB
			10'd9 : rdata = 48'b000110110000100101000001001000000000000100000000;
			// PEs: 47, 47 -> 40
			// srcs: (11, 10)(193) 0, (978) 0 --> (1762) 0:ND10, NW10, *, PENB
			10'd10 : rdata = 48'b000110110000101001000001010000000000000100000000;
			// PEs: 47, 47 -> 47
			// srcs: (12, 11)(377) -2, (1162) 2 --> (1946) -4:ND11, NW11, *, NI1
			10'd11 : rdata = 48'b000110110000101101000001011100001000000000000000;
			// PEs: 47, 47 -> 40
			// srcs: (13, 12)(561) 2, (1346) -2 --> (2130) -4:ND12, NW12, *, PENB
			10'd12 : rdata = 48'b000110110000110001000001100000000000000100000000;
			// PEs: 47, 47 -> 40
			// srcs: (14, 13)(745) -2, (1530) -2 --> (2314) 4:ND13, NW13, *, PENB
			10'd13 : rdata = 48'b000110110000110101000001101000000000000100000000;
			// PEs: 40 -> 
			// srcs: (36, 14)(1780) -6 --> (1780) -6:PEGB0, pass, 
			10'd14 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 40, 47 -> 47
			// srcs: (45, 15)(1779) 0, (1780) -6 --> (2560) -6:PEGB0, ALU, +, NI2
			10'd15 : rdata = 48'b000011110000000000111111111100010000000000000000;
			// PEs: 45, 47 -> 47
			// srcs: (94, 22)(2723) 2, (1946) -4 --> (2724) -2:PEGB5, NI1, +, NI3
			10'd16 : rdata = 48'b000011110000101010100000001100011000000000000000;
			// PEs: 40 -> 
			// srcs: (126, 16)(2106) -6 --> (2106) -6:PEGB0, pass, 
			10'd17 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 47, 41 -> 42
			// srcs: (128, 17)(2106) -6, (2107) 3 --> (2885) -3:ALU, PEGB1, +, PEGB2
			10'd18 : rdata = 48'b000010011111111111100000010000000000000010100000;
			// PEs: 41 -> 
			// srcs: (129, 20)(2714) 1 --> (2714) 1:PEGB1, pass, 
			10'd19 : rdata = 48'b110001110000001000000000000000000000000000000000;
			// PEs: 47, 44 -> 
			// srcs: (131, 21)(2714) 1, (1937) 6 --> (2715) 7:ALU, PEGB4, +, 
			10'd20 : rdata = 48'b000010011111111111100001000000000000000000000000;
			// PEs: 47, 46 -> 46
			// srcs: (134, 25)(2715) 7, (2717) -4 --> (2718) 3:ALU, PENB, +, PEGB6
			10'd21 : rdata = 48'b000010011111111111011111110000000000000011100000;
			// PEs: 46, 47 -> 47
			// srcs: (135, 26)(2722) 6, (2724) -2 --> (2725) 4:PENB, NI3, +, NI1
			10'd22 : rdata = 48'b000011101111111010100000011100001000000000000000;
			// PEs: 47 -> 40
			// srcs: (157, 18)(2115) 3 --> (2115) 3:NI0, pass, PENB
			10'd23 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 47 -> 40
			// srcs: (194, 19)(2560) -6 --> (2560) -6:NI2, pass, PENB
			10'd24 : rdata = 48'b110001010000001000000000000000000000000100000000;
			// PEs: 40 -> 
			// srcs: (613, 23)(2102) 0 --> (2102) 0:PEGB0, pass, 
			10'd25 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 41, 47 -> 43
			// srcs: (615, 24)(2880) 3, (2102) 0 --> (2881) 3:PEGB1, ALU, +, PEGB3
			10'd26 : rdata = 48'b000011110000001000111111111000000000000010110000;
			// PEs: 47 -> 40
			// srcs: (755, 27)(2725) 4 --> (2725) 4:NI1, pass, PENB
			10'd27 : rdata = 48'b110001010000000100000000000000000000000100000000;
			// PEs: 40, 47 -> 
			// srcs: (1524, 28)(3140) 47, (13) -3 --> (3150) -141:PEGB0, ND9, *, 
			10'd28 : rdata = 48'b000111110000000001100001001000000000000000000000;
			// PEs: 47, 47 -> 
			// srcs: (1527, 42)(3) 1, (3150) -141 --> (3934) -141:NM0, ALU, *, 
			10'd29 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 47, 47 -> 47
			// srcs: (1530, 58)(798) 2, (3934) -141 --> (4718) 143:NW9, ALU, -, NW9
			10'd30 : rdata = 48'b000100100000100100111111111000000110010000000000;
			// PEs: 40, 47 -> 47
			// srcs: (1571, 29)(3140) 47, (61) -2 --> (3198) -94:PEGB0, ND0, *, NI0
			10'd31 : rdata = 48'b000111110000000001100000000100000000000000000000;
			// PEs: 47, 46 -> 46
			// srcs: (1573, 43)(3) 1, (3197) -94 --> (3981) -94:NM0, PENB, *, PEGB6
			10'd32 : rdata = 48'b000111000000000011011111110000000000000011100000;
			// PEs: 47, 47 -> 
			// srcs: (1574, 44)(3) 1, (3198) -94 --> (3982) -94:NM0, NI0, *, 
			10'd33 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 47, 47 -> 47
			// srcs: (1577, 59)(846) 1, (3982) -94 --> (4766) 95:NW0, ALU, -, NW0
			10'd34 : rdata = 48'b000100100000000000111111111000000100000000000000;
			// PEs: 40, 47 -> 
			// srcs: (1653, 30)(3140) 47, (143) -3 --> (3280) -141:PEGB0, ND1, *, 
			10'd35 : rdata = 48'b000111110000000001100000001000000000000000000000;
			// PEs: 47, 47 -> 
			// srcs: (1656, 45)(3) 1, (3280) -141 --> (4064) -141:NM0, ALU, *, 
			10'd36 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 47, 47 -> 47
			// srcs: (1659, 60)(928) 2, (4064) -141 --> (4848) 143:NW1, ALU, -, NW1
			10'd37 : rdata = 48'b000100100000000100111111111000000100010000000000;
			// PEs: 40, 47 -> 
			// srcs: (1703, 31)(3140) 47, (193) 0 --> (3330) 0:PEGB0, ND10, *, 
			10'd38 : rdata = 48'b000111110000000001100001010000000000000000000000;
			// PEs: 47, 47 -> 
			// srcs: (1706, 46)(3) 1, (3330) 0 --> (4114) 0:NM0, ALU, *, 
			10'd39 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 47, 47 -> 47
			// srcs: (1709, 61)(978) 0, (4114) 0 --> (4898) 0:NW10, ALU, -, NW10
			10'd40 : rdata = 48'b000100100000101000111111111000000110100000000000;
			// PEs: 40, 47 -> 
			// srcs: (1733, 32)(3140) 47, (223) 0 --> (3360) 0:PEGB0, ND2, *, 
			10'd41 : rdata = 48'b000111110000000001100000010000000000000000000000;
			// PEs: 47, 47 -> 
			// srcs: (1736, 47)(3) 1, (3360) 0 --> (4144) 0:NM0, ALU, *, 
			10'd42 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 47, 47 -> 47
			// srcs: (1739, 62)(1008) 2, (4144) 0 --> (4928) 2:NW2, ALU, -, NW2
			10'd43 : rdata = 48'b000100100000001000111111111000000100100000000000;
			// PEs: 40, 47 -> 
			// srcs: (1813, 33)(3140) 47, (303) -1 --> (3440) -47:PEGB0, ND3, *, 
			10'd44 : rdata = 48'b000111110000000001100000011000000000000000000000;
			// PEs: 47, 47 -> 
			// srcs: (1816, 48)(3) 1, (3440) -47 --> (4224) -47:NM0, ALU, *, 
			10'd45 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 47, 47 -> 47
			// srcs: (1819, 63)(1088) -3, (4224) -47 --> (5008) 44:NW3, ALU, -, NW3
			10'd46 : rdata = 48'b000100100000001100111111111000000100110000000000;
			// PEs: 40, 47 -> 
			// srcs: (1887, 34)(3140) 47, (377) -2 --> (3514) -94:PEGB0, ND11, *, 
			10'd47 : rdata = 48'b000111110000000001100001011000000000000000000000;
			// PEs: 47, 47 -> 
			// srcs: (1890, 49)(3) 1, (3514) -94 --> (4298) -94:NM0, ALU, *, 
			10'd48 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 47, 47 -> 47
			// srcs: (1893, 64)(1162) 2, (4298) -94 --> (5082) 96:NW11, ALU, -, NW11
			10'd49 : rdata = 48'b000100100000101100111111111000000110110000000000;
			// PEs: 40, 47 -> 
			// srcs: (1895, 35)(3140) 47, (385) -3 --> (3522) -141:PEGB0, ND4, *, 
			10'd50 : rdata = 48'b000111110000000001100000100000000000000000000000;
			// PEs: 47, 47 -> 
			// srcs: (1898, 50)(3) 1, (3522) -141 --> (4306) -141:NM0, ALU, *, 
			10'd51 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 47, 47 -> 47
			// srcs: (1901, 65)(1170) -1, (4306) -141 --> (5090) 140:NW4, ALU, -, NW4
			10'd52 : rdata = 48'b000100100000010000111111111000000101000000000000;
			// PEs: 40, 47 -> 47
			// srcs: (1975, 36)(3140) 47, (465) 1 --> (3602) 47:PEGB0, ND5, *, NI0
			10'd53 : rdata = 48'b000111110000000001100000101100000000000000000000;
			// PEs: 47, 46 -> 46
			// srcs: (1977, 51)(3) 1, (3601) -141 --> (4385) -141:NM0, PENB, *, PEGB6
			10'd54 : rdata = 48'b000111000000000011011111110000000000000011100000;
			// PEs: 47, 47 -> 
			// srcs: (1978, 52)(3) 1, (3602) 47 --> (4386) 47:NM0, NI0, *, 
			10'd55 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 47, 47 -> 47
			// srcs: (1981, 66)(1250) 1, (4386) 47 --> (5170) -46:NW5, ALU, -, NW5
			10'd56 : rdata = 48'b000100100000010100111111111000000101010000000000;
			// PEs: 40, 47 -> 
			// srcs: (2056, 37)(3140) 47, (546) -1 --> (3683) -47:PEGB0, ND6, *, 
			10'd57 : rdata = 48'b000111110000000001100000110000000000000000000000;
			// PEs: 47, 47 -> 
			// srcs: (2059, 53)(3) 1, (3683) -47 --> (4467) -47:NM0, ALU, *, 
			10'd58 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 47, 47 -> 47
			// srcs: (2062, 67)(1331) -3, (4467) -47 --> (5251) 44:NW6, ALU, -, NW6
			10'd59 : rdata = 48'b000100100000011000111111111000000101100000000000;
			// PEs: 40, 47 -> 
			// srcs: (2071, 38)(3140) 47, (561) 2 --> (3698) 94:PEGB0, ND12, *, 
			10'd60 : rdata = 48'b000111110000000001100001100000000000000000000000;
			// PEs: 47, 47 -> 
			// srcs: (2074, 54)(3) 1, (3698) 94 --> (4482) 94:NM0, ALU, *, 
			10'd61 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 47, 47 -> 47
			// srcs: (2077, 68)(1346) -2, (4482) 94 --> (5266) -96:NW12, ALU, -, NW12
			10'd62 : rdata = 48'b000100100000110000111111111000000111000000000000;
			// PEs: 40, 47 -> 
			// srcs: (2137, 39)(3140) 47, (627) 2 --> (3764) 94:PEGB0, ND7, *, 
			10'd63 : rdata = 48'b000111110000000001100000111000000000000000000000;
			// PEs: 47, 47 -> 
			// srcs: (2140, 55)(3) 1, (3764) 94 --> (4548) 94:NM0, ALU, *, 
			10'd64 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 47, 47 -> 47
			// srcs: (2143, 69)(1412) 1, (4548) 94 --> (5332) -93:NW7, ALU, -, NW7
			10'd65 : rdata = 48'b000100100000011100111111111000000101110000000000;
			// PEs: 40, 47 -> 
			// srcs: (2217, 40)(3140) 47, (707) 1 --> (3844) 47:PEGB0, ND8, *, 
			10'd66 : rdata = 48'b000111110000000001100001000000000000000000000000;
			// PEs: 47, 47 -> 
			// srcs: (2220, 56)(3) 1, (3844) 47 --> (4628) 47:NM0, ALU, *, 
			10'd67 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 47, 47 -> 47
			// srcs: (2223, 70)(1492) -1, (4628) 47 --> (5412) -48:NW8, ALU, -, NW8
			10'd68 : rdata = 48'b000100100000100000111111111000000110000000000000;
			// PEs: 40, 47 -> 
			// srcs: (2255, 41)(3140) 47, (745) -2 --> (3882) -94:PEGB0, ND13, *, 
			10'd69 : rdata = 48'b000111110000000001100001101000000000000000000000;
			// PEs: 47, 47 -> 
			// srcs: (2258, 57)(3) 1, (3882) -94 --> (4666) -94:NM0, ALU, *, 
			10'd70 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 47, 47 -> 47
			// srcs: (2261, 71)(1530) -2, (4666) -94 --> (5450) 92:NW13, ALU, -, NW13
			10'd71 : rdata = 48'b000100100000110100111111111000000111010000000000;
			default : rdata = 48'b000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 48) begin
	always @(*) begin
		case(address)
			// PEs: 49 -> 16
			// srcs: (6, 0)(1632) 0 --> (1632) 0:PEGB1, pass, PUGB2
			10'd0 : rdata = 48'b110001110000001000000000000000000000000000001010;
			// PEs: 50 -> 16
			// srcs: (7, 1)(1633) -6 --> (1633) -6:PEGB2, pass, PUGB2
			10'd1 : rdata = 48'b110001110000010000000000000000000000000000001010;
			// PEs: 51 -> 24
			// srcs: (8, 2)(1635) -1 --> (1635) -1:PEGB3, pass, PUGB3
			10'd2 : rdata = 48'b110001110000011000000000000000000000000000001011;
			// PEs: 52 -> 24
			// srcs: (9, 3)(1636) 0 --> (1636) 0:PEGB4, pass, PUGB3
			10'd3 : rdata = 48'b110001110000100000000000000000000000000000001011;
			// PEs: 53 -> 24
			// srcs: (10, 4)(1638) 0 --> (1638) 0:PEGB5, pass, PUGB3
			10'd4 : rdata = 48'b110001110000101000000000000000000000000000001011;
			// PEs: 54 -> 24
			// srcs: (11, 5)(1639) 3 --> (1639) 3:PEGB6, pass, PUGB3
			10'd5 : rdata = 48'b110001110000110000000000000000000000000000001011;
			// PEs: 55 -> 24
			// srcs: (12, 6)(1641) -6 --> (1641) -6:PENB, pass, PUGB3
			10'd6 : rdata = 48'b110001101111111000000000000000000000000000001011;
			// PEs: 32 -> 48
			// srcs: (13, 10)(1702) -4 --> (1702) -4:PUGB4, pass, NI0
			10'd7 : rdata = 48'b110001110000100100000000000100000000000000000000;
			// PEs: 40 -> 50
			// srcs: (14, 11)(1703) 3 --> (1703) 3:PUNB, pass, PEGB2
			10'd8 : rdata = 48'b110001101111111100000000000000000000000010100000;
			// PEs: 40 -> 48
			// srcs: (15, 13)(1705) 6 --> (1705) 6:PUNB, pass, NI1
			10'd9 : rdata = 48'b110001101111111100000000000100001000000000000000;
			// PEs: 40 -> 51
			// srcs: (16, 14)(1706) 2 --> (1706) 2:PUNB, pass, PEGB3
			10'd10 : rdata = 48'b110001101111111100000000000000000000000010110000;
			// PEs: 40 -> 48
			// srcs: (17, 16)(1708) 0 --> (1708) 0:PUNB, pass, NI2
			10'd11 : rdata = 48'b110001101111111100000000000100010000000000000000;
			// PEs: 49 -> 56
			// srcs: (18, 22)(1714) 9 --> (1714) 9:PEGB1, pass, PUNB
			10'd12 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 50 -> 56
			// srcs: (19, 23)(1715) -2 --> (1715) -2:PEGB2, pass, PUNB
			10'd13 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 51 -> 56
			// srcs: (20, 24)(1717) 0 --> (1717) 0:PEGB3, pass, PUNB
			10'd14 : rdata = 48'b110001110000011000000000000000000000001000000000;
			// PEs: 52 -> 56
			// srcs: (21, 25)(1718) 2 --> (1718) 2:PEGB4, pass, PUNB
			10'd15 : rdata = 48'b110001110000100000000000000000000000001000000000;
			// PEs: 40 -> 52
			// srcs: (22, 17)(1709) 0 --> (1709) 0:PUNB, pass, PEGB4
			10'd16 : rdata = 48'b110001101111111100000000000000000000000011000000;
			// PEs: 48 -> 50
			// srcs: (23, 12)(1702) -4 --> (1702) -4:NI0, pass, PEGB2
			10'd17 : rdata = 48'b110001010000000000000000000000000000000010100000;
			// PEs: 40 -> 48
			// srcs: (24, 19)(1711) 0 --> (1711) 0:PUNB, pass, NI0
			10'd18 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 48 -> 51
			// srcs: (25, 15)(1705) 6 --> (1705) 6:NI1, pass, PEGB3
			10'd19 : rdata = 48'b110001010000000100000000000000000000000010110000;
			// PEs: 40 -> 53
			// srcs: (26, 20)(1712) -6 --> (1712) -6:PUNB, pass, PEGB5
			10'd20 : rdata = 48'b110001101111111100000000000000000000000011010000;
			// PEs: 32 -> 48
			// srcs: (27, 26)(1782) 3 --> (1782) 3:PUGB4, pass, NI1
			10'd21 : rdata = 48'b110001110000100100000000000100001000000000000000;
			// PEs: 49 -> 56
			// srcs: (28, 32)(1794) 0 --> (1794) 0:PEGB1, pass, PUNB
			10'd22 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 50 -> 56
			// srcs: (29, 33)(1795) -4 --> (1795) -4:PEGB2, pass, PUNB
			10'd23 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 51 -> 56
			// srcs: (30, 34)(1797) -4 --> (1797) -4:PEGB3, pass, PUNB
			10'd24 : rdata = 48'b110001110000011000000000000000000000001000000000;
			// PEs: 48 -> 52
			// srcs: (31, 18)(1708) 0 --> (1708) 0:NI2, pass, PEGB4
			10'd25 : rdata = 48'b110001010000001000000000000000000000000011000000;
			// PEs: 52 -> 56
			// srcs: (32, 35)(1798) -3 --> (1798) -3:PEGB4, pass, PUNB
			10'd26 : rdata = 48'b110001110000100000000000000000000000001000000000;
			// PEs: 53 -> 56
			// srcs: (33, 36)(1800) -2 --> (1800) -2:PEGB5, pass, PUNB
			10'd27 : rdata = 48'b110001110000101000000000000000000000001000000000;
			// PEs: 40 -> 54
			// srcs: (34, 27)(1783) 2 --> (1783) 2:PUNB, pass, PEGB6
			10'd28 : rdata = 48'b110001101111111100000000000000000000000011100000;
			// PEs: 48 -> 53
			// srcs: (35, 21)(1711) 0 --> (1711) 0:NI0, pass, PEGB5
			10'd29 : rdata = 48'b110001010000000000000000000000000000000011010000;
			// PEs: 40 -> 48
			// srcs: (36, 29)(1785) 2 --> (1785) 2:PUNB, pass, NI0
			10'd30 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 54 -> 56
			// srcs: (37, 37)(1801) 0 --> (1801) 0:PEGB6, pass, PUNB
			10'd31 : rdata = 48'b110001110000110000000000000000000000001000000000;
			// PEs: 40 -> 55
			// srcs: (38, 30)(1786) 2 --> (1786) 2:PUNB, pass, PEGB7
			10'd32 : rdata = 48'b110001101111111100000000000000000000000011110000;
			// PEs: 8 -> 48
			// srcs: (39, 7)(1668) 9 --> (1668) 9:PUGB1, pass, NI2
			10'd33 : rdata = 48'b110001110000001100000000000100010000000000000000;
			// PEs: 8 -> 49
			// srcs: (40, 8)(1669) 0 --> (1669) 0:PUGB1, pass, PENB
			10'd34 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 55 -> 0
			// srcs: (41, 38)(1803) 0 --> (1803) 0:PENB, pass, PUGB0
			10'd35 : rdata = 48'b110001101111111000000000000000000000000000001000;
			// PEs: 32 -> 48
			// srcs: (42, 39)(1864) 1 --> (1864) 1:PUGB4, pass, NI3
			10'd36 : rdata = 48'b110001110000100100000000000100011000000000000000;
			// PEs: 48 -> 54
			// srcs: (43, 28)(1782) 3 --> (1782) 3:NI1, pass, PEGB6
			10'd37 : rdata = 48'b110001010000000100000000000000000000000011100000;
			// PEs: 49 -> 56
			// srcs: (44, 45)(1874) -2 --> (1874) -2:PEGB1, pass, PUNB
			10'd38 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 50 -> 56
			// srcs: (45, 46)(1875) 0 --> (1875) 0:PEGB2, pass, PUNB
			10'd39 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 48 -> 49
			// srcs: (46, 9)(1668) 9 --> (1668) 9:NI2, pass, PENB
			10'd40 : rdata = 48'b110001010000001000000000000000000000000100000000;
			// PEs: 48 -> 55
			// srcs: (47, 31)(1785) 2 --> (1785) 2:NI0, pass, PEGB7
			10'd41 : rdata = 48'b110001010000000000000000000000000000000011110000;
			// PEs: 51 -> 40
			// srcs: (48, 47)(1877) 0 --> (1877) 0:PEGB3, pass, PUGB5
			10'd42 : rdata = 48'b110001110000011000000000000000000000000000001101;
			// PEs: 52 -> 40
			// srcs: (49, 48)(1878) -2 --> (1878) -2:PEGB4, pass, PUGB5
			10'd43 : rdata = 48'b110001110000100000000000000000000000000000001101;
			// PEs: 53 -> 56
			// srcs: (50, 49)(1880) -1 --> (1880) -1:PEGB5, pass, PUNB
			10'd44 : rdata = 48'b110001110000101000000000000000000000001000000000;
			// PEs: 54 -> 56
			// srcs: (51, 50)(1881) 1 --> (1881) 1:PEGB6, pass, PUNB
			10'd45 : rdata = 48'b110001110000110000000000000000000000001000000000;
			// PEs: 56 -> 49
			// srcs: (52, 51)(1884) -1 --> (1884) -1:PUGB7, pass, PENB
			10'd46 : rdata = 48'b110001110000111100000000000000000000000100000000;
			// PEs: 40 -> 50
			// srcs: (53, 40)(1865) -3 --> (1865) -3:PUNB, pass, PEGB2
			10'd47 : rdata = 48'b110001101111111100000000000000000000000010100000;
			// PEs: 40 -> 48
			// srcs: (54, 42)(1871) 0 --> (1871) 0:PUNB, pass, NI0
			10'd48 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 40 -> 51
			// srcs: (55, 43)(1872) 3 --> (1872) 3:PUNB, pass, PEGB3
			10'd49 : rdata = 48'b110001101111111100000000000000000000000010110000;
			// PEs: 56 -> 48
			// srcs: (56, 52)(1886) -6 --> (1886) -6:PUGB7, pass, NI1
			10'd50 : rdata = 48'b110001110000111100000000000100001000000000000000;
			// PEs: 56 -> 49
			// srcs: (57, 53)(1887) -2 --> (1887) -2:PUGB7, pass, PENB
			10'd51 : rdata = 48'b110001110000111100000000000000000000000100000000;
			// PEs: 49 -> 56
			// srcs: (58, 64)(1956) -2 --> (1956) -2:PEGB1, pass, PUNB
			10'd52 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 50 -> 56
			// srcs: (59, 65)(1957) 0 --> (1957) 0:PEGB2, pass, PUNB
			10'd53 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 51 -> 56
			// srcs: (60, 66)(1959) 0 --> (1959) 0:PEGB3, pass, PUNB
			10'd54 : rdata = 48'b110001110000011000000000000000000000001000000000;
			// PEs: 52 -> 56
			// srcs: (61, 67)(1960) 0 --> (1960) 0:PEGB4, pass, PUNB
			10'd55 : rdata = 48'b110001110000100000000000000000000000001000000000;
			// PEs: 48 -> 50
			// srcs: (62, 41)(1864) 1 --> (1864) 1:NI3, pass, PEGB2
			10'd56 : rdata = 48'b110001010000001100000000000000000000000010100000;
			// PEs: 48 -> 49
			// srcs: (63, 54)(1886) -6 --> (1886) -6:NI1, pass, PENB
			10'd57 : rdata = 48'b110001010000000100000000000000000000000100000000;
			// PEs: 48 -> 51
			// srcs: (64, 44)(1871) 0 --> (1871) 0:NI0, pass, PEGB3
			10'd58 : rdata = 48'b110001010000000000000000000000000000000010110000;
			// PEs: 40 -> 48
			// srcs: (65, 55)(1947) 1 --> (1947) 1:PUNB, pass, NI0
			10'd59 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 40 -> 49
			// srcs: (66, 56)(1948) -2 --> (1948) -2:PUNB, pass, PENB
			10'd60 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 53 -> 56
			// srcs: (67, 68)(1962) 6 --> (1962) 6:PEGB5, pass, PUNB
			10'd61 : rdata = 48'b110001110000101000000000000000000000001000000000;
			// PEs: 54 -> 56
			// srcs: (68, 69)(1963) 0 --> (1963) 0:PEGB6, pass, PUNB
			10'd62 : rdata = 48'b110001110000110000000000000000000000001000000000;
			// PEs: 49 -> 56
			// srcs: (69, 79)(2036) 0 --> (2036) 0:PEGB1, pass, PUNB
			10'd63 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 50 -> 56
			// srcs: (70, 80)(2037) -1 --> (2037) -1:PEGB2, pass, PUNB
			10'd64 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 51 -> 56
			// srcs: (71, 81)(2039) 3 --> (2039) 3:PEGB3, pass, PUNB
			10'd65 : rdata = 48'b110001110000011000000000000000000000001000000000;
			// PEs: 48 -> 49
			// srcs: (72, 57)(1947) 1 --> (1947) 1:NI0, pass, PENB
			10'd66 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 40 -> 48
			// srcs: (73, 58)(1950) 9 --> (1950) 9:PUNB, pass, NI0
			10'd67 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 40 -> 49
			// srcs: (74, 59)(1951) 6 --> (1951) 6:PUNB, pass, PENB
			10'd68 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 52 -> 56
			// srcs: (75, 82)(2040) 0 --> (2040) 0:PEGB4, pass, PUNB
			10'd69 : rdata = 48'b110001110000100000000000000000000000001000000000;
			// PEs: 53 -> 56
			// srcs: (76, 83)(2042) 2 --> (2042) 2:PEGB5, pass, PUNB
			10'd70 : rdata = 48'b110001110000101000000000000000000000001000000000;
			// PEs: 54 -> 56
			// srcs: (77, 84)(2043) 3 --> (2043) 3:PEGB6, pass, PUNB
			10'd71 : rdata = 48'b110001110000110000000000000000000000001000000000;
			// PEs: 55 -> 56
			// srcs: (78, 85)(2045) -2 --> (2045) -2:PENB, pass, PUNB
			10'd72 : rdata = 48'b110001101111111000000000000000000000001000000000;
			// PEs: 49 -> 56
			// srcs: (79, 89)(2116) -2 --> (2116) -2:PEGB1, pass, PUNB
			10'd73 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 48 -> 49
			// srcs: (80, 60)(1950) 9 --> (1950) 9:NI0, pass, PENB
			10'd74 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 40 -> 48
			// srcs: (81, 61)(1953) -3 --> (1953) -3:PUNB, pass, NI0
			10'd75 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 40 -> 49
			// srcs: (82, 62)(1954) 3 --> (1954) 3:PUNB, pass, PENB
			10'd76 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 50 -> 56
			// srcs: (83, 90)(2117) 2 --> (2117) 2:PEGB2, pass, PUNB
			10'd77 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 51 -> 56
			// srcs: (84, 91)(2119) 4 --> (2119) 4:PEGB3, pass, PUNB
			10'd78 : rdata = 48'b110001110000011000000000000000000000001000000000;
			// PEs: 52 -> 56
			// srcs: (85, 92)(2120) 9 --> (2120) 9:PEGB4, pass, PUNB
			10'd79 : rdata = 48'b110001110000100000000000000000000000001000000000;
			// PEs: 53 -> 56
			// srcs: (86, 93)(2122) 0 --> (2122) 0:PEGB5, pass, PUNB
			10'd80 : rdata = 48'b110001110000101000000000000000000000001000000000;
			// PEs: 54 -> 56
			// srcs: (87, 94)(2123) 6 --> (2123) 6:PEGB6, pass, PUNB
			10'd81 : rdata = 48'b110001110000110000000000000000000000001000000000;
			// PEs: 48 -> 49
			// srcs: (88, 63)(1953) -3 --> (1953) -3:NI0, pass, PENB
			10'd82 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 40 -> 48
			// srcs: (89, 70)(2027) -6 --> (2027) -6:PUNB, pass, NI0
			10'd83 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 40 -> 49
			// srcs: (90, 71)(2028) 0 --> (2028) 0:PUNB, pass, PENB
			10'd84 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 55 -> 56
			// srcs: (91, 95)(2125) -2 --> (2125) -2:PENB, pass, PUNB
			10'd85 : rdata = 48'b110001101111111000000000000000000000001000000000;
			// PEs: 49 -> 56
			// srcs: (92, 105)(2198) 0 --> (2198) 0:PEGB1, pass, PUNB
			10'd86 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 50 -> 56
			// srcs: (93, 106)(2199) -4 --> (2199) -4:PEGB2, pass, PUNB
			10'd87 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 51 -> 56
			// srcs: (94, 107)(2201) 2 --> (2201) 2:PEGB3, pass, PUNB
			10'd88 : rdata = 48'b110001110000011000000000000000000000001000000000;
			// PEs: 52 -> 56
			// srcs: (95, 108)(2202) 2 --> (2202) 2:PEGB4, pass, PUNB
			10'd89 : rdata = 48'b110001110000100000000000000000000000001000000000;
			// PEs: 48 -> 49
			// srcs: (96, 72)(2027) -6 --> (2027) -6:NI0, pass, PENB
			10'd90 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 40 -> 48
			// srcs: (97, 73)(2030) -1 --> (2030) -1:PUNB, pass, NI0
			10'd91 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 40 -> 49
			// srcs: (98, 74)(2031) -2 --> (2031) -2:PUNB, pass, PENB
			10'd92 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 53 -> 56
			// srcs: (99, 109)(2204) -3 --> (2204) -3:PEGB5, pass, PUNB
			10'd93 : rdata = 48'b110001110000101000000000000000000000001000000000;
			// PEs: 54 -> 56
			// srcs: (100, 110)(2205) 2 --> (2205) 2:PEGB6, pass, PUNB
			10'd94 : rdata = 48'b110001110000110000000000000000000000001000000000;
			// PEs: 55 -> 56
			// srcs: (101, 111)(2207) -4 --> (2207) -4:PENB, pass, PUNB
			10'd95 : rdata = 48'b110001101111111000000000000000000000001000000000;
			// PEs: 55 -> 56
			// srcs: (102, 112)(2287) 0 --> (2287) 0:PENB, pass, PUNB
			10'd96 : rdata = 48'b110001101111111000000000000000000000001000000000;
			// PEs: 49 -> 16
			// srcs: (103, 133)(1585) -3 --> (1585) -3:PEGB1, pass, PUGB2
			10'd97 : rdata = 48'b110001110000001000000000000000000000000000001010;
			// PEs: 48 -> 49
			// srcs: (104, 75)(2030) -1 --> (2030) -1:NI0, pass, PENB
			10'd98 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 40 -> 48
			// srcs: (105, 76)(2033) 9 --> (2033) 9:PUNB, pass, NI0
			10'd99 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 40 -> 49
			// srcs: (106, 77)(2034) 1 --> (2034) 1:PUNB, pass, PENB
			10'd100 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 55 -> 0
			// srcs: (107, 118)(1722) -6 --> (1722) -6:PENB, pass, PUGB0
			10'd101 : rdata = 48'b110001101111111000000000000000000000000000001000;
			// PEs: 50 -> 32
			// srcs: (108, 134)(1588) 2 --> (1588) 2:PEGB2, pass, PUGB4
			10'd102 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 54 -> 8
			// srcs: (109, 138)(1600) -2 --> (1600) -2:PEGB6, pass, PUGB1
			10'd103 : rdata = 48'b110001110000110000000000000000000000000000001001;
			// PEs: 53 -> 56
			// srcs: (110, 116)(1720) 6 --> (1720) 6:PEGB5, pass, PUNB
			10'd104 : rdata = 48'b110001110000101000000000000000000000001000000000;
			// PEs: 50 -> 0
			// srcs: (111, 150)(2483) -1 --> (2483) -1:PEGB2, pass, PUGB0
			10'd105 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 48 -> 49
			// srcs: (112, 78)(2033) 9 --> (2033) 9:NI0, pass, PENB
			10'd106 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 40 -> 48
			// srcs: (113, 86)(2109) 6 --> (2109) 6:PUNB, pass, NI0
			10'd107 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 40 -> 49
			// srcs: (114, 87)(2110) 6 --> (2110) 6:PUNB, pass, PENB
			10'd108 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 55 -> 8
			// srcs: (115, 139)(1603) -3 --> (1603) -3:PENB, pass, PUGB1
			10'd109 : rdata = 48'b110001101111111000000000000000000000000000001001;
			// PEs: 51 -> 16
			// srcs: (116, 151)(2485) 8 --> (2485) 8:PEGB3, pass, PUGB2
			10'd110 : rdata = 48'b110001110000011000000000000000000000000000001010;
			// PEs: 49 -> 32
			// srcs: (117, 160)(1765) 0 --> (1765) 0:PEGB1, pass, PUGB4
			10'd111 : rdata = 48'b110001110000001000000000000000000000000000001100;
			// PEs: 54 -> 56
			// srcs: (118, 117)(1721) 1 --> (1721) 1:PEGB6, pass, PUNB
			10'd112 : rdata = 48'b110001110000110000000000000000000000001000000000;
			// PEs: 51 -> 8
			// srcs: (119, 169)(2652) 3 --> (2652) 3:PEGB3, pass, PUGB1
			10'd113 : rdata = 48'b110001110000011000000000000000000000000000001001;
			// PEs: 48 -> 49
			// srcs: (120, 88)(2109) 6 --> (2109) 6:NI0, pass, PENB
			10'd114 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 40 -> 48
			// srcs: (121, 96)(2189) -2 --> (2189) -2:PUNB, pass, NI0
			10'd115 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 40 -> 49
			// srcs: (122, 97)(2190) -2 --> (2190) -2:PUNB, pass, PENB
			10'd116 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 55 -> 56
			// srcs: (123, 125)(1965) -3 --> (1965) -3:PENB, pass, PUNB
			10'd117 : rdata = 48'b110001101111111000000000000000000000001000000000;
			// PEs: 52 -> 56
			// srcs: (124, 136)(1594) -1 --> (1594) -1:PEGB4, pass, PUNB
			10'd118 : rdata = 48'b110001110000100000000000000000000000001000000000;
			// PEs: 52 -> 40
			// srcs: (125, 152)(2489) 0 --> (2489) 0:PEGB4, pass, PUGB5
			10'd119 : rdata = 48'b110001110000100000000000000000000000000000001101;
			// PEs: 49 -> 0
			// srcs: (126, 173)(2663) -2 --> (2663) -2:PEGB1, pass, PUGB0
			10'd120 : rdata = 48'b110001110000001000000000000000000000000000001000;
			// PEs: 49 -> 40
			// srcs: (127, 174)(2666) -8 --> (2666) -8:PEGB1, pass, PUGB5
			10'd121 : rdata = 48'b110001110000001000000000000000000000000000001101;
			// PEs: 48 -> 49
			// srcs: (128, 98)(2189) -2 --> (2189) -2:NI0, pass, PENB
			10'd122 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 40 -> 48
			// srcs: (129, 99)(2192) -3 --> (2192) -3:PUNB, pass, NI0
			10'd123 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 40 -> 49
			// srcs: (130, 100)(2193) -6 --> (2193) -6:PUNB, pass, PENB
			10'd124 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 49 -> 0
			// srcs: (131, 194)(2808) -6 --> (2808) -6:PEGB1, pass, PUGB0
			10'd125 : rdata = 48'b110001110000001000000000000000000000000000001000;
			// PEs: 49 -> 16
			// srcs: (132, 195)(2810) -3 --> (2810) -3:PEGB1, pass, PUGB2
			10'd126 : rdata = 48'b110001110000001000000000000000000000000000001010;
			// PEs: 53 -> 56
			// srcs: (133, 153)(2491) -6 --> (2491) -6:PEGB5, pass, PUNB
			10'd127 : rdata = 48'b110001110000101000000000000000000000001000000000;
			// PEs: 50 -> 56
			// srcs: (134, 168)(2642) -2 --> (2642) -2:PEGB2, pass, PUNB
			10'd128 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 55 -> 8
			// srcs: (135, 184)(1971) -6 --> (1971) -6:PENB, pass, PUGB1
			10'd129 : rdata = 48'b110001101111111000000000000000000000000000001001;
			// PEs: 48 -> 49
			// srcs: (136, 101)(2192) -3 --> (2192) -3:NI0, pass, PENB
			10'd130 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 40 -> 48
			// srcs: (137, 102)(2195) -2 --> (2195) -2:PUNB, pass, NI0
			10'd131 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 40 -> 49
			// srcs: (138, 103)(2196) 2 --> (2196) 2:PUNB, pass, PENB
			10'd132 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 49 -> 32
			// srcs: (139, 196)(2813) 10 --> (2813) 10:PEGB1, pass, PUGB4
			10'd133 : rdata = 48'b110001110000001000000000000000000000000000001100;
			// PEs: 52 -> 56
			// srcs: (142, 181)(1958) 4 --> (1958) 4:PEGB4, pass, PUNB
			10'd134 : rdata = 48'b110001110000100000000000000000000000001000000000;
			// PEs: 49 -> 16
			// srcs: (143, 212)(2972) -9 --> (2972) -9:PEGB1, pass, PUGB2
			10'd135 : rdata = 48'b110001110000001000000000000000000000000000001010;
			// PEs: 48 -> 49
			// srcs: (144, 104)(2195) -2 --> (2195) -2:NI0, pass, PENB
			10'd136 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 55 -> 24
			// srcs: (145, 204)(2151) 0 --> (2151) 0:PENB, pass, PUGB3
			10'd137 : rdata = 48'b110001101111111000000000000000000000000000001011;
			// PEs: 52 -> 40
			// srcs: (147, 201)(2142) -2 --> (2142) -2:PEGB4, pass, PUGB5
			10'd138 : rdata = 48'b110001110000100000000000000000000000000000001101;
			// PEs: 53 -> 32
			// srcs: (148, 202)(2145) 1 --> (2145) 1:PEGB5, pass, PUGB4
			10'd139 : rdata = 48'b110001110000101000000000000000000000000000001100;
			// PEs: 50 -> 0
			// srcs: (149, 227)(2320) 0 --> (2320) 0:PEGB2, pass, PUGB0
			10'd140 : rdata = 48'b110001110000010000000000000000000000000000001000;
			// PEs: 53 -> 56
			// srcs: (150, 182)(1961) 3 --> (1961) 3:PEGB5, pass, PUNB
			10'd141 : rdata = 48'b110001110000101000000000000000000000001000000000;
			// PEs: 53 -> 24
			// srcs: (153, 218)(3059) -4 --> (3059) -4:PEGB5, pass, PUGB3
			10'd142 : rdata = 48'b110001110000101000000000000000000000000000001011;
			// PEs: 55 -> 32
			// srcs: (154, 219)(3064) -2 --> (3064) -2:PENB, pass, PUGB4
			10'd143 : rdata = 48'b110001101111111000000000000000000000000000001100;
			// PEs: 53 -> 16
			// srcs: (155, 230)(2329) -4 --> (2329) -4:PEGB5, pass, PUGB2
			10'd144 : rdata = 48'b110001110000101000000000000000000000000000001010;
			// PEs: 54 -> 56
			// srcs: (158, 183)(1964) 9 --> (1964) 9:PEGB6, pass, PUNB
			10'd145 : rdata = 48'b110001110000110000000000000000000000001000000000;
			// PEs: 55 -> 24
			// srcs: (160, 232)(2335) -2 --> (2335) -2:PENB, pass, PUGB3
			10'd146 : rdata = 48'b110001101111111000000000000000000000000000001011;
			// PEs: 51 -> 32
			// srcs: (162, 228)(2323) 2 --> (2323) 2:PEGB3, pass, PUGB4
			10'd147 : rdata = 48'b110001110000011000000000000000000000000000001100;
			// PEs: 52 -> 56
			// srcs: (166, 217)(3057) -5 --> (3057) -5:PEGB4, pass, PUNB
			10'd148 : rdata = 48'b110001110000100000000000000000000000001000000000;
			// PEs: 49 -> 56
			// srcs: (174, 226)(2317) 0 --> (2317) 0:PEGB1, pass, PUNB
			10'd149 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 52 -> 56
			// srcs: (182, 229)(2326) -2 --> (2326) -2:PEGB4, pass, PUNB
			10'd150 : rdata = 48'b110001110000100000000000000000000000001000000000;
			// PEs: 40 -> 48
			// srcs: (191, 119)(1867) 6 --> (1867) 6:PUNB, pass, NI0
			10'd151 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 40 -> 50
			// srcs: (216, 120)(1868) -1 --> (1868) -1:PUNB, pass, PEGB2
			10'd152 : rdata = 48'b110001101111111100000000000000000000000010100000;
			// PEs: 0 -> 48
			// srcs: (221, 113)(1573) 6 --> (1573) 6:PUGB0, pass, NI1
			10'd153 : rdata = 48'b110001110000000100000000000100001000000000000000;
			// PEs: 48 -> 50
			// srcs: (225, 121)(1867) 6 --> (1867) 6:NI0, pass, PEGB2
			10'd154 : rdata = 48'b110001010000000000000000000000000000000010100000;
			// PEs: 40 -> 48
			// srcs: (234, 122)(1869) 0 --> (1869) 0:PUNB, pass, NI0
			10'd155 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 0 -> 54
			// srcs: (237, 114)(1574) 3 --> (1574) 3:PUGB0, pass, PEGB6
			10'd156 : rdata = 48'b110001110000000100000000000000000000000011100000;
			// PEs: 48 -> 54
			// srcs: (246, 115)(1573) 6 --> (1573) 6:NI1, pass, PEGB6
			10'd157 : rdata = 48'b110001010000000100000000000000000000000011100000;
			// PEs: 40 -> 51
			// srcs: (251, 123)(1870) 0 --> (1870) 0:PUNB, pass, PEGB3
			10'd158 : rdata = 48'b110001101111111100000000000000000000000010110000;
			// PEs: 48 -> 51
			// srcs: (260, 124)(1869) 0 --> (1869) 0:NI0, pass, PEGB3
			10'd159 : rdata = 48'b110001010000000000000000000000000000000010110000;
			// PEs: 40 -> 48
			// srcs: (264, 126)(2112) 9 --> (2112) 9:PUNB, pass, NI0
			10'd160 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 40 -> 49
			// srcs: (280, 127)(2113) -1 --> (2113) -1:PUNB, pass, PENB
			10'd161 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 48 -> 49
			// srcs: (286, 128)(2112) 9 --> (2112) 9:NI0, pass, PENB
			10'd162 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 40 -> 48
			// srcs: (296, 129)(2114) 2 --> (2114) 2:PUNB, pass, NI0
			10'd163 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 40 -> 49
			// srcs: (309, 130)(2115) 3 --> (2115) 3:PUNB, pass, PENB
			10'd164 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 48 -> 49
			// srcs: (315, 131)(2114) 2 --> (2114) 2:NI0, pass, PENB
			10'd165 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 56 -> 49
			// srcs: (316, 132)(2358) 0 --> (2358) 0:PUGB7, pass, PENB
			10'd166 : rdata = 48'b110001110000111100000000000000000000000100000000;
			// PEs: 0 -> 49
			// srcs: (317, 135)(2371) 9 --> (2371) 9:PUGB0, pass, PENB
			10'd167 : rdata = 48'b110001110000000100000000000000000000000100000000;
			// PEs: 0 -> 49
			// srcs: (318, 137)(2376) -6 --> (2376) -6:PUGB0, pass, PENB
			10'd168 : rdata = 48'b110001110000000100000000000000000000000100000000;
			// PEs: 16 -> 48
			// srcs: (319, 140)(2399) 0 --> (2399) 0:PUGB2, pass, NI0
			10'd169 : rdata = 48'b110001110000010100000000000100000000000000000000;
			// PEs: 56 -> 49
			// srcs: (320, 141)(1621) 2 --> (1621) 2:PUGB7, pass, PENB
			10'd170 : rdata = 48'b110001110000111100000000000000000000000100000000;
			// PEs: 49 -> 16
			// srcs: (323, 233)(2359) 9 --> (2359) 9:PEGB1, pass, PUGB2
			10'd171 : rdata = 48'b110001110000001000000000000000000000000000001010;
			// PEs: 49 -> 0
			// srcs: (324, 237)(2372) 11 --> (2372) 11:PEGB1, pass, PUGB0
			10'd172 : rdata = 48'b110001110000001000000000000000000000000000001000;
			// PEs: 49 -> 56
			// srcs: (325, 238)(2377) -6 --> (2377) -6:PEGB1, pass, PUNB
			10'd173 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 48 -> 49
			// srcs: (326, 142)(2399) 0 --> (2399) 0:NI0, pass, PENB
			10'd174 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 32 -> 48
			// srcs: (327, 143)(2440) 2 --> (2440) 2:PUGB4, pass, NI0
			10'd175 : rdata = 48'b110001110000100100000000000100000000000000000000;
			// PEs: 8 -> 49
			// srcs: (328, 144)(1661) 0 --> (1661) 0:PUGB1, pass, PENB
			10'd176 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 49 -> 40
			// srcs: (333, 239)(2400) 2 --> (2400) 2:PEGB1, pass, PUGB5
			10'd177 : rdata = 48'b110001110000001000000000000000000000000000001101;
			// PEs: 48 -> 49
			// srcs: (334, 145)(2440) 2 --> (2440) 2:NI0, pass, PENB
			10'd178 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 8 -> 49
			// srcs: (335, 146)(1670) -6 --> (1670) -6:PUGB1, pass, PENB
			10'd179 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 40 -> 48
			// srcs: (336, 147)(2473) -6 --> (2473) -6:PUNB, pass, NI0
			10'd180 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 16 -> 49
			// srcs: (337, 148)(1695) 3 --> (1695) 3:PUGB2, pass, PENB
			10'd181 : rdata = 48'b110001110000010100000000000000000000000100000000;
			// PEs: 49 -> 40
			// srcs: (341, 243)(2441) 2 --> (2441) 2:PEGB1, pass, PUGB5
			10'd182 : rdata = 48'b110001110000001000000000000000000000000000001101;
			// PEs: 49 -> 56
			// srcs: (342, 244)(2448) 3 --> (2448) 3:PEGB1, pass, PUNB
			10'd183 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 48 -> 49
			// srcs: (343, 149)(2473) -6 --> (2473) -6:NI0, pass, PENB
			10'd184 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 0 -> 48
			// srcs: (344, 154)(2508) 6 --> (2508) 6:PUGB0, pass, NI0
			10'd185 : rdata = 48'b110001110000000100000000000100000000000000000000;
			// PEs: 32 -> 49
			// srcs: (345, 155)(1729) -3 --> (1729) -3:PUGB4, pass, PENB
			10'd186 : rdata = 48'b110001110000100100000000000000000000000100000000;
			// PEs: 49 -> 0
			// srcs: (350, 248)(2474) -3 --> (2474) -3:PEGB1, pass, PUGB0
			10'd187 : rdata = 48'b110001110000001000000000000000000000000000001000;
			// PEs: 48 -> 49
			// srcs: (351, 156)(2508) 6 --> (2508) 6:NI0, pass, PENB
			10'd188 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 8 -> 48
			// srcs: (352, 157)(2533) -4 --> (2533) -4:PUGB1, pass, NI0
			10'd189 : rdata = 48'b110001110000001100000000000100000000000000000000;
			// PEs: 40 -> 49
			// srcs: (353, 158)(1756) -2 --> (1756) -2:PUNB, pass, PENB
			10'd190 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 49 -> 56
			// srcs: (358, 249)(2509) 3 --> (2509) 3:PEGB1, pass, PUNB
			10'd191 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 48 -> 49
			// srcs: (359, 159)(2533) -4 --> (2533) -4:NI0, pass, PENB
			10'd192 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 32 -> 49
			// srcs: (360, 161)(2544) -3 --> (2544) -3:PUGB4, pass, PENB
			10'd193 : rdata = 48'b110001110000100100000000000000000000000100000000;
			// PEs: 40 -> 49
			// srcs: (361, 162)(2555) 1 --> (2555) 1:PUNB, pass, PENB
			10'd194 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 40 -> 49
			// srcs: (362, 163)(2558) 11 --> (2558) 11:PUNB, pass, PENB
			10'd195 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 40 -> 49
			// srcs: (363, 164)(2560) -6 --> (2560) -6:PUNB, pass, PENB
			10'd196 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 40 -> 48
			// srcs: (364, 165)(2637) -2 --> (2637) -2:PUNB, pass, NI0
			10'd197 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 16 -> 49
			// srcs: (365, 166)(1860) 0 --> (1860) 0:PUGB2, pass, PENB
			10'd198 : rdata = 48'b110001110000010100000000000000000000000100000000;
			// PEs: 40 -> 48
			// srcs: (366, 170)(2657) -2 --> (2657) -2:PUNB, pass, NI1
			10'd199 : rdata = 48'b110001101111111100000000000100001000000000000000;
			// PEs: 16 -> 52
			// srcs: (367, 171)(1879) 4 --> (1879) 4:PUGB2, pass, PEGB4
			10'd200 : rdata = 48'b110001110000010100000000000000000000000011000000;
			// PEs: 49 -> 16
			// srcs: (368, 250)(2534) -6 --> (2534) -6:PEGB1, pass, PUGB2
			10'd201 : rdata = 48'b110001110000001000000000000000000000000000001010;
			// PEs: 49 -> 40
			// srcs: (369, 251)(2545) -5 --> (2545) -5:PEGB1, pass, PUGB5
			10'd202 : rdata = 48'b110001110000001000000000000000000000000000001101;
			// PEs: 51 -> 16
			// srcs: (370, 257)(2651) 5 --> (2651) 5:PEGB3, pass, PUGB2
			10'd203 : rdata = 48'b110001110000011000000000000000000000000000001010;
			// PEs: 48 -> 49
			// srcs: (371, 167)(2637) -2 --> (2637) -2:NI0, pass, PENB
			10'd204 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 0 -> 48
			// srcs: (372, 175)(2668) -2 --> (2668) -2:PUGB0, pass, NI0
			10'd205 : rdata = 48'b110001110000000100000000000100000000000000000000;
			// PEs: 24 -> 49
			// srcs: (373, 176)(1891) 2 --> (1891) 2:PUGB3, pass, PENB
			10'd206 : rdata = 48'b110001110000011100000000000000000000000100000000;
			// PEs: 48 -> 52
			// srcs: (376, 172)(2657) -2 --> (2657) -2:NI1, pass, PEGB4
			10'd207 : rdata = 48'b110001010000000100000000000000000000000011000000;
			// PEs: 48 -> 49
			// srcs: (379, 177)(2668) -2 --> (2668) -2:NI0, pass, PENB
			10'd208 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 16 -> 48
			// srcs: (380, 178)(2691) -2 --> (2691) -2:PUGB2, pass, NI0
			10'd209 : rdata = 48'b110001110000010100000000000100000000000000000000;
			// PEs: 32 -> 49
			// srcs: (381, 179)(1915) 0 --> (1915) 0:PUGB4, pass, PENB
			10'd210 : rdata = 48'b110001110000100100000000000000000000000100000000;
			// PEs: 53 -> 56
			// srcs: (382, 264)(2733) 0 --> (2733) 0:PEGB5, pass, PUNB
			10'd211 : rdata = 48'b110001110000101000000000000000000000001000000000;
			// PEs: 52 -> 32
			// srcs: (386, 258)(2658) 2 --> (2658) 2:PEGB4, pass, PUGB4
			10'd212 : rdata = 48'b110001110000100000000000000000000000000000001100;
			// PEs: 48 -> 49
			// srcs: (387, 180)(2691) -2 --> (2691) -2:NI0, pass, PENB
			10'd213 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 16 -> 48
			// srcs: (388, 185)(2767) 2 --> (2767) 2:PUGB2, pass, NI0
			10'd214 : rdata = 48'b110001110000010100000000000100000000000000000000;
			// PEs: 56 -> 49
			// srcs: (389, 186)(1989) 4 --> (1989) 4:PUGB7, pass, PENB
			10'd215 : rdata = 48'b110001110000111100000000000000000000000100000000;
			// PEs: 48 -> 49
			// srcs: (395, 187)(2767) 2 --> (2767) 2:NI0, pass, PENB
			10'd216 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 24 -> 48
			// srcs: (396, 188)(2785) 4 --> (2785) 4:PUGB3, pass, NI0
			10'd217 : rdata = 48'b110001110000011100000000000100000000000000000000;
			// PEs: 0 -> 49
			// srcs: (397, 189)(2007) 0 --> (2007) 0:PUGB0, pass, PENB
			10'd218 : rdata = 48'b110001110000000100000000000000000000000100000000;
			// PEs: 49 -> 16
			// srcs: (402, 265)(2768) 6 --> (2768) 6:PEGB1, pass, PUGB2
			10'd219 : rdata = 48'b110001110000001000000000000000000000000000001010;
			// PEs: 48 -> 49
			// srcs: (403, 190)(2785) 4 --> (2785) 4:NI0, pass, PENB
			10'd220 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 40 -> 48
			// srcs: (404, 191)(2804) 0 --> (2804) 0:PUNB, pass, NI0
			10'd221 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 8 -> 49
			// srcs: (405, 192)(2026) -1 --> (2026) -1:PUGB1, pass, PENB
			10'd222 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 49 -> 56
			// srcs: (410, 266)(2786) 4 --> (2786) 4:PEGB1, pass, PUNB
			10'd223 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 48 -> 49
			// srcs: (411, 193)(2804) 0 --> (2804) 0:NI0, pass, PENB
			10'd224 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 0 -> 49
			// srcs: (412, 198)(2910) 0 --> (2910) 0:PUGB0, pass, PENB
			10'd225 : rdata = 48'b110001110000000100000000000000000000000100000000;
			// PEs: 0 -> 49
			// srcs: (413, 199)(2912) -1 --> (2912) -1:PUGB0, pass, PENB
			10'd226 : rdata = 48'b110001110000000100000000000000000000000100000000;
			// PEs: 8 -> 49
			// srcs: (414, 200)(2917) 0 --> (2917) 0:PUGB1, pass, PENB
			10'd227 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 49
			// srcs: (415, 203)(2924) -3 --> (2924) -3:PUGB1, pass, PENB
			10'd228 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 24 -> 48
			// srcs: (416, 205)(2935) -3 --> (2935) -3:PUGB3, pass, NI0
			10'd229 : rdata = 48'b110001110000011100000000000100000000000000000000;
			// PEs: 50 -> 56
			// srcs: (417, 272)(2895) 13 --> (2895) 13:PEGB2, pass, PUNB
			10'd230 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 49 -> 32
			// srcs: (429, 274)(2925) -3 --> (2925) -3:PEGB1, pass, PUGB4
			10'd231 : rdata = 48'b110001110000001000000000000000000000000000001100;
			// PEs: 40 -> 51
			// srcs: (440, 197)(2111) 0 --> (2111) 0:PUNB, pass, PEGB3
			10'd232 : rdata = 48'b110001101111111100000000000000000000000010110000;
			// PEs: 56 -> 49
			// srcs: (531, 206)(2160) 4 --> (2160) 4:PUGB7, pass, PENB
			10'd233 : rdata = 48'b110001110000111100000000000000000000000100000000;
			// PEs: 48 -> 49
			// srcs: (537, 207)(2935) -3 --> (2935) -3:NI0, pass, PENB
			10'd234 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 40 -> 48
			// srcs: (538, 208)(2957) 3 --> (2957) 3:PUNB, pass, NI0
			10'd235 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 0 -> 49
			// srcs: (539, 209)(2179) -3 --> (2179) -3:PUGB0, pass, PENB
			10'd236 : rdata = 48'b110001110000000100000000000000000000000100000000;
			// PEs: 48 -> 49
			// srcs: (545, 210)(2957) 3 --> (2957) 3:NI0, pass, PENB
			10'd237 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 0 -> 49
			// srcs: (546, 211)(2191) 6 --> (2191) 6:PUGB0, pass, PENB
			10'd238 : rdata = 48'b110001110000000100000000000000000000000100000000;
			// PEs: 0 -> 49
			// srcs: (547, 213)(2197) 0 --> (2197) 0:PUGB0, pass, PENB
			10'd239 : rdata = 48'b110001110000000100000000000000000000000100000000;
			// PEs: 40 -> 48
			// srcs: (548, 214)(3046) 1 --> (3046) 1:PUNB, pass, NI0
			10'd240 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 24 -> 49
			// srcs: (549, 215)(2268) 1 --> (2268) 1:PUGB3, pass, PENB
			10'd241 : rdata = 48'b110001110000011100000000000000000000000100000000;
			// PEs: 49 -> 8
			// srcs: (552, 276)(2958) 0 --> (2958) 0:PEGB1, pass, PUGB1
			10'd242 : rdata = 48'b110001110000001000000000000000000000000000001001;
			// PEs: 49 -> 56
			// srcs: (553, 277)(2970) 2 --> (2970) 2:PEGB1, pass, PUNB
			10'd243 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 49 -> 32
			// srcs: (554, 278)(2975) 0 --> (2975) 0:PEGB1, pass, PUGB4
			10'd244 : rdata = 48'b110001110000001000000000000000000000000000001100;
			// PEs: 48 -> 49
			// srcs: (555, 216)(3046) 1 --> (3046) 1:NI0, pass, PENB
			10'd245 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 56 -> 48
			// srcs: (556, 220)(3069) 6 --> (3069) 6:PUGB7, pass, NI0
			10'd246 : rdata = 48'b110001110000111100000000000100000000000000000000;
			// PEs: 40 -> 49
			// srcs: (557, 221)(2292) -2 --> (2292) -2:PUNB, pass, PENB
			10'd247 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 48 -> 49
			// srcs: (563, 222)(3069) 6 --> (3069) 6:NI0, pass, PENB
			10'd248 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 0 -> 48
			// srcs: (564, 223)(3082) -4 --> (3082) -4:PUGB0, pass, NI0
			10'd249 : rdata = 48'b110001110000000100000000000100000000000000000000;
			// PEs: 40 -> 49
			// srcs: (565, 224)(2307) 2 --> (2307) 2:PUNB, pass, PENB
			10'd250 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 49 -> 32
			// srcs: (570, 280)(3070) 4 --> (3070) 4:PEGB1, pass, PUGB4
			10'd251 : rdata = 48'b110001110000001000000000000000000000000000001100;
			// PEs: 48 -> 49
			// srcs: (571, 225)(3082) -4 --> (3082) -4:NI0, pass, PENB
			10'd252 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 24 -> 49
			// srcs: (572, 231)(3107) -6 --> (3107) -6:PUGB3, pass, PENB
			10'd253 : rdata = 48'b110001110000011100000000000000000000000100000000;
			// PEs: 0 -> 48
			// srcs: (573, 234)(2364) -11 --> (2364) -11:PUGB0, pass, NI0
			10'd254 : rdata = 48'b110001110000000100000000000100000000000000000000;
			// PEs: 16 -> 49
			// srcs: (574, 235)(2366) -11 --> (2366) -11:PUGB2, pass, PENB
			10'd255 : rdata = 48'b110001110000010100000000000000000000000100000000;
			// PEs: 49 -> 40
			// srcs: (578, 281)(3083) -2 --> (3083) -2:PEGB1, pass, PUGB5
			10'd256 : rdata = 48'b110001110000001000000000000000000000000000001101;
			// PEs: 48 -> 49
			// srcs: (585, 236)(2364) -11 --> (2364) -11:NI0, pass, PENB
			10'd257 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 40 -> 48
			// srcs: (586, 240)(2412) 0 --> (2412) 0:PUNB, pass, NI0
			10'd258 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 8 -> 49
			// srcs: (587, 241)(2414) -3 --> (2414) -3:PUGB1, pass, PENB
			10'd259 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 40 -> 54
			// srcs: (588, 256)(2636) 2 --> (2636) 2:PUNB, pass, PEGB6
			10'd260 : rdata = 48'b110001101111111100000000000000000000000011100000;
			// PEs: 40 -> 51
			// srcs: (589, 259)(2667) -10 --> (2667) -10:PUNB, pass, PEGB3
			10'd261 : rdata = 48'b110001101111111100000000000000000000000010110000;
			// PEs: 40 -> 52
			// srcs: (590, 263)(2690) 1 --> (2690) 1:PUNB, pass, PEGB4
			10'd262 : rdata = 48'b110001101111111100000000000000000000000011000000;
			// PEs: 49 -> 56
			// srcs: (591, 282)(3108) -9 --> (3108) -9:PEGB1, pass, PUNB
			10'd263 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 49 -> 40
			// srcs: (592, 283)(2367) -22 --> (2367) -22:PEGB1, pass, PUGB5
			10'd264 : rdata = 48'b110001110000001000000000000000000000000000001101;
			// PEs: 48 -> 49
			// srcs: (593, 242)(2412) 0 --> (2412) 0:NI0, pass, PENB
			10'd265 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 24 -> 48
			// srcs: (594, 245)(2467) 0 --> (2467) 0:PUGB3, pass, NI0
			10'd266 : rdata = 48'b110001110000011100000000000100000000000000000000;
			// PEs: 56 -> 49
			// srcs: (595, 246)(2469) -5 --> (2469) -5:PUGB7, pass, PENB
			10'd267 : rdata = 48'b110001110000111100000000000000000000000100000000;
			// PEs: 49 -> 32
			// srcs: (600, 287)(2415) -3 --> (2415) -3:PEGB1, pass, PUGB4
			10'd268 : rdata = 48'b110001110000001000000000000000000000000000001100;
			// PEs: 48 -> 49
			// srcs: (601, 247)(2467) 0 --> (2467) 0:NI0, pass, PENB
			10'd269 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 32 -> 49
			// srcs: (602, 252)(2554) -1 --> (2554) -1:PUGB4, pass, PENB
			10'd270 : rdata = 48'b110001110000100100000000000000000000000100000000;
			// PEs: 16 -> 48
			// srcs: (603, 253)(2618) -2 --> (2618) -2:PUGB2, pass, NI0
			10'd271 : rdata = 48'b110001110000010100000000000100000000000000000000;
			// PEs: 56 -> 49
			// srcs: (604, 254)(2620) 1 --> (2620) 1:PUGB7, pass, PENB
			10'd272 : rdata = 48'b110001110000111100000000000000000000000100000000;
			// PEs: 55 -> 56
			// srcs: (605, 292)(2568) 8 --> (2568) 8:PENB, pass, PUNB
			10'd273 : rdata = 48'b110001101111111000000000000000000000001000000000;
			// PEs: 51 -> 0
			// srcs: (606, 295)(2670) -10 --> (2670) -10:PEGB3, pass, PUGB0
			10'd274 : rdata = 48'b110001110000011000000000000000000000000000001000;
			// PEs: 52 -> 16
			// srcs: (607, 297)(2693) -1 --> (2693) -1:PEGB4, pass, PUGB2
			10'd275 : rdata = 48'b110001110000100000000000000000000000000000001010;
			// PEs: 50 -> 16
			// srcs: (608, 302)(2914) -9 --> (2914) -9:PEGB2, pass, PUGB2
			10'd276 : rdata = 48'b110001110000010000000000000000000000000000001010;
			// PEs: 48 -> 49
			// srcs: (610, 255)(2618) -2 --> (2618) -2:NI0, pass, PENB
			10'd277 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 16 -> 48
			// srcs: (611, 260)(2679) 4 --> (2679) 4:PUGB2, pass, NI0
			10'd278 : rdata = 48'b110001110000010100000000000100000000000000000000;
			// PEs: 0 -> 49
			// srcs: (612, 261)(2681) -5 --> (2681) -5:PUGB0, pass, PENB
			10'd279 : rdata = 48'b110001110000000100000000000000000000000100000000;
			// PEs: 49 -> 56
			// srcs: (617, 293)(2621) -1 --> (2621) -1:PEGB1, pass, PUNB
			10'd280 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 48 -> 49
			// srcs: (618, 262)(2679) 4 --> (2679) 4:NI0, pass, PENB
			10'd281 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 16 -> 49
			// srcs: (619, 267)(2803) 3 --> (2803) 3:PUGB2, pass, PENB
			10'd282 : rdata = 48'b110001110000010100000000000000000000000100000000;
			// PEs: 32 -> 48
			// srcs: (620, 268)(2814) 9 --> (2814) 9:PUGB4, pass, NI0
			10'd283 : rdata = 48'b110001110000100100000000000100000000000000000000;
			// PEs: 0 -> 49
			// srcs: (621, 269)(2816) -3 --> (2816) -3:PUGB0, pass, PENB
			10'd284 : rdata = 48'b110001110000000100000000000000000000000100000000;
			// PEs: 49 -> 56
			// srcs: (625, 296)(2682) -1 --> (2682) -1:PEGB1, pass, PUNB
			10'd285 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 49 -> 24
			// srcs: (626, 299)(2806) 2 --> (2806) 2:PEGB1, pass, PUGB3
			10'd286 : rdata = 48'b110001110000001000000000000000000000000000001011;
			// PEs: 48 -> 49
			// srcs: (627, 270)(2814) 9 --> (2814) 9:NI0, pass, PENB
			10'd287 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 40 -> 49
			// srcs: (661, 271)(2886) -9 --> (2886) -9:PUNB, pass, PENB
			10'd288 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 40 -> 49
			// srcs: (662, 273)(2920) -2 --> (2920) -2:PUNB, pass, PENB
			10'd289 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 40 -> 49
			// srcs: (663, 275)(2934) 8 --> (2934) 8:PUNB, pass, PENB
			10'd290 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 49 -> 24
			// srcs: (669, 303)(2921) -1 --> (2921) -1:PEGB1, pass, PUGB3
			10'd291 : rdata = 48'b110001110000001000000000000000000000000000001011;
			// PEs: 49 -> 56
			// srcs: (670, 304)(2937) 9 --> (2937) 9:PEGB1, pass, PUNB
			10'd292 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 40 -> 49
			// srcs: (674, 279)(3049) -2 --> (3049) -2:PUNB, pass, PENB
			10'd293 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 8 -> 48
			// srcs: (675, 284)(2385) -3 --> (2385) -3:PUGB1, pass, NI0
			10'd294 : rdata = 48'b110001110000001100000000000100000000000000000000;
			// PEs: 32 -> 49
			// srcs: (676, 285)(2390) 7 --> (2390) 7:PUGB4, pass, PENB
			10'd295 : rdata = 48'b110001110000100100000000000000000000000100000000;
			// PEs: 48 -> 49
			// srcs: (682, 286)(2385) -3 --> (2385) -3:NI0, pass, PENB
			10'd296 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 0 -> 49
			// srcs: (683, 288)(2475) 12 --> (2475) 12:PUGB0, pass, PENB
			10'd297 : rdata = 48'b110001110000000100000000000000000000000100000000;
			// PEs: 49 -> 32
			// srcs: (689, 306)(2391) 4 --> (2391) 4:PEGB1, pass, PUGB4
			10'd298 : rdata = 48'b110001110000001000000000000000000000000000001100;
			// PEs: 49 -> 56
			// srcs: (690, 310)(2476) 7 --> (2476) 7:PEGB1, pass, PUNB
			10'd299 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 50 -> 56
			// srcs: (691, 312)(2563) 3 --> (2563) 3:PEGB2, pass, PUNB
			10'd300 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 24 -> 48
			// srcs: (725, 289)(2541) -7 --> (2541) -7:PUGB3, pass, NI0
			10'd301 : rdata = 48'b110001110000011100000000000100000000000000000000;
			// PEs: 40 -> 49
			// srcs: (741, 290)(2546) -5 --> (2546) -5:PUNB, pass, PENB
			10'd302 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 48 -> 49
			// srcs: (751, 291)(2541) -7 --> (2541) -7:NI0, pass, PENB
			10'd303 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 40 -> 49
			// srcs: (752, 294)(2644) 2 --> (2644) 2:PUNB, pass, PENB
			10'd304 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 49 -> 0
			// srcs: (758, 311)(2547) -12 --> (2547) -12:PEGB1, pass, PUGB0
			10'd305 : rdata = 48'b110001110000001000000000000000000000000000001000;
			// PEs: 49 -> 32
			// srcs: (759, 313)(2645) 2 --> (2645) 2:PEGB1, pass, PUGB4
			10'd306 : rdata = 48'b110001110000001000000000000000000000000000001100;
			// PEs: 40 -> 49
			// srcs: (1377, 298)(2725) 4 --> (2725) 4:PUNB, pass, PENB
			10'd307 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 40 -> 49
			// srcs: (1378, 300)(2812) -9 --> (2812) -9:PUNB, pass, PENB
			10'd308 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 40 -> 49
			// srcs: (1379, 301)(2884) 2 --> (2884) 2:PUNB, pass, PENB
			10'd309 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 32 -> 49
			// srcs: (1380, 305)(3045) -9 --> (3045) -9:PUGB4, pass, PENB
			10'd310 : rdata = 48'b110001110000100100000000000000000000000100000000;
			// PEs: 32 -> 48
			// srcs: (1381, 307)(2439) 10 --> (2439) 10:PUGB4, pass, NI0
			10'd311 : rdata = 48'b110001110000100100000000000100000000000000000000;
			// PEs: 8 -> 49
			// srcs: (1382, 308)(2450) 8 --> (2450) 8:PUGB1, pass, PENB
			10'd312 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 49 -> 56
			// srcs: (1391, 317)(2731) 18 --> (2731) 18:PEGB1, pass, PUNB
			10'd313 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 49 -> 8
			// srcs: (1392, 318)(2818) -3 --> (2818) -3:PEGB1, pass, PUGB1
			10'd314 : rdata = 48'b110001110000001000000000000000000000000000001001;
			// PEs: 48 -> 49
			// srcs: (1393, 309)(2439) 10 --> (2439) 10:NI0, pass, PENB
			10'd315 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 56 -> 48
			// srcs: (1394, 314)(2683) -4 --> (2683) -4:PUGB7, pass, NI0
			10'd316 : rdata = 48'b110001110000111100000000000100000000000000000000;
			// PEs: 16 -> 49
			// srcs: (1395, 315)(2694) -4 --> (2694) -4:PUGB2, pass, PENB
			10'd317 : rdata = 48'b110001110000010100000000000000000000000100000000;
			// PEs: 49 -> 56
			// srcs: (1396, 320)(3051) -9 --> (3051) -9:PEGB1, pass, PUNB
			10'd318 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 48 -> 49
			// srcs: (1401, 316)(2683) -4 --> (2683) -4:NI0, pass, PENB
			10'd319 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 40 -> 49
			// srcs: (1402, 319)(2879) 12 --> (2879) 12:PUNB, pass, PENB
			10'd320 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 40 -> 49
			// srcs: (1403, 321)(2428) -4 --> (2428) -4:PUNB, pass, PENB
			10'd321 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 40 -> 49
			// srcs: (1404, 322)(2672) -6 --> (2672) -6:PUNB, pass, PENB
			10'd322 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 40 -> 49
			// srcs: (1405, 323)(2868) 11 --> (2868) 11:PUNB, pass, PENB
			10'd323 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 49 -> 24
			// srcs: (1410, 324)(2452) 14 --> (2452) 14:PEGB1, pass, PUGB3
			10'd324 : rdata = 48'b110001110000001000000000000000000000000000001011;
			// PEs: 8 -> 48
			// srcs: (1418, 325)(2599) 4 --> (2599) 4:PUGB1, pass, NI0
			10'd325 : rdata = 48'b110001110000001100000000000100000000000000000000;
			// PEs: 40 -> 49
			// srcs: (1419, 326)(2647) 48 --> (2647) 48:PUNB, pass, PENB
			10'd326 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 49 -> 56
			// srcs: (1420, 328)(2696) -14 --> (2696) -14:PEGB1, pass, PUNB
			10'd327 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 49 -> 24
			// srcs: (1421, 329)(2892) 28 --> (2892) 28:PEGB1, pass, PUGB3
			10'd328 : rdata = 48'b110001110000001000000000000000000000000000001011;
			// PEs: 48 -> 49
			// srcs: (1425, 327)(2599) 4 --> (2599) 4:NI0, pass, PENB
			10'd329 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 49 -> 56
			// srcs: (1432, 330)(2648) 52 --> (2648) 52:PEGB1, pass, PUNB
			10'd330 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 24 -> 48
			// srcs: (1458, 331)(2942) 24 --> (2942) 24:PUGB3, pass, NI0
			10'd331 : rdata = 48'b110001110000011100000000000100000000000000000000;
			// PEs: 40 -> 49
			// srcs: (1463, 332)(3137) -63 --> (3137) -63:PUNB, pass, PENB
			10'd332 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 48 -> 49
			// srcs: (1473, 333)(2942) 24 --> (2942) 24:NI0, pass, PENB
			10'd333 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 49 -> 8
			// srcs: (1480, 334)(3138) -39 --> (3138) -39:PEGB1, pass, PUGB1
			10'd334 : rdata = 48'b110001110000001000000000000000000000000000001001;
			// PEs: 8 -> 49
			// srcs: (1521, 335)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd335 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 50
			// srcs: (1524, 336)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd336 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 51
			// srcs: (1527, 337)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd337 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 52
			// srcs: (1530, 338)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd338 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 53
			// srcs: (1533, 339)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd339 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 54
			// srcs: (1536, 340)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd340 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 55
			// srcs: (1539, 341)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd341 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 49
			// srcs: (1568, 342)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd342 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 50
			// srcs: (1569, 343)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd343 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 51
			// srcs: (1571, 344)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd344 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 52
			// srcs: (1572, 345)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd345 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 53
			// srcs: (1574, 346)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd346 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 54
			// srcs: (1575, 347)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd347 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 55
			// srcs: (1577, 348)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd348 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 49
			// srcs: (1650, 349)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd349 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 50
			// srcs: (1651, 350)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd350 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 51
			// srcs: (1653, 351)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd351 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 52
			// srcs: (1654, 352)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd352 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 53
			// srcs: (1656, 353)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd353 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 54
			// srcs: (1657, 354)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd354 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 55
			// srcs: (1658, 355)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd355 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 49
			// srcs: (1701, 356)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd356 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 50
			// srcs: (1704, 357)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd357 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 51
			// srcs: (1711, 358)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd358 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 52
			// srcs: (1714, 359)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd359 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 53
			// srcs: (1717, 360)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd360 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 54
			// srcs: (1720, 361)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd361 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 55
			// srcs: (1723, 362)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd362 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 49
			// srcs: (1730, 363)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd363 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 50
			// srcs: (1731, 364)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd364 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 51
			// srcs: (1733, 365)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd365 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 52
			// srcs: (1734, 366)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd366 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 53
			// srcs: (1736, 367)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd367 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 54
			// srcs: (1737, 368)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd368 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 55
			// srcs: (1739, 369)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd369 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 49
			// srcs: (1810, 370)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd370 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 50
			// srcs: (1811, 371)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd371 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 51
			// srcs: (1813, 372)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd372 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 52
			// srcs: (1814, 373)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd373 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 53
			// srcs: (1816, 374)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd374 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 54
			// srcs: (1817, 375)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd375 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 55
			// srcs: (1819, 376)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd376 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 49
			// srcs: (1885, 377)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd377 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 50
			// srcs: (1888, 378)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd378 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 51
			// srcs: (1891, 379)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd379 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 49
			// srcs: (1892, 380)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd380 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 50
			// srcs: (1893, 381)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd381 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 52
			// srcs: (1894, 382)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd382 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 51
			// srcs: (1895, 383)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd383 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 52
			// srcs: (1896, 384)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd384 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 53
			// srcs: (1897, 385)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd385 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 53
			// srcs: (1898, 386)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd386 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 54
			// srcs: (1899, 387)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd387 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 54
			// srcs: (1900, 388)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd388 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 55
			// srcs: (1901, 389)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd389 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 55
			// srcs: (1907, 390)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd390 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 49
			// srcs: (1972, 391)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd391 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 50
			// srcs: (1973, 392)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd392 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 51
			// srcs: (1975, 393)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd393 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 52
			// srcs: (1976, 394)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd394 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 53
			// srcs: (1978, 395)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd395 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 54
			// srcs: (1979, 396)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd396 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 55
			// srcs: (1981, 397)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd397 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 49
			// srcs: (2052, 398)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd398 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 50
			// srcs: (2053, 399)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd399 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 51
			// srcs: (2055, 400)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd400 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 52
			// srcs: (2056, 401)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd401 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 53
			// srcs: (2058, 402)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd402 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 54
			// srcs: (2059, 403)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd403 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 55
			// srcs: (2061, 404)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd404 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 49
			// srcs: (2069, 405)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd405 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 50
			// srcs: (2072, 406)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd406 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 51
			// srcs: (2075, 407)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd407 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 52
			// srcs: (2078, 408)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd408 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 53
			// srcs: (2081, 409)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd409 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 54
			// srcs: (2084, 410)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd410 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 55
			// srcs: (2087, 411)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd411 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 49
			// srcs: (2134, 412)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd412 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 50
			// srcs: (2135, 413)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd413 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 51
			// srcs: (2137, 414)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd414 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 52
			// srcs: (2138, 415)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd415 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 53
			// srcs: (2140, 416)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd416 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 54
			// srcs: (2141, 417)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd417 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 55
			// srcs: (2143, 418)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd418 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 49
			// srcs: (2214, 419)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd419 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 50
			// srcs: (2215, 420)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd420 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 51
			// srcs: (2217, 421)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd421 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 52
			// srcs: (2218, 422)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd422 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 53
			// srcs: (2220, 423)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd423 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 54
			// srcs: (2221, 424)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd424 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 55
			// srcs: (2223, 425)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd425 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 49
			// srcs: (2253, 426)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd426 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 50
			// srcs: (2256, 427)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd427 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 51
			// srcs: (2259, 428)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd428 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 52
			// srcs: (2262, 429)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd429 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 53
			// srcs: (2265, 430)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd430 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 54
			// srcs: (2268, 431)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd431 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 55
			// srcs: (2271, 432)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd432 : rdata = 48'b110001110000001100000000000000000000000011110000;
			default : rdata = 48'b000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 49) begin
	always @(*) begin
		case(address)
			// PEs: 49, 49 -> 48
			// srcs: (1, 0)(63) 0, (848) 2 --> (1632) 0:ND0, NW0, *, PEGB0
			10'd0 : rdata = 48'b000110110000000001000000000000000000000010000000;
			// PEs: 49, 49 -> 48
			// srcs: (2, 1)(145) -3, (930) -3 --> (1714) 9:ND1, NW1, *, PEGB0
			10'd1 : rdata = 48'b000110110000000101000000001000000000000010000000;
			// PEs: 49, 49 -> 48
			// srcs: (3, 2)(225) -2, (1010) 0 --> (1794) 0:ND2, NW2, *, PEGB0
			10'd2 : rdata = 48'b000110110000001001000000010000000000000010000000;
			// PEs: 49, 49 -> 48
			// srcs: (4, 3)(305) 1, (1090) -2 --> (1874) -2:ND3, NW3, *, PEGB0
			10'd3 : rdata = 48'b000110110000001101000000011000000000000010000000;
			// PEs: 49, 49 -> 48
			// srcs: (5, 4)(387) 2, (1172) -1 --> (1956) -2:ND4, NW4, *, PEGB0
			10'd4 : rdata = 48'b000110110000010001000000100000000000000010000000;
			// PEs: 49, 49 -> 48
			// srcs: (6, 5)(467) 0, (1252) 1 --> (2036) 0:ND5, NW5, *, PEGB0
			10'd5 : rdata = 48'b000110110000010101000000101000000000000010000000;
			// PEs: 49, 49 -> 48
			// srcs: (7, 6)(547) -1, (1332) 2 --> (2116) -2:ND6, NW6, *, PEGB0
			10'd6 : rdata = 48'b000110110000011001000000110000000000000010000000;
			// PEs: 49, 49 -> 48
			// srcs: (8, 7)(629) 2, (1414) 0 --> (2198) 0:ND7, NW7, *, PEGB0
			10'd7 : rdata = 48'b000110110000011101000000111000000000000010000000;
			// PEs: 49, 49 -> 52
			// srcs: (9, 8)(709) 1, (1494) -1 --> (2278) -1:ND8, NW8, *, PEGB4
			10'd8 : rdata = 48'b000110110000100001000001000000000000000011000000;
			// PEs: 49, 49 -> 48
			// srcs: (10, 9)(16) -3, (801) 1 --> (1585) -3:ND9, NW9, *, PEGB0
			10'd9 : rdata = 48'b000110110000100101000001001000000000000010000000;
			// PEs: 49, 49 -> 48
			// srcs: (11, 10)(196) 0, (981) -3 --> (1765) 0:ND10, NW10, *, PEGB0
			10'd10 : rdata = 48'b000110110000101001000001010000000000000010000000;
			// PEs: 49, 49 -> 49
			// srcs: (12, 11)(380) -2, (1165) -3 --> (1949) 6:ND11, NW11, *, NI0
			10'd11 : rdata = 48'b000110110000101101000001011100000000000000000000;
			// PEs: 49, 49 -> 49
			// srcs: (13, 12)(564) 2, (1349) -1 --> (2133) -2:ND12, NW12, *, NI1
			10'd12 : rdata = 48'b000110110000110001000001100100001000000000000000;
			// PEs: 49, 49 -> 49
			// srcs: (14, 13)(748) 2, (1533) 0 --> (2317) 0:ND13, NW13, *, NI2
			10'd13 : rdata = 48'b000110110000110101000001101100010000000000000000;
			// PEs: 48 -> 
			// srcs: (42, 14)(1669) 0 --> (1669) 0:PENB, pass, 
			10'd14 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 48, 49 -> 49
			// srcs: (48, 15)(1668) 9, (1669) 0 --> (2447) 9:PENB, ALU, +, NI3
			10'd15 : rdata = 48'b000011101111111000111111111100011000000000000000;
			// PEs: 55, 48 -> 48
			// srcs: (54, 16)(1883) -1, (1884) -1 --> (2663) -2:PEGB7, PENB, +, PEGB0
			10'd16 : rdata = 48'b000011110000111011011111110000000000000010000000;
			// PEs: 48 -> 
			// srcs: (59, 17)(1887) -2 --> (1887) -2:PENB, pass, 
			10'd17 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 48, 49 -> 48
			// srcs: (65, 18)(1886) -6, (1887) -2 --> (2666) -8:PENB, ALU, +, PEGB0
			10'd18 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 48 -> 
			// srcs: (68, 19)(1948) -2 --> (1948) -2:PENB, pass, 
			10'd19 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 48, 49 -> 50
			// srcs: (74, 20)(1947) 1, (1948) -2 --> (2726) -1:PENB, ALU, +, PENB
			10'd20 : rdata = 48'b000011101111111000111111111000000000000100000000;
			// PEs: 48 -> 49
			// srcs: (76, 21)(1951) 6 --> (1951) 6:PENB, pass, NI4
			10'd21 : rdata = 48'b110001101111111000000000000100100000000000000000;
			// PEs: 49 -> 50
			// srcs: (81, 67)(1949) 6 --> (1949) 6:NI0, pass, PENB
			10'd22 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 48, 49 -> 50
			// srcs: (82, 22)(1950) 9, (1951) 6 --> (2728) 15:PENB, NI4, +, PENB
			10'd23 : rdata = 48'b000011101111111010100000100000000000000100000000;
			// PEs: 48 -> 
			// srcs: (84, 23)(1954) 3 --> (1954) 3:PENB, pass, 
			10'd24 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 48, 49 -> 53
			// srcs: (90, 24)(1953) -3, (1954) 3 --> (2732) 0:PENB, ALU, +, PEGB5
			10'd25 : rdata = 48'b000011101111111000111111111000000000000011010000;
			// PEs: 48 -> 
			// srcs: (92, 25)(2028) 0 --> (2028) 0:PENB, pass, 
			10'd26 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 48, 49 -> 48
			// srcs: (98, 26)(2027) -6, (2028) 0 --> (2808) -6:PENB, ALU, +, PEGB0
			10'd27 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 48 -> 
			// srcs: (100, 27)(2031) -2 --> (2031) -2:PENB, pass, 
			10'd28 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 48, 49 -> 48
			// srcs: (106, 28)(2030) -1, (2031) -2 --> (2810) -3:PENB, ALU, +, PEGB0
			10'd29 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 48 -> 
			// srcs: (108, 29)(2034) 1 --> (2034) 1:PENB, pass, 
			10'd30 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 48, 49 -> 48
			// srcs: (114, 30)(2033) 9, (2034) 1 --> (2813) 10:PENB, ALU, +, PEGB0
			10'd31 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 48 -> 
			// srcs: (116, 31)(2110) 6 --> (2110) 6:PENB, pass, 
			10'd32 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 48, 49 -> 51
			// srcs: (122, 32)(2109) 6, (2110) 6 --> (2887) 12:PENB, ALU, +, PEGB3
			10'd33 : rdata = 48'b000011101111111000111111111000000000000010110000;
			// PEs: 48 -> 
			// srcs: (124, 33)(2190) -2 --> (2190) -2:PENB, pass, 
			10'd34 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 48, 49 -> 49
			// srcs: (130, 34)(2189) -2, (2190) -2 --> (2969) -4:PENB, ALU, +, NI0
			10'd35 : rdata = 48'b000011101111111000111111111100000000000000000000;
			// PEs: 48 -> 
			// srcs: (132, 35)(2193) -6 --> (2193) -6:PENB, pass, 
			10'd36 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 48, 49 -> 48
			// srcs: (138, 36)(2192) -3, (2193) -6 --> (2972) -9:PENB, ALU, +, PEGB0
			10'd37 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 48 -> 
			// srcs: (140, 37)(2196) 2 --> (2196) 2:PENB, pass, 
			10'd38 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 48, 49 -> 49
			// srcs: (146, 38)(2195) -2, (2196) 2 --> (2974) 0:PENB, ALU, +, NI4
			10'd39 : rdata = 48'b000011101111111000111111111100100000000000000000;
			// PEs: 49 -> 48
			// srcs: (169, 91)(2317) 0 --> (2317) 0:NI2, pass, PEGB0
			10'd40 : rdata = 48'b110001010000001000000000000000000000000010000000;
			// PEs: 48 -> 
			// srcs: (282, 39)(2113) -1 --> (2113) -1:PENB, pass, 
			10'd41 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 48, 49 -> 49
			// srcs: (288, 40)(2112) 9, (2113) -1 --> (2893) 8:PENB, ALU, +, NI2
			10'd42 : rdata = 48'b000011101111111000111111111100010000000000000000;
			// PEs: 48 -> 
			// srcs: (311, 41)(2115) 3 --> (2115) 3:PENB, pass, 
			10'd43 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 48, 49 -> 50
			// srcs: (317, 42)(2114) 2, (2115) 3 --> (2894) 5:PENB, ALU, +, PENB
			10'd44 : rdata = 48'b000011101111111000111111111000000000000100000000;
			// PEs: 54, 48 -> 48
			// srcs: (318, 43)(2357) 9, (2358) 0 --> (2359) 9:PEGB6, PENB, +, PEGB0
			10'd45 : rdata = 48'b000011110000110011011111110000000000000010000000;
			// PEs: 48, 51 -> 48
			// srcs: (319, 44)(2371) 9, (1591) 2 --> (2372) 11:PENB, PEGB3, +, PEGB0
			10'd46 : rdata = 48'b000011101111111011100000110000000000000010000000;
			// PEs: 48, 53 -> 48
			// srcs: (320, 45)(2376) -6, (1597) 0 --> (2377) -6:PENB, PEGB5, +, PEGB0
			10'd47 : rdata = 48'b000011101111111011100001010000000000000010000000;
			// PEs: 48 -> 49
			// srcs: (322, 46)(1621) 2 --> (1621) 2:PENB, pass, NI5
			10'd48 : rdata = 48'b110001101111111000000000000100101000000000000000;
			// PEs: 49 -> 50
			// srcs: (324, 74)(2893) 8 --> (2893) 8:NI2, pass, PENB
			10'd49 : rdata = 48'b110001010000001000000000000000000000000100000000;
			// PEs: 48, 49 -> 48
			// srcs: (328, 47)(2399) 0, (1621) 2 --> (2400) 2:PENB, NI5, +, PEGB0
			10'd50 : rdata = 48'b000011101111111010100000101000000000000010000000;
			// PEs: 48 -> 
			// srcs: (330, 48)(1661) 0 --> (1661) 0:PENB, pass, 
			10'd51 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 48, 49 -> 48
			// srcs: (336, 49)(2440) 2, (1661) 0 --> (2441) 2:PENB, ALU, +, PEGB0
			10'd52 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 49, 48 -> 48
			// srcs: (337, 50)(2447) 9, (1670) -6 --> (2448) 3:NI3, PENB, +, PEGB0
			10'd53 : rdata = 48'b000011010000001111011111110000000000000010000000;
			// PEs: 48 -> 
			// srcs: (339, 51)(1695) 3 --> (1695) 3:PENB, pass, 
			10'd54 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 48, 49 -> 48
			// srcs: (345, 52)(2473) -6, (1695) 3 --> (2474) -3:PENB, ALU, +, PEGB0
			10'd55 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 48 -> 
			// srcs: (347, 53)(1729) -3 --> (1729) -3:PENB, pass, 
			10'd56 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 48, 49 -> 48
			// srcs: (353, 54)(2508) 6, (1729) -3 --> (2509) 3:PENB, ALU, +, PEGB0
			10'd57 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 48 -> 
			// srcs: (355, 55)(1756) -2 --> (1756) -2:PENB, pass, 
			10'd58 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 48, 49 -> 48
			// srcs: (361, 56)(2533) -4, (1756) -2 --> (2534) -6:PENB, ALU, +, PEGB0
			10'd59 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 48, 50 -> 48
			// srcs: (362, 57)(2544) -3, (1768) -2 --> (2545) -5:PENB, PEGB2, +, PEGB0
			10'd60 : rdata = 48'b000011101111111011100000100000000000000010000000;
			// PEs: 48, 51 -> 49
			// srcs: (363, 58)(2555) 1, (1775) 0 --> (2556) 1:PENB, PEGB3, +, NI2
			10'd61 : rdata = 48'b000011101111111011100000110100010000000000000000;
			// PEs: 48, 52 -> 49
			// srcs: (364, 59)(2558) 11, (1778) -6 --> (2559) 5:PENB, PEGB4, +, NI3
			10'd62 : rdata = 48'b000011101111111011100001000100011000000000000000;
			// PEs: 48, 53 -> 50
			// srcs: (365, 60)(2560) -6, (1781) 4 --> (2561) -2:PENB, PEGB5, +, PENB
			10'd63 : rdata = 48'b000011101111111011100001010000000000000100000000;
			// PEs: 48 -> 49
			// srcs: (367, 61)(1860) 0 --> (1860) 0:PENB, pass, NI5
			10'd64 : rdata = 48'b110001101111111000000000000100101000000000000000;
			// PEs: 49 -> 50
			// srcs: (372, 100)(2559) 5 --> (2559) 5:NI3, pass, PENB
			10'd65 : rdata = 48'b110001010000001100000000000000000000000100000000;
			// PEs: 48, 49 -> 54
			// srcs: (373, 62)(2637) -2, (1860) 0 --> (2638) -2:PENB, NI5, +, PEGB6
			10'd66 : rdata = 48'b000011101111111010100000101000000000000011100000;
			// PEs: 48 -> 
			// srcs: (375, 63)(1891) 2 --> (1891) 2:PENB, pass, 
			10'd67 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 48, 49 -> 51
			// srcs: (381, 64)(2668) -2, (1891) 2 --> (2669) 0:PENB, ALU, +, PEGB3
			10'd68 : rdata = 48'b000011101111111000111111111000000000000010110000;
			// PEs: 48 -> 
			// srcs: (383, 65)(1915) 0 --> (1915) 0:PENB, pass, 
			10'd69 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 48, 49 -> 52
			// srcs: (389, 66)(2691) -2, (1915) 0 --> (2692) -2:PENB, ALU, +, PEGB4
			10'd70 : rdata = 48'b000011101111111000111111111000000000000011000000;
			// PEs: 48 -> 
			// srcs: (391, 68)(1989) 4 --> (1989) 4:PENB, pass, 
			10'd71 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 48, 49 -> 48
			// srcs: (397, 69)(2767) 2, (1989) 4 --> (2768) 6:PENB, ALU, +, PEGB0
			10'd72 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 48 -> 
			// srcs: (399, 70)(2007) 0 --> (2007) 0:PENB, pass, 
			10'd73 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 48, 49 -> 48
			// srcs: (405, 71)(2785) 4, (2007) 0 --> (2786) 4:PENB, ALU, +, PEGB0
			10'd74 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 48 -> 
			// srcs: (407, 72)(2026) -1 --> (2026) -1:PENB, pass, 
			10'd75 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 48, 49 -> 49
			// srcs: (413, 73)(2804) 0, (2026) -1 --> (2805) -1:PENB, ALU, +, NI3
			10'd76 : rdata = 48'b000011101111111000111111111100011000000000000000;
			// PEs: 48, 49 -> 49
			// srcs: (414, 75)(2910) 0, (2133) -2 --> (2911) -2:PENB, NI1, +, NI5
			10'd77 : rdata = 48'b000011101111111010100000001100101000000000000000;
			// PEs: 48, 50 -> 50
			// srcs: (415, 76)(2912) -1, (2136) -6 --> (2913) -7:PENB, PEGB2, +, PENB
			10'd78 : rdata = 48'b000011101111111011100000100000000000000100000000;
			// PEs: 48, 51 -> 49
			// srcs: (416, 77)(2917) 0, (2139) 1 --> (2918) 1:PENB, PEGB3, +, NI1
			10'd79 : rdata = 48'b000011101111111011100000110100001000000000000000;
			// PEs: 49 -> 50
			// srcs: (422, 109)(2911) -2 --> (2911) -2:NI5, pass, PENB
			10'd80 : rdata = 48'b110001010000010100000000000000000000000100000000;
			// PEs: 48, 54 -> 48
			// srcs: (424, 78)(2924) -3, (2148) 0 --> (2925) -3:PENB, PEGB6, +, PEGB0
			10'd81 : rdata = 48'b000011101111111011100001100000000000000010000000;
			// PEs: 48 -> 
			// srcs: (533, 79)(2160) 4 --> (2160) 4:PENB, pass, 
			10'd82 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 48, 49 -> 49
			// srcs: (539, 80)(2935) -3, (2160) 4 --> (2936) 1:PENB, ALU, +, NI5
			10'd83 : rdata = 48'b000011101111111000111111111100101000000000000000;
			// PEs: 48 -> 
			// srcs: (541, 81)(2179) -3 --> (2179) -3:PENB, pass, 
			10'd84 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 48, 49 -> 48
			// srcs: (547, 82)(2957) 3, (2179) -3 --> (2958) 0:PENB, ALU, +, PEGB0
			10'd85 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 49, 48 -> 48
			// srcs: (548, 83)(2969) -4, (2191) 6 --> (2970) 2:NI0, PENB, +, PEGB0
			10'd86 : rdata = 48'b000011010000000011011111110000000000000010000000;
			// PEs: 49, 48 -> 48
			// srcs: (549, 84)(2974) 0, (2197) 0 --> (2975) 0:NI4, PENB, +, PEGB0
			10'd87 : rdata = 48'b000011010000010011011111110000000000000010000000;
			// PEs: 48 -> 
			// srcs: (551, 85)(2268) 1 --> (2268) 1:PENB, pass, 
			10'd88 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 48, 49 -> 49
			// srcs: (557, 86)(3046) 1, (2268) 1 --> (3047) 2:PENB, ALU, +, NI0
			10'd89 : rdata = 48'b000011101111111000111111111100000000000000000000;
			// PEs: 48 -> 
			// srcs: (559, 87)(2292) -2 --> (2292) -2:PENB, pass, 
			10'd90 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 48, 49 -> 48
			// srcs: (565, 88)(3069) 6, (2292) -2 --> (3070) 4:PENB, ALU, +, PEGB0
			10'd91 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 48 -> 
			// srcs: (567, 89)(2307) 2 --> (2307) 2:PENB, pass, 
			10'd92 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 48, 49 -> 48
			// srcs: (573, 90)(3082) -4, (2307) 2 --> (3083) -2:PENB, ALU, +, PEGB0
			10'd93 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 48, 54 -> 48
			// srcs: (581, 92)(3107) -6, (2332) -3 --> (3108) -9:PENB, PEGB6, +, PEGB0
			10'd94 : rdata = 48'b000011101111111011100001100000000000000010000000;
			// PEs: 48 -> 
			// srcs: (582, 93)(2366) -11 --> (2366) -11:PENB, pass, 
			10'd95 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 48, 49 -> 48
			// srcs: (587, 94)(2364) -11, (2366) -11 --> (2367) -22:PENB, ALU, +, PEGB0
			10'd96 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 48 -> 
			// srcs: (589, 95)(2414) -3 --> (2414) -3:PENB, pass, 
			10'd97 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 48, 49 -> 48
			// srcs: (595, 96)(2412) 0, (2414) -3 --> (2415) -3:PENB, ALU, +, PEGB0
			10'd98 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 48 -> 
			// srcs: (597, 97)(2469) -5 --> (2469) -5:PENB, pass, 
			10'd99 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 48, 49 -> 49
			// srcs: (603, 98)(2467) 0, (2469) -5 --> (2470) -5:PENB, ALU, +, NI4
			10'd100 : rdata = 48'b000011101111111000111111111100100000000000000000;
			// PEs: 48, 49 -> 50
			// srcs: (604, 99)(2554) -1, (2556) 1 --> (2557) 0:PENB, NI2, +, PENB
			10'd101 : rdata = 48'b000011101111111010100000010000000000000100000000;
			// PEs: 48 -> 
			// srcs: (606, 101)(2620) 1 --> (2620) 1:PENB, pass, 
			10'd102 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 48, 49 -> 48
			// srcs: (612, 102)(2618) -2, (2620) 1 --> (2621) -1:PENB, ALU, +, PEGB0
			10'd103 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 48 -> 
			// srcs: (614, 103)(2681) -5 --> (2681) -5:PENB, pass, 
			10'd104 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 48, 49 -> 48
			// srcs: (620, 104)(2679) 4, (2681) -5 --> (2682) -1:PENB, ALU, +, PEGB0
			10'd105 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 48, 49 -> 48
			// srcs: (621, 105)(2803) 3, (2805) -1 --> (2806) 2:PENB, NI3, +, PEGB0
			10'd106 : rdata = 48'b000011101111111010100000011000000000000010000000;
			// PEs: 48 -> 
			// srcs: (623, 106)(2816) -3 --> (2816) -3:PENB, pass, 
			10'd107 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 48, 49 -> 49
			// srcs: (629, 107)(2814) 9, (2816) -3 --> (2817) 6:PENB, ALU, +, NI2
			10'd108 : rdata = 48'b000011101111111000111111111100010000000000000000;
			// PEs: 48, 51 -> 49
			// srcs: (663, 108)(2886) -9, (2888) 12 --> (2889) 3:PENB, PEGB3, +, NI3
			10'd109 : rdata = 48'b000011101111111011100000110100011000000000000000;
			// PEs: 49, 48 -> 48
			// srcs: (664, 110)(2918) 1, (2920) -2 --> (2921) -1:NI1, PENB, +, PEGB0
			10'd110 : rdata = 48'b000011010000000111011111110000000000000010000000;
			// PEs: 48, 49 -> 48
			// srcs: (665, 111)(2934) 8, (2936) 1 --> (2937) 9:PENB, NI5, +, PEGB0
			10'd111 : rdata = 48'b000011101111111010100000101000000000000010000000;
			// PEs: 49, 48 -> 49
			// srcs: (677, 112)(3047) 2, (3049) -2 --> (3050) 0:NI0, PENB, +, NI1
			10'd112 : rdata = 48'b000011010000000011011111110100001000000000000000;
			// PEs: 48 -> 
			// srcs: (678, 113)(2390) 7 --> (2390) 7:PENB, pass, 
			10'd113 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 48, 49 -> 48
			// srcs: (684, 114)(2385) -3, (2390) 7 --> (2391) 4:PENB, ALU, +, PEGB0
			10'd114 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 49, 48 -> 48
			// srcs: (685, 115)(2470) -5, (2475) 12 --> (2476) 7:NI4, PENB, +, PEGB0
			10'd115 : rdata = 48'b000011010000010011011111110000000000000010000000;
			// PEs: 48 -> 
			// srcs: (743, 116)(2546) -5 --> (2546) -5:PENB, pass, 
			10'd116 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 48, 49 -> 48
			// srcs: (753, 117)(2541) -7, (2546) -5 --> (2547) -12:PENB, ALU, +, PEGB0
			10'd117 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 54, 48 -> 48
			// srcs: (754, 118)(2639) 0, (2644) 2 --> (2645) 2:PEGB6, PENB, +, PEGB0
			10'd118 : rdata = 48'b000011110000110011011111110000000000000010000000;
			// PEs: 48, 51 -> 48
			// srcs: (1386, 119)(2725) 4, (2730) 14 --> (2731) 18:PENB, PEGB3, +, PEGB0
			10'd119 : rdata = 48'b000011101111111011100000110000000000000010000000;
			// PEs: 48, 49 -> 48
			// srcs: (1387, 120)(2812) -9, (2817) 6 --> (2818) -3:PENB, NI2, +, PEGB0
			10'd120 : rdata = 48'b000011101111111010100000010000000000000010000000;
			// PEs: 48, 49 -> 49
			// srcs: (1388, 121)(2884) 2, (2889) 3 --> (2890) 5:PENB, NI3, +, NI0
			10'd121 : rdata = 48'b000011101111111010100000011100000000000000000000;
			// PEs: 48, 49 -> 48
			// srcs: (1389, 122)(3045) -9, (3050) 0 --> (3051) -9:PENB, NI1, +, PEGB0
			10'd122 : rdata = 48'b000011101111111010100000001000000000000010000000;
			// PEs: 48 -> 
			// srcs: (1390, 123)(2450) 8 --> (2450) 8:PENB, pass, 
			10'd123 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 48, 49 -> 49
			// srcs: (1395, 124)(2439) 10, (2450) 8 --> (2451) 18:PENB, ALU, +, NI1
			10'd124 : rdata = 48'b000011101111111000111111111100001000000000000000;
			// PEs: 48 -> 
			// srcs: (1397, 125)(2694) -4 --> (2694) -4:PENB, pass, 
			10'd125 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 48, 49 -> 49
			// srcs: (1403, 126)(2683) -4, (2694) -4 --> (2695) -8:PENB, ALU, +, NI2
			10'd126 : rdata = 48'b000011101111111000111111111100010000000000000000;
			// PEs: 48, 49 -> 49
			// srcs: (1404, 127)(2879) 12, (2890) 5 --> (2891) 17:PENB, NI0, +, NI3
			10'd127 : rdata = 48'b000011101111111010100000000100011000000000000000;
			// PEs: 48, 49 -> 48
			// srcs: (1405, 128)(2428) -4, (2451) 18 --> (2452) 14:PENB, NI1, +, PEGB0
			10'd128 : rdata = 48'b000011101111111010100000001000000000000010000000;
			// PEs: 48, 49 -> 48
			// srcs: (1413, 129)(2672) -6, (2695) -8 --> (2696) -14:PENB, NI2, +, PEGB0
			10'd129 : rdata = 48'b000011101111111010100000010000000000000010000000;
			// PEs: 48, 49 -> 48
			// srcs: (1414, 130)(2868) 11, (2891) 17 --> (2892) 28:PENB, NI3, +, PEGB0
			10'd130 : rdata = 48'b000011101111111010100000011000000000000010000000;
			// PEs: 48 -> 
			// srcs: (1421, 131)(2647) 48 --> (2647) 48:PENB, pass, 
			10'd131 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 48, 49 -> 48
			// srcs: (1427, 132)(2599) 4, (2647) 48 --> (2648) 52:PENB, ALU, +, PEGB0
			10'd132 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 48 -> 
			// srcs: (1465, 133)(3137) -63 --> (3137) -63:PENB, pass, 
			10'd133 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 48, 49 -> 48
			// srcs: (1475, 134)(2942) 24, (3137) -63 --> (3138) -39:PENB, ALU, +, PEGB0
			10'd134 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 48, 49 -> 50
			// srcs: (1523, 135)(3140) 47, (16) -3 --> (3153) -141:PENB, ND9, *, PENB
			10'd135 : rdata = 48'b000111101111111001100001001000000000000100000000;
			// PEs: 49, 50 -> 49
			// srcs: (1532, 149)(801) 1, (3937) -141 --> (4721) 142:NW9, PEGB2, -, NW9
			10'd136 : rdata = 48'b000100100000100111100000100000000110010000000000;
			// PEs: 48, 49 -> 50
			// srcs: (1570, 136)(3140) 47, (63) 0 --> (3200) 0:PENB, ND0, *, PENB
			10'd137 : rdata = 48'b000111101111111001100000000000000000000100000000;
			// PEs: 49, 50 -> 49
			// srcs: (1579, 150)(848) 2, (3984) 0 --> (4768) 2:NW0, PEGB2, -, NW0
			10'd138 : rdata = 48'b000100100000000011100000100000000100000000000000;
			// PEs: 48, 49 -> 50
			// srcs: (1652, 137)(3140) 47, (145) -3 --> (3282) -141:PENB, ND1, *, PENB
			10'd139 : rdata = 48'b000111101111111001100000001000000000000100000000;
			// PEs: 49, 50 -> 49
			// srcs: (1661, 151)(930) -3, (4066) -141 --> (4850) 138:NW1, PEGB2, -, NW1
			10'd140 : rdata = 48'b000100100000000111100000100000000100010000000000;
			// PEs: 48, 49 -> 50
			// srcs: (1703, 138)(3140) 47, (196) 0 --> (3333) 0:PENB, ND10, *, PENB
			10'd141 : rdata = 48'b000111101111111001100001010000000000000100000000;
			// PEs: 49, 50 -> 49
			// srcs: (1712, 152)(981) -3, (4117) 0 --> (4901) -3:NW10, PEGB2, -, NW10
			10'd142 : rdata = 48'b000100100000101011100000100000000110100000000000;
			// PEs: 48, 49 -> 50
			// srcs: (1732, 139)(3140) 47, (225) -2 --> (3362) -94:PENB, ND2, *, PENB
			10'd143 : rdata = 48'b000111101111111001100000010000000000000100000000;
			// PEs: 49, 50 -> 49
			// srcs: (1741, 153)(1010) 0, (4146) -94 --> (4930) 94:NW2, PEGB2, -, NW2
			10'd144 : rdata = 48'b000100100000001011100000100000000100100000000000;
			// PEs: 48, 49 -> 50
			// srcs: (1812, 140)(3140) 47, (305) 1 --> (3442) 47:PENB, ND3, *, PENB
			10'd145 : rdata = 48'b000111101111111001100000011000000000000100000000;
			// PEs: 49, 50 -> 49
			// srcs: (1821, 154)(1090) -2, (4226) 47 --> (5010) -49:NW3, PEGB2, -, NW3
			10'd146 : rdata = 48'b000100100000001111100000100000000100110000000000;
			// PEs: 48, 49 -> 50
			// srcs: (1887, 141)(3140) 47, (380) -2 --> (3517) -94:PENB, ND11, *, PENB
			10'd147 : rdata = 48'b000111101111111001100001011000000000000100000000;
			// PEs: 48, 49 -> 50
			// srcs: (1894, 142)(3140) 47, (387) 2 --> (3524) 94:PENB, ND4, *, PENB
			10'd148 : rdata = 48'b000111101111111001100000100000000000000100000000;
			// PEs: 49, 50 -> 49
			// srcs: (1896, 155)(1165) -3, (4301) -94 --> (5085) 91:NW11, PEGB2, -, NW11
			10'd149 : rdata = 48'b000100100000101111100000100000000110110000000000;
			// PEs: 49, 50 -> 49
			// srcs: (1903, 156)(1172) -1, (4308) 94 --> (5092) -95:NW4, PEGB2, -, NW4
			10'd150 : rdata = 48'b000100100000010011100000100000000101000000000000;
			// PEs: 48, 49 -> 50
			// srcs: (1974, 143)(3140) 47, (467) 0 --> (3604) 0:PENB, ND5, *, PENB
			10'd151 : rdata = 48'b000111101111111001100000101000000000000100000000;
			// PEs: 49, 50 -> 49
			// srcs: (1983, 157)(1252) 1, (4388) 0 --> (5172) 1:NW5, PEGB2, -, NW5
			10'd152 : rdata = 48'b000100100000010111100000100000000101010000000000;
			// PEs: 48, 49 -> 50
			// srcs: (2054, 144)(3140) 47, (547) -1 --> (3684) -47:PENB, ND6, *, PENB
			10'd153 : rdata = 48'b000111101111111001100000110000000000000100000000;
			// PEs: 49, 50 -> 49
			// srcs: (2063, 158)(1332) 2, (4468) -47 --> (5252) 49:NW6, PEGB2, -, NW6
			10'd154 : rdata = 48'b000100100000011011100000100000000101100000000000;
			// PEs: 48, 49 -> 50
			// srcs: (2071, 145)(3140) 47, (564) 2 --> (3701) 94:PENB, ND12, *, PENB
			10'd155 : rdata = 48'b000111101111111001100001100000000000000100000000;
			// PEs: 49, 50 -> 49
			// srcs: (2080, 159)(1349) -1, (4485) 94 --> (5269) -95:NW12, PEGB2, -, NW12
			10'd156 : rdata = 48'b000100100000110011100000100000000111000000000000;
			// PEs: 48, 49 -> 50
			// srcs: (2136, 146)(3140) 47, (629) 2 --> (3766) 94:PENB, ND7, *, PENB
			10'd157 : rdata = 48'b000111101111111001100000111000000000000100000000;
			// PEs: 49, 50 -> 49
			// srcs: (2145, 160)(1414) 0, (4550) 94 --> (5334) -94:NW7, PEGB2, -, NW7
			10'd158 : rdata = 48'b000100100000011111100000100000000101110000000000;
			// PEs: 48, 49 -> 50
			// srcs: (2216, 147)(3140) 47, (709) 1 --> (3846) 47:PENB, ND8, *, PENB
			10'd159 : rdata = 48'b000111101111111001100001000000000000000100000000;
			// PEs: 49, 50 -> 49
			// srcs: (2225, 161)(1494) -1, (4630) 47 --> (5414) -48:NW8, PEGB2, -, NW8
			10'd160 : rdata = 48'b000100100000100011100000100000000110000000000000;
			// PEs: 48, 49 -> 50
			// srcs: (2255, 148)(3140) 47, (748) 2 --> (3885) 94:PENB, ND13, *, PENB
			10'd161 : rdata = 48'b000111101111111001100001101000000000000100000000;
			// PEs: 49, 50 -> 49
			// srcs: (2264, 162)(1533) 0, (4669) 94 --> (5453) -94:NW13, PEGB2, -, NW13
			10'd162 : rdata = 48'b000100100000110111100000100000000111010000000000;
			default : rdata = 48'b000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 50) begin
	always @(*) begin
		case(address)
			// PEs: 50, 50 -> 48
			// srcs: (1, 0)(64) 2, (849) -3 --> (1633) -6:ND0, NW0, *, PEGB0
			10'd0 : rdata = 48'b000110110000000001000000000000000000000010000000;
			// PEs: 50, 50 -> 48
			// srcs: (2, 1)(146) -2, (931) 1 --> (1715) -2:ND1, NW1, *, PEGB0
			10'd1 : rdata = 48'b000110110000000101000000001000000000000010000000;
			// PEs: 50, 50 -> 48
			// srcs: (3, 2)(226) -2, (1011) 2 --> (1795) -4:ND2, NW2, *, PEGB0
			10'd2 : rdata = 48'b000110110000001001000000010000000000000010000000;
			// PEs: 50, 50 -> 48
			// srcs: (4, 3)(306) 0, (1091) 1 --> (1875) 0:ND3, NW3, *, PEGB0
			10'd3 : rdata = 48'b000110110000001101000000011000000000000010000000;
			// PEs: 50, 50 -> 48
			// srcs: (5, 4)(388) -2, (1173) 0 --> (1957) 0:ND4, NW4, *, PEGB0
			10'd4 : rdata = 48'b000110110000010001000000100000000000000010000000;
			// PEs: 50, 50 -> 48
			// srcs: (6, 5)(468) 1, (1253) -1 --> (2037) -1:ND5, NW5, *, PEGB0
			10'd5 : rdata = 48'b000110110000010101000000101000000000000010000000;
			// PEs: 50, 50 -> 48
			// srcs: (7, 6)(548) 1, (1333) 2 --> (2117) 2:ND6, NW6, *, PEGB0
			10'd6 : rdata = 48'b000110110000011001000000110000000000000010000000;
			// PEs: 50, 50 -> 48
			// srcs: (8, 7)(630) -2, (1415) 2 --> (2199) -4:ND7, NW7, *, PEGB0
			10'd7 : rdata = 48'b000110110000011101000000111000000000000010000000;
			// PEs: 50, 50 -> 52
			// srcs: (9, 8)(710) -2, (1495) 2 --> (2279) -4:ND8, NW8, *, PEGB4
			10'd8 : rdata = 48'b000110110000100001000001000000000000000011000000;
			// PEs: 50, 50 -> 48
			// srcs: (10, 9)(19) -1, (804) -2 --> (1588) 2:ND9, NW9, *, PEGB0
			10'd9 : rdata = 48'b000110110000100101000001001000000000000010000000;
			// PEs: 50, 50 -> 49
			// srcs: (11, 10)(199) 1, (984) -2 --> (1768) -2:ND10, NW10, *, PEGB1
			10'd10 : rdata = 48'b000110110000101001000001010000000000000010010000;
			// PEs: 50, 50 -> 50
			// srcs: (12, 11)(383) -3, (1168) 2 --> (1952) -6:ND11, NW11, *, NI0
			10'd11 : rdata = 48'b000110110000101101000001011100000000000000000000;
			// PEs: 50, 50 -> 49
			// srcs: (13, 12)(567) -3, (1352) 2 --> (2136) -6:ND12, NW12, *, PEGB1
			10'd12 : rdata = 48'b000110110000110001000001100000000000000010010000;
			// PEs: 50, 50 -> 50
			// srcs: (14, 13)(751) 2, (1536) 0 --> (2320) 0:ND13, NW13, *, NI1
			10'd13 : rdata = 48'b000110110000110101000001101100001000000000000000;
			// PEs: 48 -> 
			// srcs: (19, 14)(1703) 3 --> (1703) 3:PEGB0, pass, 
			10'd14 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 48, 50 -> 48
			// srcs: (28, 15)(1702) -4, (1703) 3 --> (2483) -1:PEGB0, ALU, +, PEGB0
			10'd15 : rdata = 48'b000011110000000000111111111000000000000010000000;
			// PEs: 48 -> 
			// srcs: (58, 16)(1865) -3 --> (1865) -3:PEGB0, pass, 
			10'd16 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 48, 50 -> 48
			// srcs: (67, 17)(1864) 1, (1865) -3 --> (2642) -2:PEGB0, ALU, +, PEGB0
			10'd17 : rdata = 48'b000011110000000000111111111000000000000010000000;
			// PEs: 49 -> 
			// srcs: (76, 20)(2726) -1 --> (2726) -1:PENB, pass, 
			10'd18 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 50, 49 -> 50
			// srcs: (83, 21)(2726) -1, (1949) 6 --> (2727) 5:ALU, PENB, +, NI2
			10'd19 : rdata = 48'b000010011111111111011111110100010000000000000000;
			// PEs: 49, 50 -> 51
			// srcs: (85, 22)(2728) 15, (1952) -6 --> (2729) 9:PENB, NI0, +, PENB
			10'd20 : rdata = 48'b000011101111111010100000000000000000000100000000;
			// PEs: 50 -> 51
			// srcs: (92, 28)(2727) 5 --> (2727) 5:NI2, pass, PENB
			10'd21 : rdata = 48'b110001010000001000000000000000000000000100000000;
			// PEs: 50 -> 48
			// srcs: (142, 25)(2320) 0 --> (2320) 0:NI1, pass, PEGB0
			10'd22 : rdata = 48'b110001010000000100000000000000000000000010000000;
			// PEs: 48 -> 
			// srcs: (221, 18)(1868) -1 --> (1868) -1:PEGB0, pass, 
			10'd23 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 48, 50 -> 51
			// srcs: (230, 19)(1867) 6, (1868) -1 --> (2649) 5:PEGB0, ALU, +, PENB
			10'd24 : rdata = 48'b000011110000000000111111111000000000000100000000;
			// PEs: 49 -> 
			// srcs: (319, 23)(2894) 5 --> (2894) 5:PENB, pass, 
			10'd25 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 49, 50 -> 48
			// srcs: (326, 24)(2893) 8, (2894) 5 --> (2895) 13:PENB, ALU, +, PEGB0
			10'd26 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 49 -> 
			// srcs: (367, 26)(2561) -2 --> (2561) -2:PENB, pass, 
			10'd27 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 49, 50 -> 50
			// srcs: (374, 27)(2559) 5, (2561) -2 --> (2562) 3:PENB, ALU, +, NI0
			10'd28 : rdata = 48'b000011101111111000111111111100000000000000000000;
			// PEs: 49 -> 
			// srcs: (417, 29)(2913) -7 --> (2913) -7:PENB, pass, 
			10'd29 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 49, 50 -> 48
			// srcs: (424, 30)(2911) -2, (2913) -7 --> (2914) -9:PENB, ALU, +, PEGB0
			10'd30 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 49, 50 -> 48
			// srcs: (607, 31)(2557) 0, (2562) 3 --> (2563) 3:PENB, NI0, +, PEGB0
			10'd31 : rdata = 48'b000011101111111010100000000000000000000010000000;
			// PEs: 50, 49 -> 49
			// srcs: (1526, 46)(3) 1, (3153) -141 --> (3937) -141:NM0, PENB, *, PEGB1
			10'd32 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 48, 50 -> 
			// srcs: (1529, 32)(3140) 47, (19) -1 --> (3156) -47:PEGB0, ND9, *, 
			10'd33 : rdata = 48'b000111110000000001100001001000000000000000000000;
			// PEs: 50, 50 -> 
			// srcs: (1532, 47)(3) 1, (3156) -47 --> (3940) -47:NM0, ALU, *, 
			10'd34 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 50, 50 -> 50
			// srcs: (1535, 64)(804) -2, (3940) -47 --> (4724) 45:NW9, ALU, -, NW9
			10'd35 : rdata = 48'b000100100000100100111111111000000110010000000000;
			// PEs: 50, 49 -> 49
			// srcs: (1573, 48)(3) 1, (3200) 0 --> (3984) 0:NM0, PENB, *, PEGB1
			10'd36 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 48, 50 -> 51
			// srcs: (1574, 33)(3140) 47, (64) 2 --> (3201) 94:PEGB0, ND0, *, PENB
			10'd37 : rdata = 48'b000111110000000001100000000000000000000100000000;
			// PEs: 50, 51 -> 50
			// srcs: (1583, 65)(849) -3, (3985) 94 --> (4769) -97:NW0, PEGB3, -, NW0
			10'd38 : rdata = 48'b000100100000000011100000110000000100000000000000;
			// PEs: 50, 49 -> 49
			// srcs: (1655, 49)(3) 1, (3282) -141 --> (4066) -141:NM0, PENB, *, PEGB1
			10'd39 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 48, 50 -> 51
			// srcs: (1656, 34)(3140) 47, (146) -2 --> (3283) -94:PEGB0, ND1, *, PENB
			10'd40 : rdata = 48'b000111110000000001100000001000000000000100000000;
			// PEs: 50, 51 -> 50
			// srcs: (1665, 66)(931) 1, (4067) -94 --> (4851) 95:NW1, PEGB3, -, NW1
			10'd41 : rdata = 48'b000100100000000111100000110000000100010000000000;
			// PEs: 50, 49 -> 49
			// srcs: (1706, 50)(3) 1, (3333) 0 --> (4117) 0:NM0, PENB, *, PEGB1
			10'd42 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 48, 50 -> 51
			// srcs: (1709, 35)(3140) 47, (199) 1 --> (3336) 47:PEGB0, ND10, *, PENB
			10'd43 : rdata = 48'b000111110000000001100001010000000000000100000000;
			// PEs: 50, 51 -> 50
			// srcs: (1718, 67)(984) -2, (4120) 47 --> (4904) -49:NW10, PEGB3, -, NW10
			10'd44 : rdata = 48'b000100100000101011100000110000000110100000000000;
			// PEs: 50, 49 -> 49
			// srcs: (1735, 51)(3) 1, (3362) -94 --> (4146) -94:NM0, PENB, *, PEGB1
			10'd45 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 48, 50 -> 51
			// srcs: (1736, 36)(3140) 47, (226) -2 --> (3363) -94:PEGB0, ND2, *, PENB
			10'd46 : rdata = 48'b000111110000000001100000010000000000000100000000;
			// PEs: 50, 51 -> 50
			// srcs: (1745, 68)(1011) 2, (4147) -94 --> (4931) 96:NW2, PEGB3, -, NW2
			10'd47 : rdata = 48'b000100100000001011100000110000000100100000000000;
			// PEs: 50, 49 -> 49
			// srcs: (1815, 52)(3) 1, (3442) 47 --> (4226) 47:NM0, PENB, *, PEGB1
			10'd48 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 48, 50 -> 51
			// srcs: (1816, 37)(3140) 47, (306) 0 --> (3443) 0:PEGB0, ND3, *, PENB
			10'd49 : rdata = 48'b000111110000000001100000011000000000000100000000;
			// PEs: 50, 51 -> 50
			// srcs: (1825, 69)(1091) 1, (4227) 0 --> (5011) 1:NW3, PEGB3, -, NW3
			10'd50 : rdata = 48'b000100100000001111100000110000000100110000000000;
			// PEs: 50, 49 -> 49
			// srcs: (1890, 53)(3) 1, (3517) -94 --> (4301) -94:NM0, PENB, *, PEGB1
			10'd51 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 48, 50 -> 
			// srcs: (1893, 38)(3140) 47, (383) -3 --> (3520) -141:PEGB0, ND11, *, 
			10'd52 : rdata = 48'b000111110000000001100001011000000000000000000000;
			// PEs: 50, 50 -> 50
			// srcs: (1896, 54)(3) 1, (3520) -141 --> (4304) -141:NM0, ALU, *, NI0
			10'd53 : rdata = 48'b000111000000000000111111111100000000000000000000;
			// PEs: 50, 49 -> 49
			// srcs: (1897, 55)(3) 1, (3524) 94 --> (4308) 94:NM0, PENB, *, PEGB1
			10'd54 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 48, 50 -> 51
			// srcs: (1898, 39)(3140) 47, (388) -2 --> (3525) -94:PEGB0, ND4, *, PENB
			10'd55 : rdata = 48'b000111110000000001100000100000000000000100000000;
			// PEs: 50, 50 -> 50
			// srcs: (1899, 70)(1168) 2, (4304) -141 --> (5088) 143:NW11, NI0, -, NW11
			10'd56 : rdata = 48'b000100100000101110100000000000000110110000000000;
			// PEs: 50, 51 -> 50
			// srcs: (1907, 71)(1173) 0, (4309) -94 --> (5093) 94:NW4, PEGB3, -, NW4
			10'd57 : rdata = 48'b000100100000010011100000110000000101000000000000;
			// PEs: 50, 49 -> 49
			// srcs: (1977, 56)(3) 1, (3604) 0 --> (4388) 0:NM0, PENB, *, PEGB1
			10'd58 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 48, 50 -> 51
			// srcs: (1978, 40)(3140) 47, (468) 1 --> (3605) 47:PEGB0, ND5, *, PENB
			10'd59 : rdata = 48'b000111110000000001100000101000000000000100000000;
			// PEs: 50, 51 -> 50
			// srcs: (1987, 72)(1253) -1, (4389) 47 --> (5173) -48:NW5, PEGB3, -, NW5
			10'd60 : rdata = 48'b000100100000010111100000110000000101010000000000;
			// PEs: 50, 49 -> 49
			// srcs: (2057, 57)(3) 1, (3684) -47 --> (4468) -47:NM0, PENB, *, PEGB1
			10'd61 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 48, 50 -> 51
			// srcs: (2058, 41)(3140) 47, (548) 1 --> (3685) 47:PEGB0, ND6, *, PENB
			10'd62 : rdata = 48'b000111110000000001100000110000000000000100000000;
			// PEs: 50, 51 -> 50
			// srcs: (2067, 73)(1333) 2, (4469) 47 --> (5253) -45:NW6, PEGB3, -, NW6
			10'd63 : rdata = 48'b000100100000011011100000110000000101100000000000;
			// PEs: 50, 49 -> 49
			// srcs: (2074, 58)(3) 1, (3701) 94 --> (4485) 94:NM0, PENB, *, PEGB1
			10'd64 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 48, 50 -> 
			// srcs: (2077, 42)(3140) 47, (567) -3 --> (3704) -141:PEGB0, ND12, *, 
			10'd65 : rdata = 48'b000111110000000001100001100000000000000000000000;
			// PEs: 50, 50 -> 
			// srcs: (2080, 59)(3) 1, (3704) -141 --> (4488) -141:NM0, ALU, *, 
			10'd66 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 50, 50 -> 50
			// srcs: (2083, 74)(1352) 2, (4488) -141 --> (5272) 143:NW12, ALU, -, NW12
			10'd67 : rdata = 48'b000100100000110000111111111000000111000000000000;
			// PEs: 50, 49 -> 49
			// srcs: (2139, 60)(3) 1, (3766) 94 --> (4550) 94:NM0, PENB, *, PEGB1
			10'd68 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 48, 50 -> 51
			// srcs: (2140, 43)(3140) 47, (630) -2 --> (3767) -94:PEGB0, ND7, *, PENB
			10'd69 : rdata = 48'b000111110000000001100000111000000000000100000000;
			// PEs: 50, 51 -> 50
			// srcs: (2149, 75)(1415) 2, (4551) -94 --> (5335) 96:NW7, PEGB3, -, NW7
			10'd70 : rdata = 48'b000100100000011111100000110000000101110000000000;
			// PEs: 50, 49 -> 49
			// srcs: (2219, 61)(3) 1, (3846) 47 --> (4630) 47:NM0, PENB, *, PEGB1
			10'd71 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 48, 50 -> 51
			// srcs: (2220, 44)(3140) 47, (710) -2 --> (3847) -94:PEGB0, ND8, *, PENB
			10'd72 : rdata = 48'b000111110000000001100001000000000000000100000000;
			// PEs: 50, 51 -> 50
			// srcs: (2229, 76)(1495) 2, (4631) -94 --> (5415) 96:NW8, PEGB3, -, NW8
			10'd73 : rdata = 48'b000100100000100011100000110000000110000000000000;
			// PEs: 50, 49 -> 49
			// srcs: (2258, 62)(3) 1, (3885) 94 --> (4669) 94:NM0, PENB, *, PEGB1
			10'd74 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 48, 50 -> 
			// srcs: (2261, 45)(3140) 47, (751) 2 --> (3888) 94:PEGB0, ND13, *, 
			10'd75 : rdata = 48'b000111110000000001100001101000000000000000000000;
			// PEs: 50, 50 -> 
			// srcs: (2264, 63)(3) 1, (3888) 94 --> (4672) 94:NM0, ALU, *, 
			10'd76 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 50, 50 -> 50
			// srcs: (2267, 77)(1536) 0, (4672) 94 --> (5456) -94:NW13, ALU, -, NW13
			10'd77 : rdata = 48'b000100100000110100111111111000000111010000000000;
			default : rdata = 48'b000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 51) begin
	always @(*) begin
		case(address)
			// PEs: 51, 51 -> 48
			// srcs: (1, 0)(66) 1, (851) -1 --> (1635) -1:ND0, NW0, *, PEGB0
			10'd0 : rdata = 48'b000110110000000001000000000000000000000010000000;
			// PEs: 51, 51 -> 48
			// srcs: (2, 1)(148) -3, (933) 0 --> (1717) 0:ND1, NW1, *, PEGB0
			10'd1 : rdata = 48'b000110110000000101000000001000000000000010000000;
			// PEs: 51, 51 -> 48
			// srcs: (3, 2)(228) 2, (1013) -2 --> (1797) -4:ND2, NW2, *, PEGB0
			10'd2 : rdata = 48'b000110110000001001000000010000000000000010000000;
			// PEs: 51, 51 -> 48
			// srcs: (4, 3)(308) 0, (1093) 0 --> (1877) 0:ND3, NW3, *, PEGB0
			10'd3 : rdata = 48'b000110110000001101000000011000000000000010000000;
			// PEs: 51, 51 -> 48
			// srcs: (5, 4)(390) 0, (1175) 2 --> (1959) 0:ND4, NW4, *, PEGB0
			10'd4 : rdata = 48'b000110110000010001000000100000000000000010000000;
			// PEs: 51, 51 -> 48
			// srcs: (6, 5)(470) -3, (1255) -1 --> (2039) 3:ND5, NW5, *, PEGB0
			10'd5 : rdata = 48'b000110110000010101000000101000000000000010000000;
			// PEs: 51, 51 -> 48
			// srcs: (7, 6)(550) -2, (1335) -2 --> (2119) 4:ND6, NW6, *, PEGB0
			10'd6 : rdata = 48'b000110110000011001000000110000000000000010000000;
			// PEs: 51, 51 -> 48
			// srcs: (8, 7)(632) -1, (1417) -2 --> (2201) 2:ND7, NW7, *, PEGB0
			10'd7 : rdata = 48'b000110110000011101000000111000000000000010000000;
			// PEs: 51, 51 -> 53
			// srcs: (9, 8)(712) 2, (1497) -3 --> (2281) -6:ND8, NW8, *, PEGB5
			10'd8 : rdata = 48'b000110110000100001000001000000000000000011010000;
			// PEs: 51, 51 -> 49
			// srcs: (10, 9)(22) -2, (807) -1 --> (1591) 2:ND9, NW9, *, PEGB1
			10'd9 : rdata = 48'b000110110000100101000001001000000000000010010000;
			// PEs: 51, 51 -> 49
			// srcs: (11, 10)(206) -3, (991) 0 --> (1775) 0:ND10, NW10, *, PEGB1
			10'd10 : rdata = 48'b000110110000101001000001010000000000000010010000;
			// PEs: 51, 51 -> 53
			// srcs: (12, 11)(386) 0, (1171) 0 --> (1955) 0:ND11, NW11, *, PEGB5
			10'd11 : rdata = 48'b000110110000101101000001011000000000000011010000;
			// PEs: 51, 51 -> 49
			// srcs: (13, 12)(570) -1, (1355) -1 --> (2139) 1:ND12, NW12, *, PEGB1
			10'd12 : rdata = 48'b000110110000110001000001100000000000000010010000;
			// PEs: 51, 51 -> 51
			// srcs: (14, 13)(754) -2, (1539) -1 --> (2323) 2:ND13, NW13, *, NI0
			10'd13 : rdata = 48'b000110110000110101000001101100000000000000000000;
			// PEs: 48 -> 
			// srcs: (21, 14)(1706) 2 --> (1706) 2:PEGB0, pass, 
			10'd14 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 48, 51 -> 48
			// srcs: (30, 15)(1705) 6, (1706) 2 --> (2485) 8:PEGB0, ALU, +, PEGB0
			10'd15 : rdata = 48'b000011110000000000111111111000000000000010000000;
			// PEs: 48 -> 
			// srcs: (60, 16)(1872) 3 --> (1872) 3:PEGB0, pass, 
			10'd16 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 48, 51 -> 48
			// srcs: (69, 17)(1871) 0, (1872) 3 --> (2652) 3:PEGB0, ALU, +, PEGB0
			10'd17 : rdata = 48'b000011110000000000111111111000000000000010000000;
			// PEs: 50 -> 
			// srcs: (87, 26)(2729) 9 --> (2729) 9:PENB, pass, 
			10'd18 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 50, 51 -> 51
			// srcs: (94, 27)(2727) 5, (2729) 9 --> (2730) 14:PENB, ALU, +, NI1
			10'd19 : rdata = 48'b000011101111111000111111111100001000000000000000;
			// PEs: 51 -> 48
			// srcs: (157, 23)(2323) 2 --> (2323) 2:NI0, pass, PEGB0
			10'd20 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 48 -> 
			// srcs: (256, 18)(1870) 0 --> (1870) 0:PEGB0, pass, 
			10'd21 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 48, 51 -> 
			// srcs: (265, 19)(1869) 0, (1870) 0 --> (2650) 0:PEGB0, ALU, +, 
			10'd22 : rdata = 48'b000011110000000000111111111000000000000000000000;
			// PEs: 50, 51 -> 48
			// srcs: (268, 20)(2649) 5, (2650) 0 --> (2651) 5:PENB, ALU, +, PEGB0
			10'd23 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 48 -> 
			// srcs: (445, 21)(2111) 0 --> (2111) 0:PEGB0, pass, 
			10'd24 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 49, 51 -> 49
			// srcs: (447, 22)(2887) 12, (2111) 0 --> (2888) 12:PEGB1, ALU, +, PEGB1
			10'd25 : rdata = 48'b000011110000001000111111111000000000000010010000;
			// PEs: 48 -> 
			// srcs: (594, 24)(2667) -10 --> (2667) -10:PEGB0, pass, 
			10'd26 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 51, 49 -> 48
			// srcs: (596, 25)(2667) -10, (2669) 0 --> (2670) -10:ALU, PEGB1, +, PEGB0
			10'd27 : rdata = 48'b000010011111111111100000010000000000000010000000;
			// PEs: 51 -> 49
			// srcs: (1381, 28)(2730) 14 --> (2730) 14:NI1, pass, PEGB1
			10'd28 : rdata = 48'b110001010000000100000000000000000000000010010000;
			// PEs: 48, 51 -> 
			// srcs: (1532, 29)(3140) 47, (22) -2 --> (3159) -94:PEGB0, ND9, *, 
			10'd29 : rdata = 48'b000111110000000001100001001000000000000000000000;
			// PEs: 51, 51 -> 
			// srcs: (1535, 43)(3) 1, (3159) -94 --> (3943) -94:NM0, ALU, *, 
			10'd30 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 51, 51 -> 51
			// srcs: (1538, 58)(807) -1, (3943) -94 --> (4727) 93:NW9, ALU, -, NW9
			10'd31 : rdata = 48'b000100100000100100111111111000000110010000000000;
			// PEs: 48, 51 -> 52
			// srcs: (1576, 30)(3140) 47, (66) 1 --> (3203) 47:PEGB0, ND0, *, PENB
			10'd32 : rdata = 48'b000111110000000001100000000000000000000100000000;
			// PEs: 51, 50 -> 50
			// srcs: (1577, 44)(3) 1, (3201) 94 --> (3985) 94:NM0, PENB, *, PEGB2
			10'd33 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 51, 52 -> 51
			// srcs: (1585, 59)(851) -1, (3987) 47 --> (4771) -48:NW0, PEGB4, -, NW0
			10'd34 : rdata = 48'b000100100000000011100001000000000100000000000000;
			// PEs: 48, 51 -> 52
			// srcs: (1658, 31)(3140) 47, (148) -3 --> (3285) -141:PEGB0, ND1, *, PENB
			10'd35 : rdata = 48'b000111110000000001100000001000000000000100000000;
			// PEs: 51, 50 -> 50
			// srcs: (1659, 45)(3) 1, (3283) -94 --> (4067) -94:NM0, PENB, *, PEGB2
			10'd36 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 51, 52 -> 51
			// srcs: (1667, 60)(933) 0, (4069) -141 --> (4853) 141:NW1, PEGB4, -, NW1
			10'd37 : rdata = 48'b000100100000000111100001000000000100010000000000;
			// PEs: 51, 50 -> 50
			// srcs: (1712, 46)(3) 1, (3336) 47 --> (4120) 47:NM0, PENB, *, PEGB2
			10'd38 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 48, 51 -> 
			// srcs: (1716, 32)(3140) 47, (206) -3 --> (3343) -141:PEGB0, ND10, *, 
			10'd39 : rdata = 48'b000111110000000001100001010000000000000000000000;
			// PEs: 51, 51 -> 
			// srcs: (1719, 47)(3) 1, (3343) -141 --> (4127) -141:NM0, ALU, *, 
			10'd40 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 51, 51 -> 51
			// srcs: (1722, 61)(991) 0, (4127) -141 --> (4911) 141:NW10, ALU, -, NW10
			10'd41 : rdata = 48'b000100100000101000111111111000000110100000000000;
			// PEs: 48, 51 -> 52
			// srcs: (1738, 33)(3140) 47, (228) 2 --> (3365) 94:PEGB0, ND2, *, PENB
			10'd42 : rdata = 48'b000111110000000001100000010000000000000100000000;
			// PEs: 51, 50 -> 50
			// srcs: (1739, 48)(3) 1, (3363) -94 --> (4147) -94:NM0, PENB, *, PEGB2
			10'd43 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 51, 52 -> 51
			// srcs: (1747, 62)(1013) -2, (4149) 94 --> (4933) -96:NW2, PEGB4, -, NW2
			10'd44 : rdata = 48'b000100100000001011100001000000000100100000000000;
			// PEs: 48, 51 -> 52
			// srcs: (1818, 34)(3140) 47, (308) 0 --> (3445) 0:PEGB0, ND3, *, PENB
			10'd45 : rdata = 48'b000111110000000001100000011000000000000100000000;
			// PEs: 51, 50 -> 50
			// srcs: (1819, 49)(3) 1, (3443) 0 --> (4227) 0:NM0, PENB, *, PEGB2
			10'd46 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 51, 52 -> 51
			// srcs: (1827, 63)(1093) 0, (4229) 0 --> (5013) 0:NW3, PEGB4, -, NW3
			10'd47 : rdata = 48'b000100100000001111100001000000000100110000000000;
			// PEs: 48, 51 -> 
			// srcs: (1896, 35)(3140) 47, (386) 0 --> (3523) 0:PEGB0, ND11, *, 
			10'd48 : rdata = 48'b000111110000000001100001011000000000000000000000;
			// PEs: 51, 51 -> 51
			// srcs: (1899, 50)(3) 1, (3523) 0 --> (4307) 0:NM0, ALU, *, NI0
			10'd49 : rdata = 48'b000111000000000000111111111100000000000000000000;
			// PEs: 48, 51 -> 52
			// srcs: (1900, 36)(3140) 47, (390) 0 --> (3527) 0:PEGB0, ND4, *, PENB
			10'd50 : rdata = 48'b000111110000000001100000100000000000000100000000;
			// PEs: 51, 50 -> 50
			// srcs: (1901, 51)(3) 1, (3525) -94 --> (4309) -94:NM0, PENB, *, PEGB2
			10'd51 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 51, 51 -> 51
			// srcs: (1902, 64)(1171) 0, (4307) 0 --> (5091) 0:NW11, NI0, -, NW11
			10'd52 : rdata = 48'b000100100000101110100000000000000110110000000000;
			// PEs: 51, 52 -> 51
			// srcs: (1909, 65)(1175) 2, (4311) 0 --> (5095) 2:NW4, PEGB4, -, NW4
			10'd53 : rdata = 48'b000100100000010011100001000000000101000000000000;
			// PEs: 48, 51 -> 52
			// srcs: (1980, 37)(3140) 47, (470) -3 --> (3607) -141:PEGB0, ND5, *, PENB
			10'd54 : rdata = 48'b000111110000000001100000101000000000000100000000;
			// PEs: 51, 50 -> 50
			// srcs: (1981, 52)(3) 1, (3605) 47 --> (4389) 47:NM0, PENB, *, PEGB2
			10'd55 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 51, 52 -> 51
			// srcs: (1989, 66)(1255) -1, (4391) -141 --> (5175) 140:NW5, PEGB4, -, NW5
			10'd56 : rdata = 48'b000100100000010111100001000000000101010000000000;
			// PEs: 48, 51 -> 52
			// srcs: (2060, 38)(3140) 47, (550) -2 --> (3687) -94:PEGB0, ND6, *, PENB
			10'd57 : rdata = 48'b000111110000000001100000110000000000000100000000;
			// PEs: 51, 50 -> 50
			// srcs: (2061, 53)(3) 1, (3685) 47 --> (4469) 47:NM0, PENB, *, PEGB2
			10'd58 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 51, 52 -> 51
			// srcs: (2069, 67)(1335) -2, (4471) -94 --> (5255) 92:NW6, PEGB4, -, NW6
			10'd59 : rdata = 48'b000100100000011011100001000000000101100000000000;
			// PEs: 48, 51 -> 
			// srcs: (2080, 39)(3140) 47, (570) -1 --> (3707) -47:PEGB0, ND12, *, 
			10'd60 : rdata = 48'b000111110000000001100001100000000000000000000000;
			// PEs: 51, 51 -> 
			// srcs: (2083, 54)(3) 1, (3707) -47 --> (4491) -47:NM0, ALU, *, 
			10'd61 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 51, 51 -> 51
			// srcs: (2086, 68)(1355) -1, (4491) -47 --> (5275) 46:NW12, ALU, -, NW12
			10'd62 : rdata = 48'b000100100000110000111111111000000111000000000000;
			// PEs: 48, 51 -> 52
			// srcs: (2142, 40)(3140) 47, (632) -1 --> (3769) -47:PEGB0, ND7, *, PENB
			10'd63 : rdata = 48'b000111110000000001100000111000000000000100000000;
			// PEs: 51, 50 -> 50
			// srcs: (2143, 55)(3) 1, (3767) -94 --> (4551) -94:NM0, PENB, *, PEGB2
			10'd64 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 51, 52 -> 51
			// srcs: (2151, 69)(1417) -2, (4553) -47 --> (5337) 45:NW7, PEGB4, -, NW7
			10'd65 : rdata = 48'b000100100000011111100001000000000101110000000000;
			// PEs: 48, 51 -> 52
			// srcs: (2222, 41)(3140) 47, (712) 2 --> (3849) 94:PEGB0, ND8, *, PENB
			10'd66 : rdata = 48'b000111110000000001100001000000000000000100000000;
			// PEs: 51, 50 -> 50
			// srcs: (2223, 56)(3) 1, (3847) -94 --> (4631) -94:NM0, PENB, *, PEGB2
			10'd67 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 51, 52 -> 51
			// srcs: (2231, 70)(1497) -3, (4633) 94 --> (5417) -97:NW8, PEGB4, -, NW8
			10'd68 : rdata = 48'b000100100000100011100001000000000110000000000000;
			// PEs: 48, 51 -> 
			// srcs: (2264, 42)(3140) 47, (754) -2 --> (3891) -94:PEGB0, ND13, *, 
			10'd69 : rdata = 48'b000111110000000001100001101000000000000000000000;
			// PEs: 51, 51 -> 
			// srcs: (2267, 57)(3) 1, (3891) -94 --> (4675) -94:NM0, ALU, *, 
			10'd70 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 51, 51 -> 51
			// srcs: (2270, 71)(1539) -1, (4675) -94 --> (5459) 93:NW13, ALU, -, NW13
			10'd71 : rdata = 48'b000100100000110100111111111000000111010000000000;
			default : rdata = 48'b000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 52) begin
	always @(*) begin
		case(address)
			// PEs: 52, 52 -> 48
			// srcs: (1, 0)(67) 1, (852) 0 --> (1636) 0:ND0, NW0, *, PEGB0
			10'd0 : rdata = 48'b000110110000000001000000000000000000000010000000;
			// PEs: 52, 52 -> 48
			// srcs: (2, 1)(149) 2, (934) 1 --> (1718) 2:ND1, NW1, *, PEGB0
			10'd1 : rdata = 48'b000110110000000101000000001000000000000010000000;
			// PEs: 52, 52 -> 48
			// srcs: (3, 2)(229) 1, (1014) -3 --> (1798) -3:ND2, NW2, *, PEGB0
			10'd2 : rdata = 48'b000110110000001001000000010000000000000010000000;
			// PEs: 52, 52 -> 48
			// srcs: (4, 3)(309) 1, (1094) -2 --> (1878) -2:ND3, NW3, *, PEGB0
			10'd3 : rdata = 48'b000110110000001101000000011000000000000010000000;
			// PEs: 52, 52 -> 48
			// srcs: (5, 4)(391) -3, (1176) 0 --> (1960) 0:ND4, NW4, *, PEGB0
			10'd4 : rdata = 48'b000110110000010001000000100000000000000010000000;
			// PEs: 52, 52 -> 48
			// srcs: (6, 5)(471) -2, (1256) 0 --> (2040) 0:ND5, NW5, *, PEGB0
			10'd5 : rdata = 48'b000110110000010101000000101000000000000010000000;
			// PEs: 52, 52 -> 48
			// srcs: (7, 6)(551) -3, (1336) -3 --> (2120) 9:ND6, NW6, *, PEGB0
			10'd6 : rdata = 48'b000110110000011001000000110000000000000010000000;
			// PEs: 52, 52 -> 48
			// srcs: (8, 7)(633) -2, (1418) -1 --> (2202) 2:ND7, NW7, *, PEGB0
			10'd7 : rdata = 48'b000110110000011101000000111000000000000010000000;
			// PEs: 52, 52 -> 53
			// srcs: (9, 8)(713) -2, (1498) -1 --> (2282) 2:ND8, NW8, *, PENB
			10'd8 : rdata = 48'b000110110000100001000001000000000000000100000000;
			// PEs: 52, 52 -> 48
			// srcs: (10, 9)(25) 1, (810) -1 --> (1594) -1:ND9, NW9, *, PEGB0
			10'd9 : rdata = 48'b000110110000100101000001001000000000000010000000;
			// PEs: 52, 52 -> 49
			// srcs: (11, 10)(209) -3, (994) 2 --> (1778) -6:ND10, NW10, *, PEGB1
			10'd10 : rdata = 48'b000110110000101001000001010000000000000010010000;
			// PEs: 52, 52 -> 52
			// srcs: (12, 11)(389) -2, (1174) -2 --> (1958) 4:ND11, NW11, *, NI0
			10'd11 : rdata = 48'b000110110000101101000001011100000000000000000000;
			// PEs: 52, 52 -> 52
			// srcs: (13, 12)(573) 1, (1358) -2 --> (2142) -2:ND12, NW12, *, NI1
			10'd12 : rdata = 48'b000110110000110001000001100100001000000000000000;
			// PEs: 52, 52 -> 52
			// srcs: (14, 13)(757) -2, (1542) 1 --> (2326) -2:ND13, NW13, *, NI2
			10'd13 : rdata = 48'b000110110000110101000001101100010000000000000000;
			// PEs: 50 -> 
			// srcs: (15, 16)(2279) -4 --> (2279) -4:PEGB2, pass, 
			10'd14 : rdata = 48'b110001110000010000000000000000000000000000000000;
			// PEs: 49, 52 -> 52
			// srcs: (17, 17)(2278) -1, (2279) -4 --> (3057) -5:PEGB1, ALU, +, NI3
			10'd15 : rdata = 48'b000011110000001000111111111100011000000000000000;
			// PEs: 48 -> 
			// srcs: (27, 14)(1709) 0 --> (1709) 0:PEGB0, pass, 
			10'd16 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 48, 52 -> 48
			// srcs: (36, 15)(1708) 0, (1709) 0 --> (2489) 0:PEGB0, ALU, +, PEGB0
			10'd17 : rdata = 48'b000011110000000000111111111000000000000010000000;
			// PEs: 52 -> 48
			// srcs: (137, 20)(1958) 4 --> (1958) 4:NI0, pass, PEGB0
			10'd18 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 52 -> 48
			// srcs: (142, 21)(2142) -2 --> (2142) -2:NI1, pass, PEGB0
			10'd19 : rdata = 48'b110001010000000100000000000000000000000010000000;
			// PEs: 52 -> 48
			// srcs: (161, 22)(3057) -5 --> (3057) -5:NI3, pass, PEGB0
			10'd20 : rdata = 48'b110001010000001100000000000000000000000010000000;
			// PEs: 52 -> 48
			// srcs: (177, 23)(2326) -2 --> (2326) -2:NI2, pass, PEGB0
			10'd21 : rdata = 48'b110001010000001000000000000000000000000010000000;
			// PEs: 48 -> 
			// srcs: (372, 18)(1879) 4 --> (1879) 4:PEGB0, pass, 
			10'd22 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 48, 52 -> 48
			// srcs: (381, 19)(2657) -2, (1879) 4 --> (2658) 2:PEGB0, ALU, +, PEGB0
			10'd23 : rdata = 48'b000011110000000000111111111000000000000010000000;
			// PEs: 48 -> 
			// srcs: (595, 24)(2690) 1 --> (2690) 1:PEGB0, pass, 
			10'd24 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 52, 49 -> 48
			// srcs: (597, 25)(2690) 1, (2692) -2 --> (2693) -1:ALU, PEGB1, +, PEGB0
			10'd25 : rdata = 48'b000010011111111111100000010000000000000010000000;
			// PEs: 48, 52 -> 
			// srcs: (1535, 26)(3140) 47, (25) 1 --> (3162) 47:PEGB0, ND9, *, 
			10'd26 : rdata = 48'b000111110000000001100001001000000000000000000000;
			// PEs: 52, 52 -> 
			// srcs: (1538, 40)(3) 1, (3162) 47 --> (3946) 47:NM0, ALU, *, 
			10'd27 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 52, 52 -> 52
			// srcs: (1541, 56)(810) -1, (3946) 47 --> (4730) -48:NW9, ALU, -, NW9
			10'd28 : rdata = 48'b000100100000100100111111111000000110010000000000;
			// PEs: 48, 52 -> 53
			// srcs: (1577, 27)(3140) 47, (67) 1 --> (3204) 47:PEGB0, ND0, *, PENB
			10'd29 : rdata = 48'b000111110000000001100000000000000000000100000000;
			// PEs: 52, 51 -> 51
			// srcs: (1579, 41)(3) 1, (3203) 47 --> (3987) 47:NM0, PENB, *, PEGB3
			10'd30 : rdata = 48'b000111000000000011011111110000000000000010110000;
			// PEs: 52, 53 -> 52
			// srcs: (1586, 57)(852) 0, (3988) 47 --> (4772) -47:NW0, PEGB5, -, NW0
			10'd31 : rdata = 48'b000100100000000011100001010000000100000000000000;
			// PEs: 48, 52 -> 53
			// srcs: (1659, 28)(3140) 47, (149) 2 --> (3286) 94:PEGB0, ND1, *, PENB
			10'd32 : rdata = 48'b000111110000000001100000001000000000000100000000;
			// PEs: 52, 51 -> 51
			// srcs: (1661, 42)(3) 1, (3285) -141 --> (4069) -141:NM0, PENB, *, PEGB3
			10'd33 : rdata = 48'b000111000000000011011111110000000000000010110000;
			// PEs: 52, 53 -> 52
			// srcs: (1668, 58)(934) 1, (4070) 94 --> (4854) -93:NW1, PEGB5, -, NW1
			10'd34 : rdata = 48'b000100100000000111100001010000000100010000000000;
			// PEs: 48, 52 -> 
			// srcs: (1719, 29)(3140) 47, (209) -3 --> (3346) -141:PEGB0, ND10, *, 
			10'd35 : rdata = 48'b000111110000000001100001010000000000000000000000;
			// PEs: 52, 52 -> 
			// srcs: (1722, 43)(3) 1, (3346) -141 --> (4130) -141:NM0, ALU, *, 
			10'd36 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 52, 52 -> 52
			// srcs: (1725, 59)(994) 2, (4130) -141 --> (4914) 143:NW10, ALU, -, NW10
			10'd37 : rdata = 48'b000100100000101000111111111000000110100000000000;
			// PEs: 48, 52 -> 53
			// srcs: (1739, 30)(3140) 47, (229) 1 --> (3366) 47:PEGB0, ND2, *, PENB
			10'd38 : rdata = 48'b000111110000000001100000010000000000000100000000;
			// PEs: 52, 51 -> 51
			// srcs: (1741, 44)(3) 1, (3365) 94 --> (4149) 94:NM0, PENB, *, PEGB3
			10'd39 : rdata = 48'b000111000000000011011111110000000000000010110000;
			// PEs: 52, 53 -> 52
			// srcs: (1748, 60)(1014) -3, (4150) 47 --> (4934) -50:NW2, PEGB5, -, NW2
			10'd40 : rdata = 48'b000100100000001011100001010000000100100000000000;
			// PEs: 48, 52 -> 52
			// srcs: (1819, 31)(3140) 47, (309) 1 --> (3446) 47:PEGB0, ND3, *, NI0
			10'd41 : rdata = 48'b000111110000000001100000011100000000000000000000;
			// PEs: 52, 51 -> 51
			// srcs: (1821, 45)(3) 1, (3445) 0 --> (4229) 0:NM0, PENB, *, PEGB3
			10'd42 : rdata = 48'b000111000000000011011111110000000000000010110000;
			// PEs: 52, 52 -> 
			// srcs: (1822, 46)(3) 1, (3446) 47 --> (4230) 47:NM0, NI0, *, 
			10'd43 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 52, 52 -> 52
			// srcs: (1825, 61)(1094) -2, (4230) 47 --> (5014) -49:NW3, ALU, -, NW3
			10'd44 : rdata = 48'b000100100000001100111111111000000100110000000000;
			// PEs: 48, 52 -> 52
			// srcs: (1899, 32)(3140) 47, (389) -2 --> (3526) -94:PEGB0, ND11, *, NI0
			10'd45 : rdata = 48'b000111110000000001100001011100000000000000000000;
			// PEs: 48, 52 -> 53
			// srcs: (1901, 33)(3140) 47, (391) -3 --> (3528) -141:PEGB0, ND4, *, PENB
			10'd46 : rdata = 48'b000111110000000001100000100000000000000100000000;
			// PEs: 52, 52 -> 52
			// srcs: (1902, 47)(3) 1, (3526) -94 --> (4310) -94:NM0, NI0, *, NI1
			10'd47 : rdata = 48'b000111000000000010100000000100001000000000000000;
			// PEs: 52, 51 -> 51
			// srcs: (1903, 48)(3) 1, (3527) 0 --> (4311) 0:NM0, PENB, *, PEGB3
			10'd48 : rdata = 48'b000111000000000011011111110000000000000010110000;
			// PEs: 52, 52 -> 52
			// srcs: (1905, 62)(1174) -2, (4310) -94 --> (5094) 92:NW11, NI1, -, NW11
			10'd49 : rdata = 48'b000100100000101110100000001000000110110000000000;
			// PEs: 52, 53 -> 52
			// srcs: (1910, 63)(1176) 0, (4312) -141 --> (5096) 141:NW4, PEGB5, -, NW4
			10'd50 : rdata = 48'b000100100000010011100001010000000101000000000000;
			// PEs: 48, 52 -> 53
			// srcs: (1981, 34)(3140) 47, (471) -2 --> (3608) -94:PEGB0, ND5, *, PENB
			10'd51 : rdata = 48'b000111110000000001100000101000000000000100000000;
			// PEs: 52, 51 -> 51
			// srcs: (1983, 49)(3) 1, (3607) -141 --> (4391) -141:NM0, PENB, *, PEGB3
			10'd52 : rdata = 48'b000111000000000011011111110000000000000010110000;
			// PEs: 52, 53 -> 52
			// srcs: (1990, 64)(1256) 0, (4392) -94 --> (5176) 94:NW5, PEGB5, -, NW5
			10'd53 : rdata = 48'b000100100000010111100001010000000101010000000000;
			// PEs: 48, 52 -> 53
			// srcs: (2061, 35)(3140) 47, (551) -3 --> (3688) -141:PEGB0, ND6, *, PENB
			10'd54 : rdata = 48'b000111110000000001100000110000000000000100000000;
			// PEs: 52, 51 -> 51
			// srcs: (2063, 50)(3) 1, (3687) -94 --> (4471) -94:NM0, PENB, *, PEGB3
			10'd55 : rdata = 48'b000111000000000011011111110000000000000010110000;
			// PEs: 52, 53 -> 52
			// srcs: (2070, 65)(1336) -3, (4472) -141 --> (5256) 138:NW6, PEGB5, -, NW6
			10'd56 : rdata = 48'b000100100000011011100001010000000101100000000000;
			// PEs: 48, 52 -> 
			// srcs: (2083, 36)(3140) 47, (573) 1 --> (3710) 47:PEGB0, ND12, *, 
			10'd57 : rdata = 48'b000111110000000001100001100000000000000000000000;
			// PEs: 52, 52 -> 
			// srcs: (2086, 51)(3) 1, (3710) 47 --> (4494) 47:NM0, ALU, *, 
			10'd58 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 52, 52 -> 52
			// srcs: (2089, 66)(1358) -2, (4494) 47 --> (5278) -49:NW12, ALU, -, NW12
			10'd59 : rdata = 48'b000100100000110000111111111000000111000000000000;
			// PEs: 48, 52 -> 52
			// srcs: (2143, 37)(3140) 47, (633) -2 --> (3770) -94:PEGB0, ND7, *, NI0
			10'd60 : rdata = 48'b000111110000000001100000111100000000000000000000;
			// PEs: 52, 51 -> 51
			// srcs: (2145, 52)(3) 1, (3769) -47 --> (4553) -47:NM0, PENB, *, PEGB3
			10'd61 : rdata = 48'b000111000000000011011111110000000000000010110000;
			// PEs: 52, 52 -> 
			// srcs: (2146, 53)(3) 1, (3770) -94 --> (4554) -94:NM0, NI0, *, 
			10'd62 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 52, 52 -> 52
			// srcs: (2149, 67)(1418) -1, (4554) -94 --> (5338) 93:NW7, ALU, -, NW7
			10'd63 : rdata = 48'b000100100000011100111111111000000101110000000000;
			// PEs: 48, 52 -> 53
			// srcs: (2223, 38)(3140) 47, (713) -2 --> (3850) -94:PEGB0, ND8, *, PENB
			10'd64 : rdata = 48'b000111110000000001100001000000000000000100000000;
			// PEs: 52, 51 -> 51
			// srcs: (2225, 54)(3) 1, (3849) 94 --> (4633) 94:NM0, PENB, *, PEGB3
			10'd65 : rdata = 48'b000111000000000011011111110000000000000010110000;
			// PEs: 52, 53 -> 52
			// srcs: (2232, 68)(1498) -1, (4634) -94 --> (5418) 93:NW8, PEGB5, -, NW8
			10'd66 : rdata = 48'b000100100000100011100001010000000110000000000000;
			// PEs: 48, 52 -> 
			// srcs: (2267, 39)(3140) 47, (757) -2 --> (3894) -94:PEGB0, ND13, *, 
			10'd67 : rdata = 48'b000111110000000001100001101000000000000000000000;
			// PEs: 52, 52 -> 
			// srcs: (2270, 55)(3) 1, (3894) -94 --> (4678) -94:NM0, ALU, *, 
			10'd68 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 52, 52 -> 52
			// srcs: (2273, 69)(1542) 1, (4678) -94 --> (5462) 95:NW13, ALU, -, NW13
			10'd69 : rdata = 48'b000100100000110100111111111000000111010000000000;
			default : rdata = 48'b000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 53) begin
	always @(*) begin
		case(address)
			// PEs: 53, 53 -> 48
			// srcs: (1, 0)(69) 1, (854) 0 --> (1638) 0:ND0, NW0, *, PEGB0
			10'd0 : rdata = 48'b000110110000000001000000000000000000000010000000;
			// PEs: 53, 53 -> 53
			// srcs: (2, 1)(151) -2, (936) -3 --> (1720) 6:ND1, NW1, *, NI0
			10'd1 : rdata = 48'b000110110000000101000000001100000000000000000000;
			// PEs: 53, 53 -> 48
			// srcs: (3, 2)(231) 2, (1016) -1 --> (1800) -2:ND2, NW2, *, PEGB0
			10'd2 : rdata = 48'b000110110000001001000000010000000000000010000000;
			// PEs: 53, 53 -> 48
			// srcs: (4, 3)(311) 1, (1096) -1 --> (1880) -1:ND3, NW3, *, PEGB0
			10'd3 : rdata = 48'b000110110000001101000000011000000000000010000000;
			// PEs: 53, 53 -> 48
			// srcs: (5, 4)(393) -3, (1178) -2 --> (1962) 6:ND4, NW4, *, PEGB0
			10'd4 : rdata = 48'b000110110000010001000000100000000000000010000000;
			// PEs: 53, 53 -> 48
			// srcs: (6, 5)(473) -2, (1258) -1 --> (2042) 2:ND5, NW5, *, PEGB0
			10'd5 : rdata = 48'b000110110000010101000000101000000000000010000000;
			// PEs: 53, 53 -> 48
			// srcs: (7, 6)(553) -1, (1338) 0 --> (2122) 0:ND6, NW6, *, PEGB0
			10'd6 : rdata = 48'b000110110000011001000000110000000000000010000000;
			// PEs: 53, 53 -> 48
			// srcs: (8, 7)(635) 1, (1420) -3 --> (2204) -3:ND7, NW7, *, PEGB0
			10'd7 : rdata = 48'b000110110000011101000000111000000000000010000000;
			// PEs: 53, 53 -> 55
			// srcs: (9, 8)(715) 2, (1500) -1 --> (2284) -2:ND8, NW8, *, PEGB7
			10'd8 : rdata = 48'b000110110000100001000001000000000000000011110000;
			// PEs: 53, 53 -> 49
			// srcs: (10, 9)(28) 0, (813) 0 --> (1597) 0:ND9, NW9, *, PEGB1
			10'd9 : rdata = 48'b000110110000100101000001001000000000000010010000;
			// PEs: 53, 53 -> 49
			// srcs: (11, 10)(212) 2, (997) 2 --> (1781) 4:ND10, NW10, *, PEGB1
			10'd10 : rdata = 48'b000110110000101001000001010000000000000010010000;
			// PEs: 53, 53 -> 53
			// srcs: (12, 11)(392) -1, (1177) -3 --> (1961) 3:ND11, NW11, *, NI1
			10'd11 : rdata = 48'b000110110000101101000001011100001000000000000000;
			// PEs: 53, 53 -> 53
			// srcs: (13, 12)(576) -1, (1361) -1 --> (2145) 1:ND12, NW12, *, NI2
			10'd12 : rdata = 48'b000110110000110001000001100100010000000000000000;
			// PEs: 53, 53 -> 53
			// srcs: (14, 13)(760) 2, (1545) -2 --> (2329) -4:ND13, NW13, *, NI3
			10'd13 : rdata = 48'b000110110000110101000001101100011000000000000000;
			// PEs: 51, 52 -> 53
			// srcs: (15, 16)(2281) -6, (2282) 2 --> (3059) -4:PEGB3, PENB, +, NI4
			10'd14 : rdata = 48'b000011110000011011011111110100100000000000000000;
			// PEs: 48 -> 
			// srcs: (31, 14)(1712) -6 --> (1712) -6:PEGB0, pass, 
			10'd15 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 48, 53 -> 53
			// srcs: (40, 15)(1711) 0, (1712) -6 --> (2491) -6:PEGB0, ALU, +, NI5
			10'd16 : rdata = 48'b000011110000000000111111111100101000000000000000;
			// PEs: 49 -> 
			// srcs: (95, 19)(2732) 0 --> (2732) 0:PEGB1, pass, 
			10'd17 : rdata = 48'b110001110000001000000000000000000000000000000000;
			// PEs: 53, 51 -> 53
			// srcs: (98, 20)(2732) 0, (1955) 0 --> (2733) 0:ALU, PEGB3, +, NI6
			10'd18 : rdata = 48'b000010011111111111100000110100110000000000000000;
			// PEs: 53 -> 48
			// srcs: (105, 17)(1720) 6 --> (1720) 6:NI0, pass, PEGB0
			10'd19 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 53 -> 48
			// srcs: (128, 18)(2491) -6 --> (2491) -6:NI5, pass, PEGB0
			10'd20 : rdata = 48'b110001010000010100000000000000000000000010000000;
			// PEs: 53 -> 48
			// srcs: (142, 22)(2145) 1 --> (2145) 1:NI2, pass, PEGB0
			10'd21 : rdata = 48'b110001010000001000000000000000000000000010000000;
			// PEs: 53 -> 48
			// srcs: (145, 21)(1961) 3 --> (1961) 3:NI1, pass, PEGB0
			10'd22 : rdata = 48'b110001010000000100000000000000000000000010000000;
			// PEs: 53 -> 48
			// srcs: (148, 23)(3059) -4 --> (3059) -4:NI4, pass, PEGB0
			10'd23 : rdata = 48'b110001010000010000000000000000000000000010000000;
			// PEs: 53 -> 48
			// srcs: (149, 24)(2329) -4 --> (2329) -4:NI3, pass, PEGB0
			10'd24 : rdata = 48'b110001010000001100000000000000000000000010000000;
			// PEs: 53 -> 48
			// srcs: (376, 25)(2733) 0 --> (2733) 0:NI6, pass, PEGB0
			10'd25 : rdata = 48'b110001010000011000000000000000000000000010000000;
			// PEs: 48, 53 -> 
			// srcs: (1538, 26)(3140) 47, (28) 0 --> (3165) 0:PEGB0, ND9, *, 
			10'd26 : rdata = 48'b000111110000000001100001001000000000000000000000;
			// PEs: 53, 53 -> 
			// srcs: (1541, 40)(3) 1, (3165) 0 --> (3949) 0:NM0, ALU, *, 
			10'd27 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 53, 53 -> 53
			// srcs: (1544, 56)(813) 0, (3949) 0 --> (4733) 0:NW9, ALU, -, NW9
			10'd28 : rdata = 48'b000100100000100100111111111000000110010000000000;
			// PEs: 48, 53 -> 54
			// srcs: (1579, 27)(3140) 47, (69) 1 --> (3206) 47:PEGB0, ND0, *, PENB
			10'd29 : rdata = 48'b000111110000000001100000000000000000000100000000;
			// PEs: 53, 52 -> 52
			// srcs: (1580, 41)(3) 1, (3204) 47 --> (3988) 47:NM0, PENB, *, PEGB4
			10'd30 : rdata = 48'b000111000000000011011111110000000000000011000000;
			// PEs: 53, 54 -> 53
			// srcs: (1588, 57)(854) 0, (3990) 47 --> (4774) -47:NW0, PEGB6, -, NW0
			10'd31 : rdata = 48'b000100100000000011100001100000000100000000000000;
			// PEs: 48, 53 -> 54
			// srcs: (1661, 28)(3140) 47, (151) -2 --> (3288) -94:PEGB0, ND1, *, PENB
			10'd32 : rdata = 48'b000111110000000001100000001000000000000100000000;
			// PEs: 53, 52 -> 52
			// srcs: (1662, 42)(3) 1, (3286) 94 --> (4070) 94:NM0, PENB, *, PEGB4
			10'd33 : rdata = 48'b000111000000000011011111110000000000000011000000;
			// PEs: 53, 54 -> 53
			// srcs: (1670, 58)(936) -3, (4072) -94 --> (4856) 91:NW1, PEGB6, -, NW1
			10'd34 : rdata = 48'b000100100000000111100001100000000100010000000000;
			// PEs: 48, 53 -> 
			// srcs: (1722, 29)(3140) 47, (212) 2 --> (3349) 94:PEGB0, ND10, *, 
			10'd35 : rdata = 48'b000111110000000001100001010000000000000000000000;
			// PEs: 53, 53 -> 
			// srcs: (1725, 43)(3) 1, (3349) 94 --> (4133) 94:NM0, ALU, *, 
			10'd36 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 53, 53 -> 53
			// srcs: (1728, 59)(997) 2, (4133) 94 --> (4917) -92:NW10, ALU, -, NW10
			10'd37 : rdata = 48'b000100100000101000111111111000000110100000000000;
			// PEs: 48, 53 -> 53
			// srcs: (1741, 30)(3140) 47, (231) 2 --> (3368) 94:PEGB0, ND2, *, NI0
			10'd38 : rdata = 48'b000111110000000001100000010100000000000000000000;
			// PEs: 53, 52 -> 52
			// srcs: (1742, 44)(3) 1, (3366) 47 --> (4150) 47:NM0, PENB, *, PEGB4
			10'd39 : rdata = 48'b000111000000000011011111110000000000000011000000;
			// PEs: 53, 53 -> 
			// srcs: (1744, 45)(3) 1, (3368) 94 --> (4152) 94:NM0, NI0, *, 
			10'd40 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 53, 53 -> 53
			// srcs: (1747, 60)(1016) -1, (4152) 94 --> (4936) -95:NW2, ALU, -, NW2
			10'd41 : rdata = 48'b000100100000001000111111111000000100100000000000;
			// PEs: 48, 53 -> 
			// srcs: (1821, 31)(3140) 47, (311) 1 --> (3448) 47:PEGB0, ND3, *, 
			10'd42 : rdata = 48'b000111110000000001100000011000000000000000000000;
			// PEs: 53, 53 -> 
			// srcs: (1824, 46)(3) 1, (3448) 47 --> (4232) 47:NM0, ALU, *, 
			10'd43 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 53, 53 -> 53
			// srcs: (1827, 61)(1096) -1, (4232) 47 --> (5016) -48:NW3, ALU, -, NW3
			10'd44 : rdata = 48'b000100100000001100111111111000000100110000000000;
			// PEs: 48, 53 -> 53
			// srcs: (1902, 32)(3140) 47, (392) -1 --> (3529) -47:PEGB0, ND11, *, NI0
			10'd45 : rdata = 48'b000111110000000001100001011100000000000000000000;
			// PEs: 48, 53 -> 54
			// srcs: (1903, 33)(3140) 47, (393) -3 --> (3530) -141:PEGB0, ND4, *, PENB
			10'd46 : rdata = 48'b000111110000000001100000100000000000000100000000;
			// PEs: 53, 52 -> 52
			// srcs: (1904, 47)(3) 1, (3528) -141 --> (4312) -141:NM0, PENB, *, PEGB4
			10'd47 : rdata = 48'b000111000000000011011111110000000000000011000000;
			// PEs: 53, 53 -> 
			// srcs: (1905, 48)(3) 1, (3529) -47 --> (4313) -47:NM0, NI0, *, 
			10'd48 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 53, 53 -> 53
			// srcs: (1908, 62)(1177) -3, (4313) -47 --> (5097) 44:NW11, ALU, -, NW11
			10'd49 : rdata = 48'b000100100000101100111111111000000110110000000000;
			// PEs: 53, 54 -> 53
			// srcs: (1912, 63)(1178) -2, (4314) -141 --> (5098) 139:NW4, PEGB6, -, NW4
			10'd50 : rdata = 48'b000100100000010011100001100000000101000000000000;
			// PEs: 48, 53 -> 54
			// srcs: (1983, 34)(3140) 47, (473) -2 --> (3610) -94:PEGB0, ND5, *, PENB
			10'd51 : rdata = 48'b000111110000000001100000101000000000000100000000;
			// PEs: 53, 52 -> 52
			// srcs: (1984, 49)(3) 1, (3608) -94 --> (4392) -94:NM0, PENB, *, PEGB4
			10'd52 : rdata = 48'b000111000000000011011111110000000000000011000000;
			// PEs: 53, 54 -> 53
			// srcs: (1992, 64)(1258) -1, (4394) -94 --> (5178) 93:NW5, PEGB6, -, NW5
			10'd53 : rdata = 48'b000100100000010111100001100000000101010000000000;
			// PEs: 48, 53 -> 53
			// srcs: (2063, 35)(3140) 47, (553) -1 --> (3690) -47:PEGB0, ND6, *, NI0
			10'd54 : rdata = 48'b000111110000000001100000110100000000000000000000;
			// PEs: 53, 52 -> 52
			// srcs: (2064, 50)(3) 1, (3688) -141 --> (4472) -141:NM0, PENB, *, PEGB4
			10'd55 : rdata = 48'b000111000000000011011111110000000000000011000000;
			// PEs: 53, 53 -> 
			// srcs: (2066, 51)(3) 1, (3690) -47 --> (4474) -47:NM0, NI0, *, 
			10'd56 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 53, 53 -> 53
			// srcs: (2069, 65)(1338) 0, (4474) -47 --> (5258) 47:NW6, ALU, -, NW6
			10'd57 : rdata = 48'b000100100000011000111111111000000101100000000000;
			// PEs: 48, 53 -> 
			// srcs: (2086, 36)(3140) 47, (576) -1 --> (3713) -47:PEGB0, ND12, *, 
			10'd58 : rdata = 48'b000111110000000001100001100000000000000000000000;
			// PEs: 53, 53 -> 
			// srcs: (2089, 52)(3) 1, (3713) -47 --> (4497) -47:NM0, ALU, *, 
			10'd59 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 53, 53 -> 53
			// srcs: (2092, 66)(1361) -1, (4497) -47 --> (5281) 46:NW12, ALU, -, NW12
			10'd60 : rdata = 48'b000100100000110000111111111000000111000000000000;
			// PEs: 48, 53 -> 
			// srcs: (2145, 37)(3140) 47, (635) 1 --> (3772) 47:PEGB0, ND7, *, 
			10'd61 : rdata = 48'b000111110000000001100000111000000000000000000000;
			// PEs: 53, 53 -> 
			// srcs: (2148, 53)(3) 1, (3772) 47 --> (4556) 47:NM0, ALU, *, 
			10'd62 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 53, 53 -> 53
			// srcs: (2151, 67)(1420) -3, (4556) 47 --> (5340) -50:NW7, ALU, -, NW7
			10'd63 : rdata = 48'b000100100000011100111111111000000101110000000000;
			// PEs: 48, 53 -> 54
			// srcs: (2225, 38)(3140) 47, (715) 2 --> (3852) 94:PEGB0, ND8, *, PENB
			10'd64 : rdata = 48'b000111110000000001100001000000000000000100000000;
			// PEs: 53, 52 -> 52
			// srcs: (2226, 54)(3) 1, (3850) -94 --> (4634) -94:NM0, PENB, *, PEGB4
			10'd65 : rdata = 48'b000111000000000011011111110000000000000011000000;
			// PEs: 53, 54 -> 53
			// srcs: (2234, 68)(1500) -1, (4636) 94 --> (5420) -95:NW8, PEGB6, -, NW8
			10'd66 : rdata = 48'b000100100000100011100001100000000110000000000000;
			// PEs: 48, 53 -> 
			// srcs: (2270, 39)(3140) 47, (760) 2 --> (3897) 94:PEGB0, ND13, *, 
			10'd67 : rdata = 48'b000111110000000001100001101000000000000000000000;
			// PEs: 53, 53 -> 
			// srcs: (2273, 55)(3) 1, (3897) 94 --> (4681) 94:NM0, ALU, *, 
			10'd68 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 53, 53 -> 53
			// srcs: (2276, 69)(1545) -2, (4681) 94 --> (5465) -96:NW13, ALU, -, NW13
			10'd69 : rdata = 48'b000100100000110100111111111000000111010000000000;
			default : rdata = 48'b000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 54) begin
	always @(*) begin
		case(address)
			// PEs: 54, 54 -> 48
			// srcs: (1, 0)(70) -1, (855) -3 --> (1639) 3:ND0, NW0, *, PEGB0
			10'd0 : rdata = 48'b000110110000000001000000000000000000000010000000;
			// PEs: 54, 54 -> 54
			// srcs: (2, 1)(152) -1, (937) -1 --> (1721) 1:ND1, NW1, *, NI0
			10'd1 : rdata = 48'b000110110000000101000000001100000000000000000000;
			// PEs: 54, 54 -> 48
			// srcs: (3, 2)(232) 0, (1017) 2 --> (1801) 0:ND2, NW2, *, PEGB0
			10'd2 : rdata = 48'b000110110000001001000000010000000000000010000000;
			// PEs: 54, 54 -> 48
			// srcs: (4, 3)(312) -1, (1097) -1 --> (1881) 1:ND3, NW3, *, PEGB0
			10'd3 : rdata = 48'b000110110000001101000000011000000000000010000000;
			// PEs: 54, 54 -> 48
			// srcs: (5, 4)(394) 0, (1179) 1 --> (1963) 0:ND4, NW4, *, PEGB0
			10'd4 : rdata = 48'b000110110000010001000000100000000000000010000000;
			// PEs: 54, 54 -> 48
			// srcs: (6, 5)(474) -3, (1259) -1 --> (2043) 3:ND5, NW5, *, PEGB0
			10'd5 : rdata = 48'b000110110000010101000000101000000000000010000000;
			// PEs: 54, 54 -> 48
			// srcs: (7, 6)(554) -2, (1339) -3 --> (2123) 6:ND6, NW6, *, PEGB0
			10'd6 : rdata = 48'b000110110000011001000000110000000000000010000000;
			// PEs: 54, 54 -> 48
			// srcs: (8, 7)(636) -1, (1421) -2 --> (2205) 2:ND7, NW7, *, PEGB0
			10'd7 : rdata = 48'b000110110000011101000000111000000000000010000000;
			// PEs: 54, 54 -> 55
			// srcs: (9, 8)(716) -2, (1501) 0 --> (2285) 0:ND8, NW8, *, PENB
			10'd8 : rdata = 48'b000110110000100001000001000000000000000100000000;
			// PEs: 54, 54 -> 48
			// srcs: (10, 9)(31) 2, (816) -1 --> (1600) -2:ND9, NW9, *, PEGB0
			10'd9 : rdata = 48'b000110110000100101000001001000000000000010000000;
			// PEs: 54, 54 -> 54
			// srcs: (11, 10)(215) -2, (1000) 0 --> (1784) 0:ND10, NW10, *, NI1
			10'd10 : rdata = 48'b000110110000101001000001010100001000000000000000;
			// PEs: 54, 54 -> 54
			// srcs: (12, 11)(395) -3, (1180) -3 --> (1964) 9:ND11, NW11, *, NI2
			10'd11 : rdata = 48'b000110110000101101000001011100010000000000000000;
			// PEs: 54, 54 -> 54
			// srcs: (13, 12)(579) 1, (1364) 0 --> (2148) 0:ND12, NW12, *, NI3
			10'd12 : rdata = 48'b000110110000110001000001100100011000000000000000;
			// PEs: 54, 54 -> 54
			// srcs: (14, 13)(763) 1, (1548) -3 --> (2332) -3:ND13, NW13, *, NI4
			10'd13 : rdata = 48'b000110110000110101000001101100100000000000000000;
			// PEs: 48 -> 
			// srcs: (39, 14)(1783) 2 --> (1783) 2:PEGB0, pass, 
			10'd14 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 48, 54 -> 
			// srcs: (48, 15)(1782) 3, (1783) 2 --> (2564) 5:PEGB0, ALU, +, 
			10'd15 : rdata = 48'b000011110000000000111111111000000000000000000000;
			// PEs: 54, 54 -> 55
			// srcs: (51, 19)(2564) 5, (1784) 0 --> (2565) 5:ALU, NI1, +, PENB
			10'd16 : rdata = 48'b000010011111111110100000001000000000000100000000;
			// PEs: 54 -> 48
			// srcs: (113, 18)(1721) 1 --> (1721) 1:NI0, pass, PEGB0
			10'd17 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 54 -> 48
			// srcs: (153, 20)(1964) 9 --> (1964) 9:NI2, pass, PEGB0
			10'd18 : rdata = 48'b110001010000001000000000000000000000000010000000;
			// PEs: 48 -> 
			// srcs: (242, 16)(1574) 3 --> (1574) 3:PEGB0, pass, 
			10'd19 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 48, 54 -> 49
			// srcs: (251, 17)(1573) 6, (1574) 3 --> (2357) 9:PEGB0, ALU, +, PEGB1
			10'd20 : rdata = 48'b000011110000000000111111111000000000000010010000;
			// PEs: 54 -> 49
			// srcs: (419, 21)(2148) 0 --> (2148) 0:NI3, pass, PEGB1
			10'd21 : rdata = 48'b110001010000001100000000000000000000000010010000;
			// PEs: 54 -> 49
			// srcs: (576, 22)(2332) -3 --> (2332) -3:NI4, pass, PEGB1
			10'd22 : rdata = 48'b110001010000010000000000000000000000000010010000;
			// PEs: 48 -> 
			// srcs: (593, 23)(2636) 2 --> (2636) 2:PEGB0, pass, 
			10'd23 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 54, 49 -> 49
			// srcs: (595, 24)(2636) 2, (2638) -2 --> (2639) 0:ALU, PEGB1, +, PEGB1
			10'd24 : rdata = 48'b000010011111111111100000010000000000000010010000;
			// PEs: 48, 54 -> 
			// srcs: (1541, 25)(3140) 47, (31) 2 --> (3168) 94:PEGB0, ND9, *, 
			10'd25 : rdata = 48'b000111110000000001100001001000000000000000000000;
			// PEs: 54, 54 -> 
			// srcs: (1544, 39)(3) 1, (3168) 94 --> (3952) 94:NM0, ALU, *, 
			10'd26 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 54, 54 -> 54
			// srcs: (1547, 56)(816) -1, (3952) 94 --> (4736) -95:NW9, ALU, -, NW9
			10'd27 : rdata = 48'b000100100000100100111111111000000110010000000000;
			// PEs: 48, 54 -> 54
			// srcs: (1580, 26)(3140) 47, (70) -1 --> (3207) -47:PEGB0, ND0, *, NI0
			10'd28 : rdata = 48'b000111110000000001100000000100000000000000000000;
			// PEs: 54, 53 -> 53
			// srcs: (1582, 40)(3) 1, (3206) 47 --> (3990) 47:NM0, PENB, *, PEGB5
			10'd29 : rdata = 48'b000111000000000011011111110000000000000011010000;
			// PEs: 54, 54 -> 
			// srcs: (1583, 41)(3) 1, (3207) -47 --> (3991) -47:NM0, NI0, *, 
			10'd30 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 54, 54 -> 54
			// srcs: (1586, 57)(855) -3, (3991) -47 --> (4775) 44:NW0, ALU, -, NW0
			10'd31 : rdata = 48'b000100100000000000111111111000000100000000000000;
			// PEs: 48, 54 -> 54
			// srcs: (1662, 27)(3140) 47, (152) -1 --> (3289) -47:PEGB0, ND1, *, NI0
			10'd32 : rdata = 48'b000111110000000001100000001100000000000000000000;
			// PEs: 54, 53 -> 53
			// srcs: (1664, 42)(3) 1, (3288) -94 --> (4072) -94:NM0, PENB, *, PEGB5
			10'd33 : rdata = 48'b000111000000000011011111110000000000000011010000;
			// PEs: 54, 54 -> 
			// srcs: (1665, 43)(3) 1, (3289) -47 --> (4073) -47:NM0, NI0, *, 
			10'd34 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 54, 54 -> 54
			// srcs: (1668, 58)(937) -1, (4073) -47 --> (4857) 46:NW1, ALU, -, NW1
			10'd35 : rdata = 48'b000100100000000100111111111000000100010000000000;
			// PEs: 48, 54 -> 
			// srcs: (1725, 28)(3140) 47, (215) -2 --> (3352) -94:PEGB0, ND10, *, 
			10'd36 : rdata = 48'b000111110000000001100001010000000000000000000000;
			// PEs: 54, 54 -> 
			// srcs: (1728, 44)(3) 1, (3352) -94 --> (4136) -94:NM0, ALU, *, 
			10'd37 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 54, 54 -> 54
			// srcs: (1731, 59)(1000) 0, (4136) -94 --> (4920) 94:NW10, ALU, -, NW10
			10'd38 : rdata = 48'b000100100000101000111111111000000110100000000000;
			// PEs: 48, 54 -> 
			// srcs: (1742, 29)(3140) 47, (232) 0 --> (3369) 0:PEGB0, ND2, *, 
			10'd39 : rdata = 48'b000111110000000001100000010000000000000000000000;
			// PEs: 54, 54 -> 
			// srcs: (1745, 45)(3) 1, (3369) 0 --> (4153) 0:NM0, ALU, *, 
			10'd40 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 54, 54 -> 54
			// srcs: (1748, 60)(1017) 2, (4153) 0 --> (4937) 2:NW2, ALU, -, NW2
			10'd41 : rdata = 48'b000100100000001000111111111000000100100000000000;
			// PEs: 48, 54 -> 
			// srcs: (1822, 30)(3140) 47, (312) -1 --> (3449) -47:PEGB0, ND3, *, 
			10'd42 : rdata = 48'b000111110000000001100000011000000000000000000000;
			// PEs: 54, 54 -> 
			// srcs: (1825, 46)(3) 1, (3449) -47 --> (4233) -47:NM0, ALU, *, 
			10'd43 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 54, 54 -> 54
			// srcs: (1828, 61)(1097) -1, (4233) -47 --> (5017) 46:NW3, ALU, -, NW3
			10'd44 : rdata = 48'b000100100000001100111111111000000100110000000000;
			// PEs: 48, 54 -> 55
			// srcs: (1904, 31)(3140) 47, (394) 0 --> (3531) 0:PEGB0, ND4, *, PENB
			10'd45 : rdata = 48'b000111110000000001100000100000000000000100000000;
			// PEs: 48, 54 -> 54
			// srcs: (1905, 32)(3140) 47, (395) -3 --> (3532) -141:PEGB0, ND11, *, NI0
			10'd46 : rdata = 48'b000111110000000001100001011100000000000000000000;
			// PEs: 54, 53 -> 53
			// srcs: (1906, 47)(3) 1, (3530) -141 --> (4314) -141:NM0, PENB, *, PEGB5
			10'd47 : rdata = 48'b000111000000000011011111110000000000000011010000;
			// PEs: 54, 54 -> 
			// srcs: (1908, 48)(3) 1, (3532) -141 --> (4316) -141:NM0, NI0, *, 
			10'd48 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 54, 54 -> 54
			// srcs: (1911, 63)(1180) -3, (4316) -141 --> (5100) 138:NW11, ALU, -, NW11
			10'd49 : rdata = 48'b000100100000101100111111111000000110110000000000;
			// PEs: 54, 55 -> 54
			// srcs: (1913, 62)(1179) 1, (4315) 0 --> (5099) 1:NW4, PEGB7, -, NW4
			10'd50 : rdata = 48'b000100100000010011100001110000000101000000000000;
			// PEs: 48, 54 -> 54
			// srcs: (1984, 33)(3140) 47, (474) -3 --> (3611) -141:PEGB0, ND5, *, NI0
			10'd51 : rdata = 48'b000111110000000001100000101100000000000000000000;
			// PEs: 54, 53 -> 53
			// srcs: (1986, 49)(3) 1, (3610) -94 --> (4394) -94:NM0, PENB, *, PEGB5
			10'd52 : rdata = 48'b000111000000000011011111110000000000000011010000;
			// PEs: 54, 54 -> 
			// srcs: (1987, 50)(3) 1, (3611) -141 --> (4395) -141:NM0, NI0, *, 
			10'd53 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 54, 54 -> 54
			// srcs: (1990, 64)(1259) -1, (4395) -141 --> (5179) 140:NW5, ALU, -, NW5
			10'd54 : rdata = 48'b000100100000010100111111111000000101010000000000;
			// PEs: 48, 54 -> 
			// srcs: (2064, 34)(3140) 47, (554) -2 --> (3691) -94:PEGB0, ND6, *, 
			10'd55 : rdata = 48'b000111110000000001100000110000000000000000000000;
			// PEs: 54, 54 -> 
			// srcs: (2067, 51)(3) 1, (3691) -94 --> (4475) -94:NM0, ALU, *, 
			10'd56 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 54, 54 -> 54
			// srcs: (2070, 65)(1339) -3, (4475) -94 --> (5259) 91:NW6, ALU, -, NW6
			10'd57 : rdata = 48'b000100100000011000111111111000000101100000000000;
			// PEs: 48, 54 -> 
			// srcs: (2089, 35)(3140) 47, (579) 1 --> (3716) 47:PEGB0, ND12, *, 
			10'd58 : rdata = 48'b000111110000000001100001100000000000000000000000;
			// PEs: 54, 54 -> 
			// srcs: (2092, 52)(3) 1, (3716) 47 --> (4500) 47:NM0, ALU, *, 
			10'd59 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 54, 54 -> 54
			// srcs: (2095, 66)(1364) 0, (4500) 47 --> (5284) -47:NW12, ALU, -, NW12
			10'd60 : rdata = 48'b000100100000110000111111111000000111000000000000;
			// PEs: 48, 54 -> 
			// srcs: (2146, 36)(3140) 47, (636) -1 --> (3773) -47:PEGB0, ND7, *, 
			10'd61 : rdata = 48'b000111110000000001100000111000000000000000000000;
			// PEs: 54, 54 -> 
			// srcs: (2149, 53)(3) 1, (3773) -47 --> (4557) -47:NM0, ALU, *, 
			10'd62 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 54, 54 -> 54
			// srcs: (2152, 67)(1421) -2, (4557) -47 --> (5341) 45:NW7, ALU, -, NW7
			10'd63 : rdata = 48'b000100100000011100111111111000000101110000000000;
			// PEs: 48, 54 -> 55
			// srcs: (2226, 37)(3140) 47, (716) -2 --> (3853) -94:PEGB0, ND8, *, PENB
			10'd64 : rdata = 48'b000111110000000001100001000000000000000100000000;
			// PEs: 54, 53 -> 53
			// srcs: (2228, 54)(3) 1, (3852) 94 --> (4636) 94:NM0, PENB, *, PEGB5
			10'd65 : rdata = 48'b000111000000000011011111110000000000000011010000;
			// PEs: 54, 55 -> 54
			// srcs: (2235, 68)(1501) 0, (4637) -94 --> (5421) 94:NW8, PEGB7, -, NW8
			10'd66 : rdata = 48'b000100100000100011100001110000000110000000000000;
			// PEs: 48, 54 -> 
			// srcs: (2273, 38)(3140) 47, (763) 1 --> (3900) 47:PEGB0, ND13, *, 
			10'd67 : rdata = 48'b000111110000000001100001101000000000000000000000;
			// PEs: 54, 54 -> 
			// srcs: (2276, 55)(3) 1, (3900) 47 --> (4684) 47:NM0, ALU, *, 
			10'd68 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 54, 54 -> 54
			// srcs: (2279, 69)(1548) -3, (4684) 47 --> (5468) -50:NW13, ALU, -, NW13
			10'd69 : rdata = 48'b000100100000110100111111111000000111010000000000;
			default : rdata = 48'b000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 55) begin
	always @(*) begin
		case(address)
			// PEs: 55, 55 -> 48
			// srcs: (1, 0)(72) 2, (857) -3 --> (1641) -6:ND0, NW0, *, PENB
			10'd0 : rdata = 48'b000110110000000001000000000000000000000100000000;
			// PEs: 55, 55 -> 55
			// srcs: (2, 1)(153) 2, (938) -3 --> (1722) -6:ND1, NW1, *, NI0
			10'd1 : rdata = 48'b000110110000000101000000001100000000000000000000;
			// PEs: 55, 55 -> 48
			// srcs: (3, 2)(234) -2, (1019) 0 --> (1803) 0:ND2, NW2, *, PENB
			10'd2 : rdata = 48'b000110110000001001000000010000000000000100000000;
			// PEs: 55, 55 -> 49
			// srcs: (4, 3)(314) 1, (1099) -1 --> (1883) -1:ND3, NW3, *, PEGB1
			10'd3 : rdata = 48'b000110110000001101000000011000000000000010010000;
			// PEs: 55, 55 -> 55
			// srcs: (5, 4)(396) -3, (1181) 1 --> (1965) -3:ND4, NW4, *, NI1
			10'd4 : rdata = 48'b000110110000010001000000100100001000000000000000;
			// PEs: 55, 55 -> 48
			// srcs: (6, 5)(476) -1, (1261) 2 --> (2045) -2:ND5, NW5, *, PENB
			10'd5 : rdata = 48'b000110110000010101000000101000000000000100000000;
			// PEs: 55, 55 -> 48
			// srcs: (7, 6)(556) 2, (1341) -1 --> (2125) -2:ND6, NW6, *, PENB
			10'd6 : rdata = 48'b000110110000011001000000110000000000000100000000;
			// PEs: 55, 55 -> 48
			// srcs: (8, 7)(638) 2, (1423) -2 --> (2207) -4:ND7, NW7, *, PENB
			10'd7 : rdata = 48'b000110110000011101000000111000000000000100000000;
			// PEs: 55, 55 -> 48
			// srcs: (9, 8)(718) 0, (1503) 2 --> (2287) 0:ND8, NW8, *, PENB
			10'd8 : rdata = 48'b000110110000100001000001000000000000000100000000;
			// PEs: 55, 55 -> 55
			// srcs: (10, 9)(34) -3, (819) 1 --> (1603) -3:ND9, NW9, *, NI2
			10'd9 : rdata = 48'b000110110000100101000001001100010000000000000000;
			// PEs: 55, 55 -> 55
			// srcs: (11, 10)(218) 1, (1003) -1 --> (1787) -1:ND10, NW10, *, NI3
			10'd10 : rdata = 48'b000110110000101001000001010100011000000000000000;
			// PEs: 55, 55 -> 55
			// srcs: (12, 11)(402) 2, (1187) -3 --> (1971) -6:ND11, NW11, *, NI4
			10'd11 : rdata = 48'b000110110000101101000001011100100000000000000000;
			// PEs: 55, 55 -> 55
			// srcs: (13, 12)(582) 0, (1367) 2 --> (2151) 0:ND12, NW12, *, NI5
			10'd12 : rdata = 48'b000110110000110001000001100100101000000000000000;
			// PEs: 55, 55 -> 55
			// srcs: (14, 13)(766) 1, (1551) -2 --> (2335) -2:ND13, NW13, *, NI6
			10'd13 : rdata = 48'b000110110000110101000001101100110000000000000000;
			// PEs: 53, 54 -> 55
			// srcs: (15, 16)(2284) -2, (2285) 0 --> (3064) -2:PEGB5, PENB, +, NI7
			10'd14 : rdata = 48'b000011110000101011011111110100111000000000000000;
			// PEs: 48 -> 
			// srcs: (43, 14)(1786) 2 --> (1786) 2:PEGB0, pass, 
			10'd15 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 48, 55 -> 
			// srcs: (52, 15)(1785) 2, (1786) 2 --> (2566) 4:PEGB0, ALU, +, 
			10'd16 : rdata = 48'b000011110000000000111111111000000000000000000000;
			// PEs: 55, 55 -> 
			// srcs: (55, 20)(2566) 4, (1787) -1 --> (2567) 3:ALU, NI3, +, 
			10'd17 : rdata = 48'b000010011111111110100000011000000000000000000000;
			// PEs: 54, 55 -> 55
			// srcs: (58, 25)(2565) 5, (2567) 3 --> (2568) 8:PENB, ALU, +, NI3
			10'd18 : rdata = 48'b000011101111111000111111111100011000000000000000;
			// PEs: 55 -> 48
			// srcs: (105, 17)(1722) -6 --> (1722) -6:NI0, pass, PENB
			10'd19 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 55 -> 48
			// srcs: (113, 19)(1603) -3 --> (1603) -3:NI2, pass, PENB
			10'd20 : rdata = 48'b110001010000001000000000000000000000000100000000;
			// PEs: 55 -> 48
			// srcs: (121, 18)(1965) -3 --> (1965) -3:NI1, pass, PENB
			10'd21 : rdata = 48'b110001010000000100000000000000000000000100000000;
			// PEs: 55 -> 48
			// srcs: (133, 21)(1971) -6 --> (1971) -6:NI4, pass, PENB
			10'd22 : rdata = 48'b110001010000010000000000000000000000000100000000;
			// PEs: 55 -> 48
			// srcs: (142, 22)(2151) 0 --> (2151) 0:NI5, pass, PENB
			10'd23 : rdata = 48'b110001010000010100000000000000000000000100000000;
			// PEs: 55 -> 48
			// srcs: (151, 23)(3064) -2 --> (3064) -2:NI7, pass, PENB
			10'd24 : rdata = 48'b110001010000011100000000000000000000000100000000;
			// PEs: 55 -> 48
			// srcs: (158, 24)(2335) -2 --> (2335) -2:NI6, pass, PENB
			10'd25 : rdata = 48'b110001010000011000000000000000000000000100000000;
			// PEs: 55 -> 48
			// srcs: (598, 26)(2568) 8 --> (2568) 8:NI3, pass, PENB
			10'd26 : rdata = 48'b110001010000001100000000000000000000000100000000;
			// PEs: 48, 55 -> 
			// srcs: (1544, 27)(3140) 47, (34) -3 --> (3171) -141:PEGB0, ND9, *, 
			10'd27 : rdata = 48'b000111110000000001100001001000000000000000000000;
			// PEs: 55, 55 -> 
			// srcs: (1547, 41)(3) 1, (3171) -141 --> (3955) -141:NM0, ALU, *, 
			10'd28 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 55, 55 -> 55
			// srcs: (1550, 57)(819) 1, (3955) -141 --> (4739) 142:NW9, ALU, -, NW9
			10'd29 : rdata = 48'b000100100000100100111111111000000110010000000000;
			// PEs: 48, 55 -> 
			// srcs: (1582, 28)(3140) 47, (72) 2 --> (3209) 94:PEGB0, ND0, *, 
			10'd30 : rdata = 48'b000111110000000001100000000000000000000000000000;
			// PEs: 55, 55 -> 
			// srcs: (1585, 42)(3) 1, (3209) 94 --> (3993) 94:NM0, ALU, *, 
			10'd31 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 55, 55 -> 55
			// srcs: (1588, 58)(857) -3, (3993) 94 --> (4777) -97:NW0, ALU, -, NW0
			10'd32 : rdata = 48'b000100100000000000111111111000000100000000000000;
			// PEs: 48, 55 -> 
			// srcs: (1663, 29)(3140) 47, (153) 2 --> (3290) 94:PEGB0, ND1, *, 
			10'd33 : rdata = 48'b000111110000000001100000001000000000000000000000;
			// PEs: 55, 55 -> 
			// srcs: (1666, 43)(3) 1, (3290) 94 --> (4074) 94:NM0, ALU, *, 
			10'd34 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 55, 55 -> 55
			// srcs: (1669, 59)(938) -3, (4074) 94 --> (4858) -97:NW1, ALU, -, NW1
			10'd35 : rdata = 48'b000100100000000100111111111000000100010000000000;
			// PEs: 48, 55 -> 
			// srcs: (1728, 30)(3140) 47, (218) 1 --> (3355) 47:PEGB0, ND10, *, 
			10'd36 : rdata = 48'b000111110000000001100001010000000000000000000000;
			// PEs: 55, 55 -> 
			// srcs: (1731, 44)(3) 1, (3355) 47 --> (4139) 47:NM0, ALU, *, 
			10'd37 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 55, 55 -> 55
			// srcs: (1734, 60)(1003) -1, (4139) 47 --> (4923) -48:NW10, ALU, -, NW10
			10'd38 : rdata = 48'b000100100000101000111111111000000110100000000000;
			// PEs: 48, 55 -> 
			// srcs: (1744, 31)(3140) 47, (234) -2 --> (3371) -94:PEGB0, ND2, *, 
			10'd39 : rdata = 48'b000111110000000001100000010000000000000000000000;
			// PEs: 55, 55 -> 
			// srcs: (1747, 45)(3) 1, (3371) -94 --> (4155) -94:NM0, ALU, *, 
			10'd40 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 55, 55 -> 55
			// srcs: (1750, 61)(1019) 0, (4155) -94 --> (4939) 94:NW2, ALU, -, NW2
			10'd41 : rdata = 48'b000100100000001000111111111000000100100000000000;
			// PEs: 48, 55 -> 
			// srcs: (1824, 32)(3140) 47, (314) 1 --> (3451) 47:PEGB0, ND3, *, 
			10'd42 : rdata = 48'b000111110000000001100000011000000000000000000000;
			// PEs: 55, 55 -> 
			// srcs: (1827, 46)(3) 1, (3451) 47 --> (4235) 47:NM0, ALU, *, 
			10'd43 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 55, 55 -> 55
			// srcs: (1830, 62)(1099) -1, (4235) 47 --> (5019) -48:NW3, ALU, -, NW3
			10'd44 : rdata = 48'b000100100000001100111111111000000100110000000000;
			// PEs: 48, 55 -> 55
			// srcs: (1906, 33)(3140) 47, (396) -3 --> (3533) -141:PEGB0, ND4, *, NI0
			10'd45 : rdata = 48'b000111110000000001100000100100000000000000000000;
			// PEs: 55, 54 -> 54
			// srcs: (1907, 47)(3) 1, (3531) 0 --> (4315) 0:NM0, PENB, *, PEGB6
			10'd46 : rdata = 48'b000111000000000011011111110000000000000011100000;
			// PEs: 55, 55 -> 55
			// srcs: (1909, 48)(3) 1, (3533) -141 --> (4317) -141:NM0, NI0, *, NI1
			10'd47 : rdata = 48'b000111000000000010100000000100001000000000000000;
			// PEs: 48, 55 -> 55
			// srcs: (1912, 34)(3140) 47, (402) 2 --> (3539) 94:PEGB0, ND11, *, NI0
			10'd48 : rdata = 48'b000111110000000001100001011100000000000000000000;
			// PEs: 55, 55 -> 55
			// srcs: (1913, 63)(1181) 1, (4317) -141 --> (5101) 142:NW4, NI1, -, NW4
			10'd49 : rdata = 48'b000100100000010010100000001000000101000000000000;
			// PEs: 55, 55 -> 
			// srcs: (1915, 49)(3) 1, (3539) 94 --> (4323) 94:NM0, NI0, *, 
			10'd50 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 55, 55 -> 55
			// srcs: (1918, 64)(1187) -3, (4323) 94 --> (5107) -97:NW11, ALU, -, NW11
			10'd51 : rdata = 48'b000100100000101100111111111000000110110000000000;
			// PEs: 48, 55 -> 
			// srcs: (1986, 35)(3140) 47, (476) -1 --> (3613) -47:PEGB0, ND5, *, 
			10'd52 : rdata = 48'b000111110000000001100000101000000000000000000000;
			// PEs: 55, 55 -> 
			// srcs: (1989, 50)(3) 1, (3613) -47 --> (4397) -47:NM0, ALU, *, 
			10'd53 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 55, 55 -> 55
			// srcs: (1992, 65)(1261) 2, (4397) -47 --> (5181) 49:NW5, ALU, -, NW5
			10'd54 : rdata = 48'b000100100000010100111111111000000101010000000000;
			// PEs: 48, 55 -> 
			// srcs: (2066, 36)(3140) 47, (556) 2 --> (3693) 94:PEGB0, ND6, *, 
			10'd55 : rdata = 48'b000111110000000001100000110000000000000000000000;
			// PEs: 55, 55 -> 
			// srcs: (2069, 51)(3) 1, (3693) 94 --> (4477) 94:NM0, ALU, *, 
			10'd56 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 55, 55 -> 55
			// srcs: (2072, 66)(1341) -1, (4477) 94 --> (5261) -95:NW6, ALU, -, NW6
			10'd57 : rdata = 48'b000100100000011000111111111000000101100000000000;
			// PEs: 48, 55 -> 
			// srcs: (2092, 37)(3140) 47, (582) 0 --> (3719) 0:PEGB0, ND12, *, 
			10'd58 : rdata = 48'b000111110000000001100001100000000000000000000000;
			// PEs: 55, 55 -> 
			// srcs: (2095, 52)(3) 1, (3719) 0 --> (4503) 0:NM0, ALU, *, 
			10'd59 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 55, 55 -> 55
			// srcs: (2098, 67)(1367) 2, (4503) 0 --> (5287) 2:NW12, ALU, -, NW12
			10'd60 : rdata = 48'b000100100000110000111111111000000111000000000000;
			// PEs: 48, 55 -> 
			// srcs: (2148, 38)(3140) 47, (638) 2 --> (3775) 94:PEGB0, ND7, *, 
			10'd61 : rdata = 48'b000111110000000001100000111000000000000000000000;
			// PEs: 55, 55 -> 
			// srcs: (2151, 53)(3) 1, (3775) 94 --> (4559) 94:NM0, ALU, *, 
			10'd62 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 55, 55 -> 55
			// srcs: (2154, 68)(1423) -2, (4559) 94 --> (5343) -96:NW7, ALU, -, NW7
			10'd63 : rdata = 48'b000100100000011100111111111000000101110000000000;
			// PEs: 48, 55 -> 55
			// srcs: (2228, 39)(3140) 47, (718) 0 --> (3855) 0:PEGB0, ND8, *, NI0
			10'd64 : rdata = 48'b000111110000000001100001000100000000000000000000;
			// PEs: 55, 54 -> 54
			// srcs: (2229, 54)(3) 1, (3853) -94 --> (4637) -94:NM0, PENB, *, PEGB6
			10'd65 : rdata = 48'b000111000000000011011111110000000000000011100000;
			// PEs: 55, 55 -> 
			// srcs: (2231, 55)(3) 1, (3855) 0 --> (4639) 0:NM0, NI0, *, 
			10'd66 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 55, 55 -> 55
			// srcs: (2234, 69)(1503) 2, (4639) 0 --> (5423) 2:NW8, ALU, -, NW8
			10'd67 : rdata = 48'b000100100000100000111111111000000110000000000000;
			// PEs: 48, 55 -> 
			// srcs: (2276, 40)(3140) 47, (766) 1 --> (3903) 47:PEGB0, ND13, *, 
			10'd68 : rdata = 48'b000111110000000001100001101000000000000000000000;
			// PEs: 55, 55 -> 
			// srcs: (2279, 56)(3) 1, (3903) 47 --> (4687) 47:NM0, ALU, *, 
			10'd69 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 55, 55 -> 55
			// srcs: (2282, 70)(1551) -2, (4687) 47 --> (5471) -49:NW13, ALU, -, NW13
			10'd70 : rdata = 48'b000100100000110100111111111000000111010000000000;
			default : rdata = 48'b000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 56) begin
	always @(*) begin
		case(address)
			// PEs: 57 -> 24
			// srcs: (6, 0)(1642) 1 --> (1642) 1:PEGB1, pass, PUGB3
			10'd0 : rdata = 48'b110001110000001000000000000000000000000000001011;
			// PEs: 58 -> 24
			// srcs: (7, 1)(1644) -1 --> (1644) -1:PEGB2, pass, PUGB3
			10'd1 : rdata = 48'b110001110000010000000000000000000000000000001011;
			// PEs: 59 -> 24
			// srcs: (8, 2)(1645) -4 --> (1645) -4:PEGB3, pass, PUGB3
			10'd2 : rdata = 48'b110001110000011000000000000000000000000000001011;
			// PEs: 60 -> 24
			// srcs: (9, 3)(1647) 2 --> (1647) 2:PEGB4, pass, PUGB3
			10'd3 : rdata = 48'b110001110000100000000000000000000000000000001011;
			// PEs: 61 -> 24
			// srcs: (10, 4)(1648) -6 --> (1648) -6:PEGB5, pass, PUGB3
			10'd4 : rdata = 48'b110001110000101000000000000000000000000000001011;
			// PEs: 62 -> 24
			// srcs: (11, 5)(1650) 9 --> (1650) 9:PEGB6, pass, PUGB3
			10'd5 : rdata = 48'b110001110000110000000000000000000000000000001011;
			// PEs: 63 -> 24
			// srcs: (12, 6)(1651) -2 --> (1651) -2:PENB, pass, PUGB3
			10'd6 : rdata = 48'b110001101111111000000000000000000000000000001011;
			// PEs: 58 -> 0
			// srcs: (13, 16)(1724) 2 --> (1724) 2:PEGB2, pass, PUNB
			10'd7 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 59 -> 0
			// srcs: (14, 17)(1725) 6 --> (1725) 6:PEGB3, pass, PUNB
			10'd8 : rdata = 48'b110001110000011000000000000000000000001000000000;
			// PEs: 60 -> 0
			// srcs: (15, 18)(1727) 0 --> (1727) 0:PEGB4, pass, PUNB
			10'd9 : rdata = 48'b110001110000100000000000000000000000001000000000;
			// PEs: 61 -> 0
			// srcs: (16, 19)(1728) 6 --> (1728) 6:PEGB5, pass, PUNB
			10'd10 : rdata = 48'b110001110000101000000000000000000000001000000000;
			// PEs: 62 -> 0
			// srcs: (17, 20)(1730) 0 --> (1730) 0:PEGB6, pass, PUNB
			10'd11 : rdata = 48'b110001110000110000000000000000000000001000000000;
			// PEs: 63 -> 0
			// srcs: (18, 21)(1731) -2 --> (1731) -2:PENB, pass, PUNB
			10'd12 : rdata = 48'b110001101111111000000000000000000000001000000000;
			// PEs: 57 -> 0
			// srcs: (19, 31)(1804) -4 --> (1804) -4:PEGB1, pass, PUNB
			10'd13 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 48 -> 56
			// srcs: (20, 10)(1714) 9 --> (1714) 9:PUNB, pass, NI0
			10'd14 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 48 -> 58
			// srcs: (21, 11)(1715) -2 --> (1715) -2:PUNB, pass, PEGB2
			10'd15 : rdata = 48'b110001101111111100000000000000000000000010100000;
			// PEs: 48 -> 56
			// srcs: (22, 13)(1717) 0 --> (1717) 0:PUNB, pass, NI1
			10'd16 : rdata = 48'b110001101111111100000000000100001000000000000000;
			// PEs: 48 -> 59
			// srcs: (23, 14)(1718) 2 --> (1718) 2:PUNB, pass, PEGB3
			10'd17 : rdata = 48'b110001101111111100000000000000000000000010110000;
			// PEs: 58 -> 0
			// srcs: (24, 32)(1806) 4 --> (1806) 4:PEGB2, pass, PUNB
			10'd18 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 59 -> 0
			// srcs: (25, 33)(1807) 4 --> (1807) 4:PEGB3, pass, PUNB
			10'd19 : rdata = 48'b110001110000011000000000000000000000001000000000;
			// PEs: 60 -> 0
			// srcs: (26, 34)(1809) 3 --> (1809) 3:PEGB4, pass, PUNB
			10'd20 : rdata = 48'b110001110000100000000000000000000000001000000000;
			// PEs: 61 -> 0
			// srcs: (27, 35)(1810) 3 --> (1810) 3:PEGB5, pass, PUNB
			10'd21 : rdata = 48'b110001110000101000000000000000000000001000000000;
			// PEs: 62 -> 32
			// srcs: (28, 36)(1812) 3 --> (1812) 3:PEGB6, pass, PUGB4
			10'd22 : rdata = 48'b110001110000110000000000000000000000000000001100;
			// PEs: 63 -> 32
			// srcs: (29, 37)(1813) 2 --> (1813) 2:PENB, pass, PUGB4
			10'd23 : rdata = 48'b110001101111111000000000000000000000000000001100;
			// PEs: 56 -> 58
			// srcs: (30, 12)(1714) 9 --> (1714) 9:NI0, pass, PEGB2
			10'd24 : rdata = 48'b110001010000000000000000000000000000000010100000;
			// PEs: 48 -> 56
			// srcs: (31, 22)(1794) 0 --> (1794) 0:PUNB, pass, NI0
			10'd25 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 56 -> 59
			// srcs: (32, 15)(1717) 0 --> (1717) 0:NI1, pass, PEGB3
			10'd26 : rdata = 48'b110001010000000100000000000000000000000010110000;
			// PEs: 48 -> 60
			// srcs: (33, 23)(1795) -4 --> (1795) -4:PUNB, pass, PEGB4
			10'd27 : rdata = 48'b110001101111111100000000000000000000000011000000;
			// PEs: 48 -> 56
			// srcs: (34, 25)(1797) -4 --> (1797) -4:PUNB, pass, NI1
			10'd28 : rdata = 48'b110001101111111100000000000100001000000000000000;
			// PEs: 48 -> 61
			// srcs: (35, 26)(1798) -3 --> (1798) -3:PUNB, pass, PEGB5
			10'd29 : rdata = 48'b110001101111111100000000000000000000000011010000;
			// PEs: 48 -> 56
			// srcs: (36, 28)(1800) -2 --> (1800) -2:PUNB, pass, NI2
			10'd30 : rdata = 48'b110001101111111100000000000100010000000000000000;
			// PEs: 57 -> 48
			// srcs: (37, 44)(1884) -1 --> (1884) -1:PEGB1, pass, PUGB6
			10'd31 : rdata = 48'b110001110000001000000000000000000000000000001110;
			// PEs: 58 -> 48
			// srcs: (38, 45)(1886) -6 --> (1886) -6:PEGB2, pass, PUGB6
			10'd32 : rdata = 48'b110001110000010000000000000000000000000000001110;
			// PEs: 16 -> 56
			// srcs: (39, 7)(1678) -1 --> (1678) -1:PUGB2, pass, NI3
			10'd33 : rdata = 48'b110001110000010100000000000100011000000000000000;
			// PEs: 48 -> 62
			// srcs: (40, 29)(1801) 0 --> (1801) 0:PUNB, pass, PEGB6
			10'd34 : rdata = 48'b110001101111111100000000000000000000000011100000;
			// PEs: 59 -> 48
			// srcs: (41, 46)(1887) -2 --> (1887) -2:PEGB3, pass, PUGB6
			10'd35 : rdata = 48'b110001110000011000000000000000000000000000001110;
			// PEs: 16 -> 57
			// srcs: (42, 8)(1679) -4 --> (1679) -4:PUGB2, pass, PENB
			10'd36 : rdata = 48'b110001110000010100000000000000000000000100000000;
			// PEs: 56 -> 60
			// srcs: (43, 24)(1794) 0 --> (1794) 0:NI0, pass, PEGB4
			10'd37 : rdata = 48'b110001010000000000000000000000000000000011000000;
			// PEs: 56 -> 61
			// srcs: (44, 27)(1797) -4 --> (1797) -4:NI1, pass, PEGB5
			10'd38 : rdata = 48'b110001010000000100000000000000000000000011010000;
			// PEs: 60 -> 0
			// srcs: (45, 47)(1889) 0 --> (1889) 0:PEGB4, pass, PUNB
			10'd39 : rdata = 48'b110001110000100000000000000000000000001000000000;
			// PEs: 48 -> 56
			// srcs: (46, 38)(1874) -2 --> (1874) -2:PUNB, pass, NI0
			10'd40 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 48 -> 63
			// srcs: (47, 39)(1875) 0 --> (1875) 0:PUNB, pass, PEGB7
			10'd41 : rdata = 48'b110001101111111100000000000000000000000011110000;
			// PEs: 56 -> 57
			// srcs: (48, 9)(1678) -1 --> (1678) -1:NI3, pass, PENB
			10'd42 : rdata = 48'b110001010000001100000000000000000000000100000000;
			// PEs: 56 -> 62
			// srcs: (49, 30)(1800) -2 --> (1800) -2:NI2, pass, PEGB6
			10'd43 : rdata = 48'b110001010000001000000000000000000000000011100000;
			// PEs: 61 -> 0
			// srcs: (50, 48)(1890) -2 --> (1890) -2:PEGB5, pass, PUNB
			10'd44 : rdata = 48'b110001110000101000000000000000000000001000000000;
			// PEs: 62 -> 0
			// srcs: (51, 49)(1892) 2 --> (1892) 2:PEGB6, pass, PUNB
			10'd45 : rdata = 48'b110001110000110000000000000000000000001000000000;
			// PEs: 48 -> 56
			// srcs: (52, 41)(1880) -1 --> (1880) -1:PUNB, pass, NI1
			10'd46 : rdata = 48'b110001101111111100000000000100001000000000000000;
			// PEs: 48 -> 58
			// srcs: (53, 42)(1881) 1 --> (1881) 1:PUNB, pass, PEGB2
			10'd47 : rdata = 48'b110001101111111100000000000000000000000010100000;
			// PEs: 63 -> 0
			// srcs: (54, 50)(1893) 0 --> (1893) 0:PENB, pass, PUNB
			10'd48 : rdata = 48'b110001101111111000000000000000000000001000000000;
			// PEs: 60 -> 0
			// srcs: (55, 60)(1969) -6 --> (1969) -6:PEGB4, pass, PUNB
			10'd49 : rdata = 48'b110001110000100000000000000000000000001000000000;
			// PEs: 56 -> 63
			// srcs: (56, 40)(1874) -2 --> (1874) -2:NI0, pass, PEGB7
			10'd50 : rdata = 48'b110001010000000000000000000000000000000011110000;
			// PEs: 61 -> 0
			// srcs: (57, 61)(1970) 2 --> (1970) 2:PEGB5, pass, PUNB
			10'd51 : rdata = 48'b110001110000101000000000000000000000001000000000;
			// PEs: 62 -> 0
			// srcs: (58, 62)(1972) -2 --> (1972) -2:PEGB6, pass, PUNB
			10'd52 : rdata = 48'b110001110000110000000000000000000000001000000000;
			// PEs: 63 -> 0
			// srcs: (59, 63)(1973) -6 --> (1973) -6:PENB, pass, PUNB
			10'd53 : rdata = 48'b110001101111111000000000000000000000001000000000;
			// PEs: 48 -> 56
			// srcs: (60, 51)(1956) -2 --> (1956) -2:PUNB, pass, NI0
			10'd54 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 48 -> 57
			// srcs: (61, 52)(1957) 0 --> (1957) 0:PUNB, pass, PENB
			10'd55 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 56 -> 58
			// srcs: (62, 43)(1880) -1 --> (1880) -1:NI1, pass, PEGB2
			10'd56 : rdata = 48'b110001010000000100000000000000000000000010100000;
			// PEs: 58 -> 0
			// srcs: (63, 74)(2048) 1 --> (2048) 1:PEGB2, pass, PUNB
			10'd57 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 59 -> 0
			// srcs: (64, 75)(2049) 0 --> (2049) 0:PEGB3, pass, PUNB
			10'd58 : rdata = 48'b110001110000011000000000000000000000001000000000;
			// PEs: 60 -> 0
			// srcs: (65, 76)(2051) -4 --> (2051) -4:PEGB4, pass, PUNB
			10'd59 : rdata = 48'b110001110000100000000000000000000000001000000000;
			// PEs: 61 -> 0
			// srcs: (66, 77)(2052) 0 --> (2052) 0:PEGB5, pass, PUNB
			10'd60 : rdata = 48'b110001110000101000000000000000000000001000000000;
			// PEs: 56 -> 57
			// srcs: (67, 53)(1956) -2 --> (1956) -2:NI0, pass, PENB
			10'd61 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 48 -> 56
			// srcs: (68, 54)(1959) 0 --> (1959) 0:PUNB, pass, NI0
			10'd62 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 48 -> 57
			// srcs: (69, 55)(1960) 0 --> (1960) 0:PUNB, pass, PENB
			10'd63 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 62 -> 0
			// srcs: (70, 78)(2054) -6 --> (2054) -6:PEGB6, pass, PUNB
			10'd64 : rdata = 48'b110001110000110000000000000000000000001000000000;
			// PEs: 63 -> 0
			// srcs: (71, 79)(2055) 0 --> (2055) 0:PENB, pass, PUNB
			10'd65 : rdata = 48'b110001101111111000000000000000000000001000000000;
			// PEs: 58 -> 0
			// srcs: (72, 90)(2128) -4 --> (2128) -4:PEGB2, pass, PUNB
			10'd66 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 59 -> 0
			// srcs: (73, 91)(2129) 6 --> (2129) 6:PEGB3, pass, PUNB
			10'd67 : rdata = 48'b110001110000011000000000000000000000001000000000;
			// PEs: 60 -> 0
			// srcs: (74, 92)(2131) 2 --> (2131) 2:PEGB4, pass, PUNB
			10'd68 : rdata = 48'b110001110000100000000000000000000000001000000000;
			// PEs: 56 -> 57
			// srcs: (75, 56)(1959) 0 --> (1959) 0:NI0, pass, PENB
			10'd69 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 48 -> 56
			// srcs: (76, 57)(1962) 6 --> (1962) 6:PUNB, pass, NI0
			10'd70 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 48 -> 57
			// srcs: (77, 58)(1963) 0 --> (1963) 0:PUNB, pass, PENB
			10'd71 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 61 -> 0
			// srcs: (78, 93)(2132) -2 --> (2132) -2:PEGB5, pass, PUNB
			10'd72 : rdata = 48'b110001110000101000000000000000000000001000000000;
			// PEs: 62 -> 0
			// srcs: (79, 94)(2134) 2 --> (2134) 2:PEGB6, pass, PUNB
			10'd73 : rdata = 48'b110001110000110000000000000000000000001000000000;
			// PEs: 63 -> 0
			// srcs: (80, 95)(2135) -3 --> (2135) -3:PENB, pass, PUNB
			10'd74 : rdata = 48'b110001101111111000000000000000000000001000000000;
			// PEs: 62 -> 0
			// srcs: (81, 106)(2214) -3 --> (2214) -3:PEGB6, pass, PUNB
			10'd75 : rdata = 48'b110001110000110000000000000000000000001000000000;
			// PEs: 63 -> 0
			// srcs: (82, 107)(2215) 2 --> (2215) 2:PENB, pass, PUNB
			10'd76 : rdata = 48'b110001101111111000000000000000000000001000000000;
			// PEs: 56 -> 57
			// srcs: (83, 59)(1962) 6 --> (1962) 6:NI0, pass, PENB
			10'd77 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 48 -> 56
			// srcs: (84, 64)(2036) 0 --> (2036) 0:PUNB, pass, NI0
			10'd78 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 48 -> 57
			// srcs: (85, 65)(2037) -1 --> (2037) -1:PUNB, pass, PENB
			10'd79 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 32 -> 56
			// srcs: (86, 112)(1622) -6 --> (1622) -6:PUGB4, pass, NI1
			10'd80 : rdata = 48'b110001110000100100000000000100001000000000000000;
			// PEs: 57 -> 24
			// srcs: (87, 130)(1606) 6 --> (1606) 6:PEGB1, pass, PUGB3
			10'd81 : rdata = 48'b110001110000001000000000000000000000000000001011;
			// PEs: 58 -> 32
			// srcs: (88, 131)(1609) 6 --> (1609) 6:PEGB2, pass, PUGB4
			10'd82 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 57 -> 32
			// srcs: (89, 141)(2460) -5 --> (2460) -5:PEGB1, pass, PUGB4
			10'd83 : rdata = 48'b110001110000001000000000000000000000000000001100;
			// PEs: 59 -> 8
			// srcs: (90, 149)(2496) 2 --> (2496) 2:PEGB3, pass, PUGB1
			10'd84 : rdata = 48'b110001110000011000000000000000000000000000001001;
			// PEs: 56 -> 57
			// srcs: (91, 66)(2036) 0 --> (2036) 0:NI0, pass, PENB
			10'd85 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 48 -> 56
			// srcs: (92, 67)(2039) 3 --> (2039) 3:PUNB, pass, NI0
			10'd86 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 48 -> 57
			// srcs: (93, 68)(2040) 0 --> (2040) 0:PUNB, pass, PENB
			10'd87 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 57 -> 0
			// srcs: (94, 118)(1723) 0 --> (1723) 0:PEGB1, pass, PUNB
			10'd88 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 58 -> 40
			// srcs: (95, 155)(1793) -1 --> (1793) -1:PEGB2, pass, PUGB5
			10'd89 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 58 -> 32
			// srcs: (96, 168)(2661) 0 --> (2661) 0:PEGB2, pass, PUGB4
			10'd90 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 56 -> 57
			// srcs: (99, 69)(2039) 3 --> (2039) 3:NI0, pass, PENB
			10'd91 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 48 -> 56
			// srcs: (100, 70)(2042) 2 --> (2042) 2:PUNB, pass, NI0
			10'd92 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 48 -> 57
			// srcs: (101, 71)(2043) 3 --> (2043) 3:PUNB, pass, PENB
			10'd93 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 48 -> 59
			// srcs: (102, 73)(2045) -2 --> (2045) -2:PUNB, pass, PEGB3
			10'd94 : rdata = 48'b110001101111111100000000000000000000000010110000;
			// PEs: 58 -> 0
			// srcs: (103, 120)(1967) 0 --> (1967) 0:PEGB2, pass, PUNB
			10'd95 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 59 -> 24
			// srcs: (104, 178)(1980) 0 --> (1980) 0:PEGB3, pass, PUGB3
			10'd96 : rdata = 48'b110001110000011000000000000000000000000000001011;
			// PEs: 58 -> 40
			// srcs: (105, 198)(2157) 4 --> (2157) 4:PEGB2, pass, PUGB5
			10'd97 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 56 -> 57
			// srcs: (107, 72)(2042) 2 --> (2042) 2:NI0, pass, PENB
			10'd98 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 48 -> 56
			// srcs: (108, 80)(2116) -2 --> (2116) -2:PUNB, pass, NI0
			10'd99 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 48 -> 57
			// srcs: (109, 81)(2117) 2 --> (2117) 2:PUNB, pass, PENB
			10'd100 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 59 -> 0
			// srcs: (111, 121)(1968) 0 --> (1968) 0:PEGB3, pass, PUNB
			10'd101 : rdata = 48'b110001110000011000000000000000000000001000000000;
			// PEs: 56 -> 57
			// srcs: (115, 82)(2116) -2 --> (2116) -2:NI0, pass, PENB
			10'd102 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 48 -> 56
			// srcs: (116, 83)(2119) 4 --> (2119) 4:PUNB, pass, NI0
			10'd103 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 48 -> 57
			// srcs: (117, 84)(2120) 9 --> (2120) 9:PUNB, pass, PENB
			10'd104 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 58 -> 0
			// srcs: (119, 122)(2210) -1 --> (2210) -1:PEGB2, pass, PUNB
			10'd105 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 56 -> 57
			// srcs: (123, 85)(2119) 4 --> (2119) 4:NI0, pass, PENB
			10'd106 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 48 -> 56
			// srcs: (124, 86)(2122) 0 --> (2122) 0:PUNB, pass, NI0
			10'd107 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 48 -> 57
			// srcs: (125, 87)(2123) 6 --> (2123) 6:PUNB, pass, PENB
			10'd108 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 48 -> 60
			// srcs: (126, 89)(2125) -2 --> (2125) -2:PUNB, pass, PEGB4
			10'd109 : rdata = 48'b110001101111111100000000000000000000000011000000;
			// PEs: 59 -> 0
			// srcs: (127, 123)(2211) -1 --> (2211) -1:PEGB3, pass, PUNB
			10'd110 : rdata = 48'b110001110000011000000000000000000000001000000000;
			// PEs: 60 -> 0
			// srcs: (128, 124)(2212) 0 --> (2212) 0:PEGB4, pass, PUNB
			10'd111 : rdata = 48'b110001110000100000000000000000000000001000000000;
			// PEs: 61 -> 0
			// srcs: (129, 125)(2213) 0 --> (2213) 0:PEGB5, pass, PUNB
			10'd112 : rdata = 48'b110001110000101000000000000000000000001000000000;
			// PEs: 61 -> 16
			// srcs: (130, 134)(1618) -6 --> (1618) -6:PEGB5, pass, PUGB2
			10'd113 : rdata = 48'b110001110000101000000000000000000000000000001010;
			// PEs: 56 -> 57
			// srcs: (131, 88)(2122) 0 --> (2122) 0:NI0, pass, PENB
			10'd114 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 48 -> 56
			// srcs: (132, 96)(2198) 0 --> (2198) 0:PUNB, pass, NI0
			10'd115 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 48 -> 57
			// srcs: (133, 97)(2199) -4 --> (2199) -4:PUNB, pass, PENB
			10'd116 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 63 -> 16
			// srcs: (134, 137)(1628) 2 --> (1628) 2:PENB, pass, PUGB2
			10'd117 : rdata = 48'b110001101111111000000000000000000000000000001010;
			// PEs: 63 -> 16
			// srcs: (135, 167)(2655) -2 --> (2655) -2:PENB, pass, PUGB2
			10'd118 : rdata = 48'b110001101111111000000000000000000000000000001010;
			// PEs: 60 -> 32
			// srcs: (136, 200)(2167) -1 --> (2167) -1:PEGB4, pass, PUGB4
			10'd119 : rdata = 48'b110001110000100000000000000000000000000000001100;
			// PEs: 59 -> 0
			// srcs: (137, 132)(1612) 0 --> (1612) 0:PEGB3, pass, PUNB
			10'd120 : rdata = 48'b110001110000011000000000000000000000001000000000;
			// PEs: 56 -> 57
			// srcs: (139, 98)(2198) 0 --> (2198) 0:NI0, pass, PENB
			10'd121 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 48 -> 56
			// srcs: (140, 99)(2201) 2 --> (2201) 2:PUNB, pass, NI0
			10'd122 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 48 -> 57
			// srcs: (141, 100)(2202) 2 --> (2202) 2:PUNB, pass, PENB
			10'd123 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 63 -> 24
			// srcs: (142, 182)(1992) 4 --> (1992) 4:PENB, pass, PUGB3
			10'd124 : rdata = 48'b110001101111111000000000000000000000000000001011;
			// PEs: 57 -> 24
			// srcs: (143, 187)(2820) 3 --> (2820) 3:PEGB1, pass, PUGB3
			10'd125 : rdata = 48'b110001110000001000000000000000000000000000001011;
			// PEs: 57 -> 8
			// srcs: (144, 195)(2901) 6 --> (2901) 6:PEGB1, pass, PUGB1
			10'd126 : rdata = 48'b110001110000001000000000000000000000000000001001;
			// PEs: 58 -> 0
			// srcs: (145, 148)(2494) 7 --> (2494) 7:PEGB2, pass, PUNB
			10'd127 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 63 -> 32
			// srcs: (146, 203)(2176) 2 --> (2176) 2:PENB, pass, PUGB4
			10'd128 : rdata = 48'b110001101111111000000000000000000000000000001100;
			// PEs: 56 -> 57
			// srcs: (147, 101)(2201) 2 --> (2201) 2:NI0, pass, PENB
			10'd129 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 48 -> 56
			// srcs: (148, 102)(2204) -3 --> (2204) -3:PUNB, pass, NI0
			10'd130 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 48 -> 57
			// srcs: (149, 103)(2205) 2 --> (2205) 2:PUNB, pass, PENB
			10'd131 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 57 -> 8
			// srcs: (150, 210)(2978) -4 --> (2978) -4:PEGB1, pass, PUGB1
			10'd132 : rdata = 48'b110001110000001000000000000000000000000000001001;
			// PEs: 56 -> 57
			// srcs: (155, 104)(2204) -3 --> (2204) -3:NI0, pass, PENB
			10'd133 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 48 -> 57
			// srcs: (156, 105)(2207) -4 --> (2207) -4:PUNB, pass, PENB
			10'd134 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 48 -> 57
			// srcs: (157, 108)(2287) 0 --> (2287) 0:PUNB, pass, PENB
			10'd135 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 58 -> 32
			// srcs: (158, 220)(3075) 4 --> (3075) 4:PEGB2, pass, PUGB4
			10'd136 : rdata = 48'b110001110000010000000000000000000000000000001100;
			// PEs: 57 -> 24
			// srcs: (162, 212)(2983) -1 --> (2983) -1:PEGB1, pass, PUGB3
			10'd137 : rdata = 48'b110001110000001000000000000000000000000000001011;
			// PEs: 60 -> 24
			// srcs: (163, 230)(2347) 2 --> (2347) 2:PEGB4, pass, PUGB3
			10'd138 : rdata = 48'b110001110000100000000000000000000000000000001011;
			// PEs: 40 -> 62
			// srcs: (195, 113)(1623) 0 --> (1623) 0:PUGB5, pass, PEGB6
			10'd139 : rdata = 48'b110001110000101100000000000000000000000011100000;
			// PEs: 56 -> 62
			// srcs: (204, 114)(1622) -6 --> (1622) -6:NI1, pass, PEGB6
			10'd140 : rdata = 48'b110001010000000100000000000000000000000011100000;
			// PEs: 48 -> 56
			// srcs: (213, 115)(1720) 6 --> (1720) 6:PUNB, pass, NI0
			10'd141 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 0 -> 56
			// srcs: (222, 109)(1575) 0 --> (1575) 0:PUGB0, pass, NI1
			10'd142 : rdata = 48'b110001110000000100000000000100001000000000000000;
			// PEs: 48 -> 59
			// srcs: (229, 116)(1721) 1 --> (1721) 1:PUNB, pass, PEGB3
			10'd143 : rdata = 48'b110001101111111100000000000000000000000010110000;
			// PEs: 56 -> 59
			// srcs: (238, 117)(1720) 6 --> (1720) 6:NI0, pass, PEGB3
			10'd144 : rdata = 48'b110001010000000000000000000000000000000010110000;
			// PEs: 48 -> 60
			// srcs: (239, 119)(1965) -3 --> (1965) -3:PUNB, pass, PEGB4
			10'd145 : rdata = 48'b110001101111111100000000000000000000000011000000;
			// PEs: 0 -> 63
			// srcs: (246, 110)(1576) 0 --> (1576) 0:PUGB0, pass, PEGB7
			10'd146 : rdata = 48'b110001110000000100000000000000000000000011110000;
			// PEs: 0 -> 56
			// srcs: (247, 127)(2374) 6 --> (2374) 6:PUGB0, pass, NI0
			10'd147 : rdata = 48'b110001110000000100000000000100000000000000000000;
			// PEs: 48 -> 57
			// srcs: (248, 128)(1594) -1 --> (1594) -1:PUNB, pass, PENB
			10'd148 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 59 -> 0
			// srcs: (249, 150)(2502) 7 --> (2502) 7:PEGB3, pass, PUNB
			10'd149 : rdata = 48'b110001110000011000000000000000000000001000000000;
			// PEs: 56 -> 57
			// srcs: (254, 129)(2374) 6 --> (2374) 6:NI0, pass, PENB
			10'd150 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 56 -> 63
			// srcs: (255, 111)(1575) 0 --> (1575) 0:NI1, pass, PEGB7
			10'd151 : rdata = 48'b110001010000000100000000000000000000000011110000;
			// PEs: 8 -> 57
			// srcs: (256, 133)(2394) 6 --> (2394) 6:PUGB1, pass, PENB
			10'd152 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 57
			// srcs: (257, 136)(2406) 4 --> (2406) 4:PUGB1, pass, PENB
			10'd153 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 40 -> 56
			// srcs: (258, 138)(2445) -1 --> (2445) -1:PUGB5, pass, NI0
			10'd154 : rdata = 48'b110001110000101100000000000100000000000000000000;
			// PEs: 63 -> 48
			// srcs: (262, 126)(2358) 0 --> (2358) 0:PENB, pass, PUGB6
			10'd155 : rdata = 48'b110001101111111000000000000000000000000000001110;
			// PEs: 62 -> 48
			// srcs: (263, 135)(1621) 2 --> (1621) 2:PEGB6, pass, PUGB6
			10'd156 : rdata = 48'b110001110000110000000000000000000000000000001110;
			// PEs: 62 -> 0
			// srcs: (264, 156)(1805) 0 --> (1805) 0:PEGB6, pass, PUNB
			10'd157 : rdata = 48'b110001110000110000000000000000000000001000000000;
			// PEs: 62 -> 48
			// srcs: (265, 181)(1989) 4 --> (1989) 4:PEGB6, pass, PUGB6
			10'd158 : rdata = 48'b110001110000110000000000000000000000000000001110;
			// PEs: 62 -> 8
			// srcs: (266, 219)(3071) -1 --> (3071) -1:PEGB6, pass, PUGB1
			10'd159 : rdata = 48'b110001110000110000000000000000000000000000001001;
			// PEs: 57 -> 24
			// srcs: (267, 236)(2407) -2 --> (2407) -2:PEGB1, pass, PUGB3
			10'd160 : rdata = 48'b110001110000001000000000000000000000000000001011;
			// PEs: 63 -> 0
			// srcs: (269, 157)(1808) 0 --> (1808) 0:PENB, pass, PUNB
			10'd161 : rdata = 48'b110001101111111000000000000000000000001000000000;
			// PEs: 60 -> 0
			// srcs: (270, 175)(2748) -1 --> (2748) -1:PEGB4, pass, PUNB
			10'd162 : rdata = 48'b110001110000100000000000000000000000001000000000;
			// PEs: 59 -> 48
			// srcs: (273, 199)(2160) 4 --> (2160) 4:PEGB3, pass, PUGB6
			10'd163 : rdata = 48'b110001110000011000000000000000000000000000001110;
			// PEs: 57 -> 8
			// srcs: (274, 227)(2338) 0 --> (2338) 0:PEGB1, pass, PUGB1
			10'd164 : rdata = 48'b110001110000001000000000000000000000000000001001;
			// PEs: 57 -> 0
			// srcs: (278, 176)(1974) 6 --> (1974) 6:PEGB1, pass, PUNB
			10'd165 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 61 -> 0
			// srcs: (279, 180)(1986) 0 --> (1986) 0:PEGB5, pass, PUNB
			10'd166 : rdata = 48'b110001110000101000000000000000000000001000000000;
			// PEs: 61 -> 40
			// srcs: (280, 201)(2170) -6 --> (2170) -6:PEGB5, pass, PUGB5
			10'd167 : rdata = 48'b110001110000101000000000000000000000000000001101;
			// PEs: 61 -> 48
			// srcs: (281, 218)(3069) 6 --> (3069) 6:PEGB5, pass, PUGB6
			10'd168 : rdata = 48'b110001110000101000000000000000000000000000001110;
			// PEs: 62 -> 8
			// srcs: (282, 232)(2353) 1 --> (2353) 1:PEGB6, pass, PUGB1
			10'd169 : rdata = 48'b110001110000110000000000000000000000000000001001;
			// PEs: 57 -> 0
			// srcs: (287, 186)(2815) -1 --> (2815) -1:PEGB1, pass, PUNB
			10'd170 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 57 -> 40
			// srcs: (288, 211)(2980) 4 --> (2980) 4:PEGB1, pass, PUGB5
			10'd171 : rdata = 48'b110001110000001000000000000000000000000000001101;
			// PEs: 61 -> 32
			// srcs: (289, 231)(2350) -3 --> (2350) -3:PEGB5, pass, PUGB4
			10'd172 : rdata = 48'b110001110000101000000000000000000000000000001100;
			// PEs: 57 -> 0
			// srcs: (296, 213)(2985) -2 --> (2985) -2:PEGB1, pass, PUNB
			10'd173 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 58 -> 40
			// srcs: (297, 228)(2341) -4 --> (2341) -4:PEGB2, pass, PUGB5
			10'd174 : rdata = 48'b110001110000010000000000000000000000000000001101;
			// PEs: 63 -> 40
			// srcs: (302, 233)(2356) 0 --> (2356) 0:PENB, pass, PUGB5
			10'd175 : rdata = 48'b110001101111111000000000000000000000000000001101;
			// PEs: 59 -> 0
			// srcs: (305, 229)(2344) 0 --> (2344) 0:PEGB3, pass, PUNB
			10'd176 : rdata = 48'b110001110000011000000000000000000000001000000000;
			// PEs: 57 -> 0
			// srcs: (313, 235)(2395) 6 --> (2395) 6:PEGB1, pass, PUNB
			10'd177 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 8 -> 57
			// srcs: (461, 139)(1667) 4 --> (1667) 4:PUGB1, pass, PENB
			10'd178 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 56 -> 57
			// srcs: (467, 140)(2445) -1 --> (2445) -1:NI0, pass, PENB
			10'd179 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 32 -> 56
			// srcs: (468, 142)(2468) -5 --> (2468) -5:PUGB4, pass, NI0
			10'd180 : rdata = 48'b110001110000100100000000000100000000000000000000;
			// PEs: 16 -> 57
			// srcs: (469, 143)(1689) 0 --> (1689) 0:PUGB2, pass, PENB
			10'd181 : rdata = 48'b110001110000010100000000000000000000000100000000;
			// PEs: 56 -> 57
			// srcs: (475, 144)(2468) -5 --> (2468) -5:NI0, pass, PENB
			10'd182 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 48 -> 56
			// srcs: (476, 145)(2491) -6 --> (2491) -6:PUNB, pass, NI0
			10'd183 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 24 -> 57
			// srcs: (477, 146)(1713) -2 --> (1713) -2:PUGB3, pass, PENB
			10'd184 : rdata = 48'b110001110000011100000000000000000000000100000000;
			// PEs: 57 -> 48
			// srcs: (482, 241)(2469) -5 --> (2469) -5:PEGB1, pass, PUGB6
			10'd185 : rdata = 48'b110001110000001000000000000000000000000000001110;
			// PEs: 56 -> 57
			// srcs: (483, 147)(2491) -6 --> (2491) -6:NI0, pass, PENB
			10'd186 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 0 -> 56
			// srcs: (484, 151)(2521) 4 --> (2521) 4:PUGB0, pass, NI0
			10'd187 : rdata = 48'b110001110000000100000000000100000000000000000000;
			// PEs: 40 -> 57
			// srcs: (485, 152)(1744) 1 --> (1744) 1:PUGB5, pass, PENB
			10'd188 : rdata = 48'b110001110000101100000000000000000000000100000000;
			// PEs: 57 -> 24
			// srcs: (490, 242)(2492) -8 --> (2492) -8:PEGB1, pass, PUGB3
			10'd189 : rdata = 48'b110001110000001000000000000000000000000000001011;
			// PEs: 56 -> 57
			// srcs: (491, 153)(2521) 4 --> (2521) 4:NI0, pass, PENB
			10'd190 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 16 -> 57
			// srcs: (492, 154)(2569) 7 --> (2569) 7:PUGB2, pass, PENB
			10'd191 : rdata = 48'b110001110000010100000000000000000000000100000000;
			// PEs: 16 -> 56
			// srcs: (493, 158)(2603) 0 --> (2603) 0:PUGB2, pass, NI0
			10'd192 : rdata = 48'b110001110000010100000000000100000000000000000000;
			// PEs: 0 -> 57
			// srcs: (494, 159)(1824) 3 --> (1824) 3:PUGB0, pass, PENB
			10'd193 : rdata = 48'b110001110000000100000000000000000000000100000000;
			// PEs: 57 -> 0
			// srcs: (498, 246)(2522) 5 --> (2522) 5:PEGB1, pass, PUNB
			10'd194 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 56 -> 57
			// srcs: (500, 160)(2603) 0 --> (2603) 0:NI0, pass, PENB
			10'd195 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 24 -> 56
			// srcs: (501, 161)(2619) -2 --> (2619) -2:PUGB3, pass, NI0
			10'd196 : rdata = 48'b110001110000011100000000000100000000000000000000;
			// PEs: 8 -> 57
			// srcs: (502, 162)(1842) 3 --> (1842) 3:PUGB1, pass, PENB
			10'd197 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 62 -> 0
			// srcs: (506, 248)(2582) 1 --> (2582) 1:PEGB6, pass, PUNB
			10'd198 : rdata = 48'b110001110000110000000000000000000000001000000000;
			// PEs: 57 -> 24
			// srcs: (507, 249)(2604) 3 --> (2604) 3:PEGB1, pass, PUGB3
			10'd199 : rdata = 48'b110001110000001000000000000000000000000000001011;
			// PEs: 56 -> 57
			// srcs: (508, 163)(2619) -2 --> (2619) -2:NI0, pass, PENB
			10'd200 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 48 -> 56
			// srcs: (509, 164)(2642) -2 --> (2642) -2:PUNB, pass, NI0
			10'd201 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 16 -> 57
			// srcs: (510, 165)(1866) -3 --> (1866) -3:PUGB2, pass, PENB
			10'd202 : rdata = 48'b110001110000010100000000000000000000000100000000;
			// PEs: 48 -> 61
			// srcs: (511, 172)(1958) 4 --> (1958) 4:PUNB, pass, PEGB5
			10'd203 : rdata = 48'b110001101111111100000000000000000000000011010000;
			// PEs: 48 -> 63
			// srcs: (512, 173)(1961) 3 --> (1961) 3:PUNB, pass, PEGB7
			10'd204 : rdata = 48'b110001101111111100000000000000000000000011110000;
			// PEs: 48 -> 62
			// srcs: (513, 174)(1964) 9 --> (1964) 9:PUNB, pass, PEGB6
			10'd205 : rdata = 48'b110001101111111100000000000000000000000011100000;
			// PEs: 57 -> 48
			// srcs: (515, 253)(2620) 1 --> (2620) 1:PEGB1, pass, PUGB6
			10'd206 : rdata = 48'b110001110000001000000000000000000000000000001110;
			// PEs: 56 -> 57
			// srcs: (516, 166)(2642) -2 --> (2642) -2:NI0, pass, PENB
			10'd207 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 0 -> 56
			// srcs: (517, 169)(2673) 2 --> (2673) 2:PUGB0, pass, NI0
			10'd208 : rdata = 48'b110001110000000100000000000100000000000000000000;
			// PEs: 24 -> 57
			// srcs: (518, 170)(1894) 4 --> (1894) 4:PUGB3, pass, PENB
			10'd209 : rdata = 48'b110001110000011100000000000000000000000100000000;
			// PEs: 57 -> 40
			// srcs: (523, 254)(2643) -5 --> (2643) -5:PEGB1, pass, PUGB5
			10'd210 : rdata = 48'b110001110000001000000000000000000000000000001101;
			// PEs: 56 -> 57
			// srcs: (524, 171)(2673) 2 --> (2673) 2:NI0, pass, PENB
			10'd211 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 8 -> 57
			// srcs: (525, 177)(2756) -5 --> (2756) -5:PUGB1, pass, PENB
			10'd212 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 57
			// srcs: (526, 179)(2762) -6 --> (2762) -6:PUGB1, pass, PENB
			10'd213 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 24 -> 56
			// srcs: (527, 183)(2779) 8 --> (2779) 8:PUGB3, pass, NI0
			10'd214 : rdata = 48'b110001110000011100000000000100000000000000000000;
			// PEs: 0 -> 57
			// srcs: (528, 184)(2001) 0 --> (2001) 0:PUGB0, pass, PENB
			10'd215 : rdata = 48'b110001110000000100000000000000000000000100000000;
			// PEs: 57 -> 0
			// srcs: (532, 257)(2757) -5 --> (2757) -5:PEGB1, pass, PUNB
			10'd216 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 57 -> 8
			// srcs: (533, 258)(2763) -4 --> (2763) -4:PEGB1, pass, PUGB1
			10'd217 : rdata = 48'b110001110000001000000000000000000000000000001001;
			// PEs: 56 -> 57
			// srcs: (534, 185)(2779) 8 --> (2779) 8:NI0, pass, PENB
			10'd218 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 16 -> 57
			// srcs: (535, 188)(2044) 0 --> (2044) 0:PUGB2, pass, PENB
			10'd219 : rdata = 48'b110001110000010100000000000000000000000100000000;
			// PEs: 16 -> 57
			// srcs: (536, 189)(2047) -4 --> (2047) -4:PUGB2, pass, PENB
			10'd220 : rdata = 48'b110001110000010100000000000000000000000100000000;
			// PEs: 0 -> 56
			// srcs: (537, 190)(2833) -6 --> (2833) -6:PUGB0, pass, NI0
			10'd221 : rdata = 48'b110001110000000100000000000100000000000000000000;
			// PEs: 16 -> 57
			// srcs: (538, 191)(2056) 0 --> (2056) 0:PUGB2, pass, PENB
			10'd222 : rdata = 48'b110001110000010100000000000000000000000100000000;
			// PEs: 57 -> 24
			// srcs: (541, 259)(2780) 8 --> (2780) 8:PEGB1, pass, PUGB3
			10'd223 : rdata = 48'b110001110000001000000000000000000000000000001011;
			// PEs: 57 -> 32
			// srcs: (542, 263)(2823) 5 --> (2823) 5:PEGB1, pass, PUGB4
			10'd224 : rdata = 48'b110001110000001000000000000000000000000000001100;
			// PEs: 56 -> 57
			// srcs: (544, 192)(2833) -6 --> (2833) -6:NI0, pass, PENB
			10'd225 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 40 -> 57
			// srcs: (545, 193)(2118) -2 --> (2118) -2:PUGB5, pass, PENB
			10'd226 : rdata = 48'b110001110000101100000000000000000000000100000000;
			// PEs: 40 -> 57
			// srcs: (546, 194)(2121) 0 --> (2121) 0:PUGB5, pass, PENB
			10'd227 : rdata = 48'b110001110000101100000000000000000000000100000000;
			// PEs: 40 -> 57
			// srcs: (547, 196)(2127) -2 --> (2127) -2:PUGB5, pass, PENB
			10'd228 : rdata = 48'b110001110000101100000000000000000000000100000000;
			// PEs: 16 -> 57
			// srcs: (548, 197)(2930) 4 --> (2930) 4:PUGB2, pass, PENB
			10'd229 : rdata = 48'b110001110000010100000000000000000000000100000000;
			// PEs: 32 -> 57
			// srcs: (549, 202)(2951) 4 --> (2951) 4:PUGB4, pass, PENB
			10'd230 : rdata = 48'b110001110000100100000000000000000000000100000000;
			// PEs: 40 -> 56
			// srcs: (550, 204)(2962) -5 --> (2962) -5:PUGB5, pass, NI0
			10'd231 : rdata = 48'b110001110000101100000000000100000000000000000000;
			// PEs: 0 -> 57
			// srcs: (551, 205)(2185) -2 --> (2185) -2:PUGB0, pass, PENB
			10'd232 : rdata = 48'b110001110000000100000000000000000000000100000000;
			// PEs: 57 -> 0
			// srcs: (552, 265)(2834) -6 --> (2834) -6:PEGB1, pass, PUNB
			10'd233 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 57 -> 8
			// srcs: (553, 267)(2900) 13 --> (2900) 13:PEGB1, pass, PUGB1
			10'd234 : rdata = 48'b110001110000001000000000000000000000000000001001;
			// PEs: 57 -> 16
			// srcs: (554, 268)(2906) 0 --> (2906) 0:PEGB1, pass, PUGB2
			10'd235 : rdata = 48'b110001110000001000000000000000000000000000001010;
			// PEs: 56 -> 57
			// srcs: (562, 206)(2962) -5 --> (2962) -5:NI0, pass, PENB
			10'd236 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 40 -> 56
			// srcs: (563, 207)(2967) 5 --> (2967) 5:PUGB5, pass, NI0
			10'd237 : rdata = 48'b110001110000101100000000000100000000000000000000;
			// PEs: 0 -> 57
			// srcs: (564, 208)(2188) 0 --> (2188) 0:PUGB0, pass, PENB
			10'd238 : rdata = 48'b110001110000000100000000000000000000000100000000;
			// PEs: 57 -> 0
			// srcs: (565, 270)(2952) 4 --> (2952) 4:PEGB1, pass, PUNB
			10'd239 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 57 -> 24
			// srcs: (569, 271)(2963) -7 --> (2963) -7:PEGB1, pass, PUGB3
			10'd240 : rdata = 48'b110001110000001000000000000000000000000000001011;
			// PEs: 56 -> 57
			// srcs: (570, 209)(2967) 5 --> (2967) 5:NI0, pass, PENB
			10'd241 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 48 -> 56
			// srcs: (571, 214)(3057) -5 --> (3057) -5:PUNB, pass, NI0
			10'd242 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 32 -> 57
			// srcs: (572, 215)(2280) 0 --> (2280) 0:PUGB4, pass, PENB
			10'd243 : rdata = 48'b110001110000100100000000000000000000000100000000;
			// PEs: 56 -> 57
			// srcs: (578, 216)(3057) -5 --> (3057) -5:NI0, pass, PENB
			10'd244 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 32 -> 57
			// srcs: (579, 217)(2289) 0 --> (2289) 0:PUGB4, pass, PENB
			10'd245 : rdata = 48'b110001110000100100000000000000000000000100000000;
			// PEs: 8 -> 56
			// srcs: (580, 221)(3094) -3 --> (3094) -3:PUGB1, pass, NI0
			10'd246 : rdata = 48'b110001110000001100000000000100000000000000000000;
			// PEs: 48 -> 57
			// srcs: (581, 222)(2317) 0 --> (2317) 0:PUNB, pass, PENB
			10'd247 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 57 -> 0
			// srcs: (586, 274)(3067) -2 --> (3067) -2:PEGB1, pass, PUNB
			10'd248 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 56 -> 57
			// srcs: (587, 223)(3094) -3 --> (3094) -3:NI0, pass, PENB
			10'd249 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 16 -> 56
			// srcs: (588, 224)(3102) 0 --> (3102) 0:PUGB2, pass, NI0
			10'd250 : rdata = 48'b110001110000010100000000000100000000000000000000;
			// PEs: 48 -> 57
			// srcs: (589, 225)(2326) -2 --> (2326) -2:PUNB, pass, PENB
			10'd251 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 57 -> 0
			// srcs: (594, 275)(3095) -3 --> (3095) -3:PEGB1, pass, PUNB
			10'd252 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 56 -> 57
			// srcs: (595, 226)(3102) 0 --> (3102) 0:NI0, pass, PENB
			10'd253 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 48 -> 57
			// srcs: (596, 234)(2377) -6 --> (2377) -6:PUNB, pass, PENB
			10'd254 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 48 -> 60
			// srcs: (597, 237)(2448) 3 --> (2448) 3:PUNB, pass, PEGB4
			10'd255 : rdata = 48'b110001101111111100000000000000000000000011000000;
			// PEs: 32 -> 56
			// srcs: (598, 238)(2461) -2 --> (2461) -2:PUGB4, pass, NI0
			10'd256 : rdata = 48'b110001110000100100000000000100000000000000000000;
			// PEs: 0 -> 57
			// srcs: (599, 239)(2463) 2 --> (2463) 2:PUGB0, pass, PENB
			10'd257 : rdata = 48'b110001110000000100000000000000000000000100000000;
			// PEs: 57 -> 0
			// srcs: (603, 280)(2378) -1 --> (2378) -1:PEGB1, pass, PUNB
			10'd258 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 56 -> 57
			// srcs: (605, 240)(2461) -2 --> (2461) -2:NI0, pass, PENB
			10'd259 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 48 -> 56
			// srcs: (606, 243)(2509) 3 --> (2509) 3:PUNB, pass, NI0
			10'd260 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 16 -> 57
			// srcs: (607, 244)(2511) -2 --> (2511) -2:PUGB2, pass, PENB
			10'd261 : rdata = 48'b110001110000010100000000000000000000000100000000;
			// PEs: 60 -> 8
			// srcs: (609, 284)(2449) 6 --> (2449) 6:PEGB4, pass, PUGB1
			10'd262 : rdata = 48'b110001110000100000000000000000000000000000001001;
			// PEs: 61 -> 0
			// srcs: (611, 288)(2580) -21 --> (2580) -21:PEGB5, pass, PUNB
			10'd263 : rdata = 48'b110001110000101000000000000000000000001000000000;
			// PEs: 57 -> 24
			// srcs: (612, 285)(2464) 0 --> (2464) 0:PEGB1, pass, PUGB3
			10'd264 : rdata = 48'b110001110000001000000000000000000000000000001011;
			// PEs: 56 -> 57
			// srcs: (613, 245)(2509) 3 --> (2509) 3:NI0, pass, PENB
			10'd265 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 40 -> 57
			// srcs: (614, 247)(2572) -1 --> (2572) -1:PUGB5, pass, PENB
			10'd266 : rdata = 48'b110001110000101100000000000000000000000100000000;
			// PEs: 24 -> 56
			// srcs: (615, 250)(2613) 6 --> (2613) 6:PUGB3, pass, NI0
			10'd267 : rdata = 48'b110001110000011100000000000100000000000000000000;
			// PEs: 40 -> 57
			// srcs: (616, 251)(2615) 4 --> (2615) 4:PUGB5, pass, PENB
			10'd268 : rdata = 48'b110001110000101100000000000000000000000100000000;
			// PEs: 57 -> 16
			// srcs: (620, 286)(2512) 1 --> (2512) 1:PEGB1, pass, PUGB2
			10'd269 : rdata = 48'b110001110000001000000000000000000000000000001010;
			// PEs: 56 -> 57
			// srcs: (622, 252)(2613) 6 --> (2613) 6:NI0, pass, PENB
			10'd270 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 8 -> 57
			// srcs: (623, 255)(2676) -9 --> (2676) -9:PUGB1, pass, PENB
			10'd271 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 56
			// srcs: (624, 260)(2784) -4 --> (2784) -4:PUGB1, pass, NI0
			10'd272 : rdata = 48'b110001110000001100000000000100000000000000000000;
			// PEs: 48 -> 60
			// srcs: (660, 256)(2733) 0 --> (2733) 0:PUNB, pass, PEGB4
			10'd273 : rdata = 48'b110001101111111100000000000000000000000011000000;
			// PEs: 48 -> 57
			// srcs: (661, 261)(2786) 4 --> (2786) 4:PUNB, pass, PENB
			10'd274 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 56 -> 57
			// srcs: (667, 262)(2784) -4 --> (2784) -4:NI0, pass, PENB
			10'd275 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 8 -> 57
			// srcs: (668, 264)(2828) 1 --> (2828) 1:PUGB1, pass, PENB
			10'd276 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 48 -> 57
			// srcs: (669, 266)(2895) 13 --> (2895) 13:PUNB, pass, PENB
			10'd277 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 24 -> 57
			// srcs: (670, 269)(2929) 5 --> (2929) 5:PUGB3, pass, PENB
			10'd278 : rdata = 48'b110001110000011100000000000000000000000100000000;
			// PEs: 48 -> 57
			// srcs: (671, 272)(2970) 2 --> (2970) 2:PUNB, pass, PENB
			10'd279 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 57 -> 32
			// srcs: (674, 291)(2787) 0 --> (2787) 0:PEGB1, pass, PUGB4
			10'd280 : rdata = 48'b110001110000001000000000000000000000000000001100;
			// PEs: 57 -> 40
			// srcs: (675, 292)(2829) -9 --> (2829) -9:PEGB1, pass, PUGB5
			10'd281 : rdata = 48'b110001110000001000000000000000000000000000001101;
			// PEs: 57 -> 8
			// srcs: (676, 296)(2898) 11 --> (2898) 11:PEGB1, pass, PUGB1
			10'd282 : rdata = 48'b110001110000001000000000000000000000000000001001;
			// PEs: 57 -> 32
			// srcs: (678, 298)(2971) 7 --> (2971) 7:PEGB1, pass, PUGB4
			10'd283 : rdata = 48'b110001110000001000000000000000000000000000001100;
			// PEs: 24 -> 57
			// srcs: (684, 273)(3060) -10 --> (3060) -10:PUGB3, pass, PENB
			10'd284 : rdata = 48'b110001110000011100000000000000000000000100000000;
			// PEs: 32 -> 57
			// srcs: (685, 276)(3101) 4 --> (3101) 4:PUGB4, pass, PENB
			10'd285 : rdata = 48'b110001110000100100000000000000000000000100000000;
			// PEs: 16 -> 56
			// srcs: (686, 277)(3106) -5 --> (3106) -5:PUGB2, pass, NI0
			10'd286 : rdata = 48'b110001110000010100000000000100000000000000000000;
			// PEs: 48 -> 57
			// srcs: (687, 278)(3108) -9 --> (3108) -9:PUNB, pass, PENB
			10'd287 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 57 -> 24
			// srcs: (692, 299)(3061) -15 --> (3061) -15:PEGB1, pass, PUGB3
			10'd288 : rdata = 48'b110001110000001000000000000000000000000000001011;
			// PEs: 56 -> 57
			// srcs: (693, 279)(3106) -5 --> (3106) -5:NI0, pass, PENB
			10'd289 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 32 -> 56
			// srcs: (694, 281)(2421) 1 --> (2421) 1:PUGB4, pass, NI0
			10'd290 : rdata = 48'b110001110000100100000000000100000000000000000000;
			// PEs: 8 -> 57
			// srcs: (695, 282)(2426) -8 --> (2426) -8:PUGB1, pass, PENB
			10'd291 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 56 -> 57
			// srcs: (701, 283)(2421) 1 --> (2421) 1:NI0, pass, PENB
			10'd292 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 57 -> 40
			// srcs: (708, 300)(2427) -7 --> (2427) -7:PEGB1, pass, PUGB5
			10'd293 : rdata = 48'b110001110000001000000000000000000000000000001101;
			// PEs: 58 -> 0
			// srcs: (709, 313)(3110) -12 --> (3110) -12:PEGB2, pass, PUNB
			10'd294 : rdata = 48'b110001110000010000000000000000000000001000000000;
			// PEs: 48 -> 57
			// srcs: (1145, 287)(2568) 8 --> (2568) 8:PUNB, pass, PENB
			10'd295 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 48 -> 57
			// srcs: (1146, 289)(2621) -1 --> (2621) -1:PUNB, pass, PENB
			10'd296 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 48 -> 57
			// srcs: (1147, 290)(2682) -1 --> (2682) -1:PUNB, pass, PENB
			10'd297 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 0 -> 56
			// srcs: (1148, 293)(2835) -6 --> (2835) -6:PUGB0, pass, NI0
			10'd298 : rdata = 48'b110001110000000100000000000100000000000000000000;
			// PEs: 24 -> 57
			// srcs: (1149, 294)(2840) -8 --> (2840) -8:PUGB3, pass, PENB
			10'd299 : rdata = 48'b110001110000011100000000000000000000000100000000;
			// PEs: 57 -> 16
			// srcs: (1153, 305)(2622) 9 --> (2622) 9:PEGB1, pass, PUGB2
			10'd300 : rdata = 48'b110001110000001000000000000000000000000000001010;
			// PEs: 57 -> 48
			// srcs: (1154, 306)(2683) -4 --> (2683) -4:PEGB1, pass, PUGB6
			10'd301 : rdata = 48'b110001110000001000000000000000000000000000001110;
			// PEs: 56 -> 57
			// srcs: (1155, 295)(2835) -6 --> (2835) -6:NI0, pass, PENB
			10'd302 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 48 -> 57
			// srcs: (1156, 297)(2937) 9 --> (2937) 9:PUNB, pass, PENB
			10'd303 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 24 -> 56
			// srcs: (1157, 301)(2465) 1 --> (2465) 1:PUGB3, pass, NI0
			10'd304 : rdata = 48'b110001110000011100000000000100000000000000000000;
			// PEs: 48 -> 57
			// srcs: (1158, 302)(2476) 7 --> (2476) 7:PUNB, pass, PENB
			10'd305 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 48 -> 60
			// srcs: (1159, 304)(2563) 3 --> (2563) 3:PUNB, pass, PEGB4
			10'd306 : rdata = 48'b110001101111111100000000000000000000000011000000;
			// PEs: 57 -> 24
			// srcs: (1162, 308)(2841) -14 --> (2841) -14:PEGB1, pass, PUGB3
			10'd307 : rdata = 48'b110001110000001000000000000000000000000000001011;
			// PEs: 56 -> 57
			// srcs: (1164, 303)(2465) 1 --> (2465) 1:NI0, pass, PENB
			10'd308 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 57 -> 0
			// srcs: (1171, 314)(2477) 8 --> (2477) 8:PEGB1, pass, PUNB
			10'd309 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 60 -> 8
			// srcs: (1172, 315)(2575) 19 --> (2575) 19:PEGB4, pass, PUGB1
			10'd310 : rdata = 48'b110001110000100000000000000000000000000000001001;
			// PEs: 48 -> 57
			// srcs: (1393, 307)(2731) 18 --> (2731) 18:PUNB, pass, PENB
			10'd311 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 24 -> 57
			// srcs: (1394, 309)(2927) -3 --> (2927) -3:PUGB3, pass, PENB
			10'd312 : rdata = 48'b110001110000011100000000000000000000000100000000;
			// PEs: 48 -> 56
			// srcs: (1398, 310)(3051) -9 --> (3051) -9:PUNB, pass, NI0
			10'd313 : rdata = 48'b110001101111111100000000000100000000000000000000;
			// PEs: 24 -> 57
			// srcs: (1399, 311)(3062) -19 --> (3062) -19:PUGB3, pass, PENB
			10'd314 : rdata = 48'b110001110000011100000000000000000000000100000000;
			// PEs: 57 -> 32
			// srcs: (1402, 317)(2939) 11 --> (2939) 11:PEGB1, pass, PUGB4
			10'd315 : rdata = 48'b110001110000001000000000000000000000000000001100;
			// PEs: 56 -> 57
			// srcs: (1406, 312)(3051) -9 --> (3051) -9:NI0, pass, PENB
			10'd316 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 40 -> 57
			// srcs: (1407, 316)(2720) -2 --> (2720) -2:PUGB5, pass, PENB
			10'd317 : rdata = 48'b110001110000101100000000000000000000000100000000;
			// PEs: 16 -> 56
			// srcs: (1408, 318)(2966) 9 --> (2966) 9:PUGB2, pass, NI0
			10'd318 : rdata = 48'b110001110000010100000000000100000000000000000000;
			// PEs: 0 -> 57
			// srcs: (1409, 319)(2989) -10 --> (2989) -10:PUGB0, pass, PENB
			10'd319 : rdata = 48'b110001110000000100000000000000000000000100000000;
			// PEs: 57 -> 0
			// srcs: (1413, 321)(3063) -28 --> (3063) -28:PEGB1, pass, PUNB
			10'd320 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 56 -> 57
			// srcs: (1415, 320)(2966) 9 --> (2966) 9:NI0, pass, PENB
			10'd321 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 48 -> 57
			// srcs: (1422, 322)(2696) -14 --> (2696) -14:PUNB, pass, PENB
			10'd322 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 57 -> 32
			// srcs: (1423, 323)(2990) -1 --> (2990) -1:PEGB1, pass, PUGB4
			10'd323 : rdata = 48'b110001110000001000000000000000000000000000001100;
			// PEs: 48 -> 57
			// srcs: (1434, 324)(2648) 52 --> (2648) 52:PUNB, pass, PENB
			10'd324 : rdata = 48'b110001101111111100000000000000000000000100000000;
			// PEs: 57 -> 0
			// srcs: (1442, 325)(2746) 74 --> (2746) 74:PEGB1, pass, PUNB
			10'd325 : rdata = 48'b110001110000001000000000000000000000001000000000;
			// PEs: 8 -> 57
			// srcs: (1542, 326)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd326 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 58
			// srcs: (1545, 327)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd327 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 59
			// srcs: (1548, 328)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd328 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 60
			// srcs: (1551, 329)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd329 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 61
			// srcs: (1554, 330)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd330 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 62
			// srcs: (1557, 331)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd331 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 63
			// srcs: (1564, 332)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd332 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 57
			// srcs: (1578, 333)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd333 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 58
			// srcs: (1580, 334)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd334 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 59
			// srcs: (1581, 335)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd335 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 60
			// srcs: (1583, 336)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd336 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 61
			// srcs: (1584, 337)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd337 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 62
			// srcs: (1586, 338)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd338 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 63
			// srcs: (1587, 339)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd339 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 57
			// srcs: (1659, 340)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd340 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 58
			// srcs: (1660, 341)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd341 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 59
			// srcs: (1661, 342)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd342 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 60
			// srcs: (1663, 343)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd343 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 61
			// srcs: (1664, 344)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd344 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 62
			// srcs: (1666, 345)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd345 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 63
			// srcs: (1667, 346)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd346 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 57
			// srcs: (1726, 347)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd347 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 58
			// srcs: (1729, 348)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd348 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 59
			// srcs: (1732, 349)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd349 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 60
			// srcs: (1735, 350)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd350 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 61
			// srcs: (1738, 351)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd351 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 57
			// srcs: (1740, 352)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd352 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 62
			// srcs: (1741, 353)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd353 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 58
			// srcs: (1742, 354)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd354 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 59
			// srcs: (1743, 355)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd355 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 63
			// srcs: (1744, 356)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd356 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 60
			// srcs: (1745, 357)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd357 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 61
			// srcs: (1746, 358)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd358 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 62
			// srcs: (1748, 359)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd359 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 63
			// srcs: (1749, 360)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd360 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 57
			// srcs: (1820, 361)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd361 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 58
			// srcs: (1822, 362)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd362 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 59
			// srcs: (1823, 363)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd363 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 60
			// srcs: (1825, 364)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd364 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 61
			// srcs: (1826, 365)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd365 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 62
			// srcs: (1828, 366)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd366 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 63
			// srcs: (1829, 367)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd367 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 57
			// srcs: (1902, 368)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd368 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 58
			// srcs: (1903, 369)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd369 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 59
			// srcs: (1904, 370)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd370 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 60
			// srcs: (1905, 371)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd371 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 61
			// srcs: (1906, 372)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd372 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 62
			// srcs: (1908, 373)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd373 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 63
			// srcs: (1909, 374)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd374 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 57
			// srcs: (1910, 375)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd375 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 58
			// srcs: (1913, 376)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd376 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 59
			// srcs: (1916, 377)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd377 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 60
			// srcs: (1919, 378)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd378 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 61
			// srcs: (1922, 379)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd379 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 62
			// srcs: (1925, 380)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd380 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 63
			// srcs: (1928, 381)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd381 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 57
			// srcs: (1982, 382)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd382 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 58
			// srcs: (1984, 383)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd383 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 59
			// srcs: (1985, 384)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd384 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 60
			// srcs: (1987, 385)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd385 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 61
			// srcs: (1988, 386)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd386 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 62
			// srcs: (1990, 387)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd387 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 63
			// srcs: (1991, 388)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd388 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 57
			// srcs: (2062, 389)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd389 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 58
			// srcs: (2064, 390)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd390 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 59
			// srcs: (2065, 391)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd391 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 60
			// srcs: (2067, 392)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd392 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 61
			// srcs: (2068, 393)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd393 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 62
			// srcs: (2070, 394)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd394 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 63
			// srcs: (2071, 395)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd395 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 57
			// srcs: (2090, 396)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd396 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 58
			// srcs: (2093, 397)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd397 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 59
			// srcs: (2096, 398)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd398 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 60
			// srcs: (2103, 399)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd399 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 61
			// srcs: (2106, 400)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd400 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 62
			// srcs: (2109, 401)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd401 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 63
			// srcs: (2112, 402)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd402 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 57
			// srcs: (2144, 403)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd403 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 58
			// srcs: (2146, 404)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd404 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 59
			// srcs: (2147, 405)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd405 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 60
			// srcs: (2148, 406)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd406 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 61
			// srcs: (2149, 407)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd407 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 62
			// srcs: (2150, 408)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd408 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 63
			// srcs: (2151, 409)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd409 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 57
			// srcs: (2224, 410)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd410 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 58
			// srcs: (2226, 411)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd411 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 59
			// srcs: (2227, 412)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd412 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 60
			// srcs: (2229, 413)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd413 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 61
			// srcs: (2230, 414)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd414 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 62
			// srcs: (2232, 415)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd415 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 63
			// srcs: (2233, 416)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd416 : rdata = 48'b110001110000001100000000000000000000000011110000;
			// PEs: 8 -> 57
			// srcs: (2274, 417)(3140) 47 --> (3140) 47:PUGB1, pass, PENB
			10'd417 : rdata = 48'b110001110000001100000000000000000000000100000000;
			// PEs: 8 -> 58
			// srcs: (2277, 418)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB2
			10'd418 : rdata = 48'b110001110000001100000000000000000000000010100000;
			// PEs: 8 -> 59
			// srcs: (2280, 419)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB3
			10'd419 : rdata = 48'b110001110000001100000000000000000000000010110000;
			// PEs: 8 -> 60
			// srcs: (2283, 420)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB4
			10'd420 : rdata = 48'b110001110000001100000000000000000000000011000000;
			// PEs: 8 -> 61
			// srcs: (2286, 421)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB5
			10'd421 : rdata = 48'b110001110000001100000000000000000000000011010000;
			// PEs: 8 -> 62
			// srcs: (2289, 422)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB6
			10'd422 : rdata = 48'b110001110000001100000000000000000000000011100000;
			// PEs: 8 -> 63
			// srcs: (2292, 423)(3140) 47 --> (3140) 47:PUGB1, pass, PEGB7
			10'd423 : rdata = 48'b110001110000001100000000000000000000000011110000;
			default : rdata = 48'b000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 57) begin
	always @(*) begin
		case(address)
			// PEs: 57, 57 -> 56
			// srcs: (1, 0)(73) 1, (858) 1 --> (1642) 1:ND0, NW0, *, PEGB0
			10'd0 : rdata = 48'b000110110000000001000000000000000000000010000000;
			// PEs: 57, 57 -> 57
			// srcs: (2, 1)(154) 0, (939) 2 --> (1723) 0:ND1, NW1, *, NI0
			10'd1 : rdata = 48'b000110110000000101000000001100000000000000000000;
			// PEs: 57, 57 -> 56
			// srcs: (3, 2)(235) -2, (1020) 2 --> (1804) -4:ND2, NW2, *, PEGB0
			10'd2 : rdata = 48'b000110110000001001000000010000000000000010000000;
			// PEs: 57, 57 -> 56
			// srcs: (4, 3)(315) 1, (1100) -1 --> (1884) -1:ND3, NW3, *, PEGB0
			10'd3 : rdata = 48'b000110110000001101000000011000000000000010000000;
			// PEs: 57, 57 -> 57
			// srcs: (5, 4)(397) -2, (1182) -1 --> (1966) 2:ND4, NW4, *, NI1
			10'd4 : rdata = 48'b000110110000010001000000100100001000000000000000;
			// PEs: 57, 57 -> 59
			// srcs: (6, 5)(477) -2, (1262) 2 --> (2046) -4:ND5, NW5, *, PEGB3
			10'd5 : rdata = 48'b000110110000010101000000101000000000000010110000;
			// PEs: 57, 57 -> 60
			// srcs: (7, 6)(557) -2, (1342) -2 --> (2126) 4:ND6, NW6, *, PEGB4
			10'd6 : rdata = 48'b000110110000011001000000110000000000000011000000;
			// PEs: 57, 57 -> 57
			// srcs: (8, 7)(639) -1, (1424) -2 --> (2208) 2:ND7, NW7, *, NI2
			10'd7 : rdata = 48'b000110110000011101000000111100010000000000000000;
			// PEs: 57, 57 -> 57
			// srcs: (9, 8)(719) -1, (1504) 2 --> (2288) -2:ND8, NW8, *, NI3
			10'd8 : rdata = 48'b000110110000100001000001000100011000000000000000;
			// PEs: 57, 57 -> 56
			// srcs: (10, 9)(37) -2, (822) -3 --> (1606) 6:ND9, NW9, *, PEGB0
			10'd9 : rdata = 48'b000110110000100101000001001000000000000010000000;
			// PEs: 57, 57 -> 57
			// srcs: (11, 10)(221) 1, (1006) 2 --> (1790) 2:ND10, NW10, *, NI4
			10'd10 : rdata = 48'b000110110000101001000001010100100000000000000000;
			// PEs: 57, 57 -> 57
			// srcs: (12, 11)(405) -3, (1190) -2 --> (1974) 6:ND11, NW11, *, NI5
			10'd11 : rdata = 48'b000110110000101101000001011100101000000000000000;
			// PEs: 57, 57 -> 57
			// srcs: (13, 12)(585) -2, (1370) 2 --> (2154) -4:ND12, NW12, *, NI6
			10'd12 : rdata = 48'b000110110000110001000001100100110000000000000000;
			// PEs: 57, 57 -> 57
			// srcs: (14, 13)(769) 0, (1554) -2 --> (2338) 0:ND13, NW13, *, NI7
			10'd13 : rdata = 48'b000110110000110101000001101100111000000000000000;
			// PEs: 56 -> 
			// srcs: (44, 14)(1679) -4 --> (1679) -4:PENB, pass, 
			10'd14 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 56, 57 -> 56
			// srcs: (50, 15)(1678) -1, (1679) -4 --> (2460) -5:PENB, ALU, +, PEGB0
			10'd15 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 56 -> 
			// srcs: (63, 16)(1957) 0 --> (1957) 0:PENB, pass, 
			10'd16 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 56, 57 -> 61
			// srcs: (69, 17)(1956) -2, (1957) 0 --> (2734) -2:PENB, ALU, +, PEGB5
			10'd17 : rdata = 48'b000011101111111000111111111000000000000011010000;
			// PEs: 56 -> 
			// srcs: (71, 18)(1960) 0 --> (1960) 0:PENB, pass, 
			10'd18 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 56, 57 -> 63
			// srcs: (77, 19)(1959) 0, (1960) 0 --> (2737) 0:PENB, ALU, +, PEGB7
			10'd19 : rdata = 48'b000011101111111000111111111000000000000011110000;
			// PEs: 56 -> 
			// srcs: (79, 20)(1963) 0 --> (1963) 0:PENB, pass, 
			10'd20 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 56, 57 -> 62
			// srcs: (85, 21)(1962) 6, (1963) 0 --> (2739) 6:PENB, ALU, +, PEGB6
			10'd21 : rdata = 48'b000011101111111000111111111000000000000011100000;
			// PEs: 56 -> 57
			// srcs: (87, 22)(2037) -1 --> (2037) -1:PENB, pass, NI8
			10'd22 : rdata = 48'b110001101111111000000000000101000000000000000000;
			// PEs: 57 -> 56
			// srcs: (89, 42)(1723) 0 --> (1723) 0:NI0, pass, PEGB0
			10'd23 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 56, 57 -> 57
			// srcs: (93, 23)(2036) 0, (2037) -1 --> (2815) -1:PENB, NI8, +, NI0
			10'd24 : rdata = 48'b000011101111111010100001000100000000000000000000;
			// PEs: 56 -> 
			// srcs: (95, 24)(2040) 0 --> (2040) 0:PENB, pass, 
			10'd25 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 56, 57 -> 56
			// srcs: (101, 25)(2039) 3, (2040) 0 --> (2820) 3:PENB, ALU, +, PEGB0
			10'd26 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 56 -> 
			// srcs: (103, 26)(2043) 3 --> (2043) 3:PENB, pass, 
			10'd27 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 56, 57 -> 57
			// srcs: (109, 27)(2042) 2, (2043) 3 --> (2822) 5:PENB, ALU, +, NI8
			10'd28 : rdata = 48'b000011101111111000111111111101000000000000000000;
			// PEs: 56 -> 
			// srcs: (111, 28)(2117) 2 --> (2117) 2:PENB, pass, 
			10'd29 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 56, 57 -> 57
			// srcs: (117, 29)(2116) -2, (2117) 2 --> (2896) 0:PENB, ALU, +, NI9
			10'd30 : rdata = 48'b000011101111111000111111111101001000000000000000;
			// PEs: 56 -> 
			// srcs: (119, 30)(2120) 9 --> (2120) 9:PENB, pass, 
			10'd31 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 56, 57 -> 57
			// srcs: (125, 31)(2119) 4, (2120) 9 --> (2899) 13:PENB, ALU, +, NI10
			10'd32 : rdata = 48'b000011101111111000111111111101010000000000000000;
			// PEs: 56 -> 
			// srcs: (127, 32)(2123) 6 --> (2123) 6:PENB, pass, 
			10'd33 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 56, 57 -> 56
			// srcs: (133, 33)(2122) 0, (2123) 6 --> (2901) 6:PENB, ALU, +, PEGB0
			10'd34 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 56 -> 
			// srcs: (135, 34)(2199) -4 --> (2199) -4:PENB, pass, 
			10'd35 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 56, 57 -> 56
			// srcs: (141, 35)(2198) 0, (2199) -4 --> (2978) -4:PENB, ALU, +, PEGB0
			10'd36 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 56 -> 
			// srcs: (143, 36)(2202) 2 --> (2202) 2:PENB, pass, 
			10'd37 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 56, 57 -> 57
			// srcs: (149, 37)(2201) 2, (2202) 2 --> (2980) 4:PENB, ALU, +, NI11
			10'd38 : rdata = 48'b000011101111111000111111111101011000000000000000;
			// PEs: 56 -> 
			// srcs: (151, 38)(2205) 2 --> (2205) 2:PENB, pass, 
			10'd39 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 56, 57 -> 56
			// srcs: (157, 39)(2204) -3, (2205) 2 --> (2983) -1:PENB, ALU, +, PEGB0
			10'd40 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 56, 57 -> 57
			// srcs: (158, 40)(2207) -4, (2208) 2 --> (2985) -2:PENB, NI2, +, NI12
			10'd41 : rdata = 48'b000011101111111010100000010101100000000000000000;
			// PEs: 56, 57 -> 57
			// srcs: (159, 41)(2287) 0, (2288) -2 --> (3066) -2:PENB, NI3, +, NI2
			10'd42 : rdata = 48'b000011101111111010100000011100010000000000000000;
			// PEs: 57 -> 60
			// srcs: (248, 43)(1966) 2 --> (1966) 2:NI1, pass, PEGB4
			10'd43 : rdata = 48'b110001010000000100000000000000000000000011000000;
			// PEs: 56 -> 
			// srcs: (250, 44)(1594) -1 --> (1594) -1:PENB, pass, 
			10'd44 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 56, 57 -> 57
			// srcs: (256, 45)(2374) 6, (1594) -1 --> (2375) 5:PENB, ALU, +, NI1
			10'd45 : rdata = 48'b000011101111111000111111111100001000000000000000;
			// PEs: 56, 60 -> 57
			// srcs: (258, 46)(2394) 6, (1615) 0 --> (2395) 6:PENB, PEGB4, +, NI3
			10'd46 : rdata = 48'b000011101111111011100001000100011000000000000000;
			// PEs: 62, 56 -> 56
			// srcs: (259, 47)(2405) -6, (2406) 4 --> (2407) -2:PEGB6, PENB, +, PEGB0
			10'd47 : rdata = 48'b000011110000110011011111110000000000000010000000;
			// PEs: 57 -> 56
			// srcs: (269, 93)(2338) 0 --> (2338) 0:NI7, pass, PEGB0
			10'd48 : rdata = 48'b110001010000011100000000000000000000000010000000;
			// PEs: 57 -> 56
			// srcs: (273, 65)(1974) 6 --> (1974) 6:NI5, pass, PEGB0
			10'd49 : rdata = 48'b110001010000010100000000000000000000000010000000;
			// PEs: 57 -> 56
			// srcs: (282, 70)(2815) -1 --> (2815) -1:NI0, pass, PEGB0
			10'd50 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 57 -> 56
			// srcs: (283, 84)(2980) 4 --> (2980) 4:NI11, pass, PEGB0
			10'd51 : rdata = 48'b110001010000101100000000000000000000000010000000;
			// PEs: 57 -> 56
			// srcs: (291, 85)(2985) -2 --> (2985) -2:NI12, pass, PEGB0
			10'd52 : rdata = 48'b110001010000110000000000000000000000000010000000;
			// PEs: 57 -> 56
			// srcs: (308, 95)(2395) 6 --> (2395) 6:NI3, pass, PEGB0
			10'd53 : rdata = 48'b110001010000001100000000000000000000000010000000;
			// PEs: 56 -> 
			// srcs: (463, 48)(1667) 4 --> (1667) 4:PENB, pass, 
			10'd54 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 56, 57 -> 60
			// srcs: (469, 49)(2445) -1, (1667) 4 --> (2446) 3:PENB, ALU, +, PEGB4
			10'd55 : rdata = 48'b000011101111111000111111111000000000000011000000;
			// PEs: 56 -> 
			// srcs: (471, 50)(1689) 0 --> (1689) 0:PENB, pass, 
			10'd56 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 56, 57 -> 56
			// srcs: (477, 51)(2468) -5, (1689) 0 --> (2469) -5:PENB, ALU, +, PEGB0
			10'd57 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 56 -> 
			// srcs: (479, 52)(1713) -2 --> (1713) -2:PENB, pass, 
			10'd58 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 56, 57 -> 56
			// srcs: (485, 53)(2491) -6, (1713) -2 --> (2492) -8:PENB, ALU, +, PEGB0
			10'd59 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 56 -> 
			// srcs: (487, 54)(1744) 1 --> (1744) 1:PENB, pass, 
			10'd60 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 56, 57 -> 56
			// srcs: (493, 55)(2521) 4, (1744) 1 --> (2522) 5:PENB, ALU, +, PEGB0
			10'd61 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 56, 57 -> 57
			// srcs: (494, 56)(2569) 7, (1790) 2 --> (2570) 9:PENB, NI4, +, NI0
			10'd62 : rdata = 48'b000011101111111010100000100100000000000000000000;
			// PEs: 56 -> 
			// srcs: (496, 57)(1824) 3 --> (1824) 3:PENB, pass, 
			10'd63 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 56, 57 -> 56
			// srcs: (502, 58)(2603) 0, (1824) 3 --> (2604) 3:PENB, ALU, +, PEGB0
			10'd64 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 56 -> 
			// srcs: (504, 59)(1842) 3 --> (1842) 3:PENB, pass, 
			10'd65 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 56, 57 -> 56
			// srcs: (510, 60)(2619) -2, (1842) 3 --> (2620) 1:PENB, ALU, +, PEGB0
			10'd66 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 56 -> 
			// srcs: (512, 61)(1866) -3 --> (1866) -3:PENB, pass, 
			10'd67 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 56, 57 -> 56
			// srcs: (518, 62)(2642) -2, (1866) -3 --> (2643) -5:PENB, ALU, +, PEGB0
			10'd68 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 56 -> 
			// srcs: (520, 63)(1894) 4 --> (1894) 4:PENB, pass, 
			10'd69 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 56, 57 -> 57
			// srcs: (526, 64)(2673) 2, (1894) 4 --> (2674) 6:PENB, ALU, +, NI3
			10'd70 : rdata = 48'b000011101111111000111111111100011000000000000000;
			// PEs: 56, 58 -> 56
			// srcs: (527, 66)(2756) -5, (1977) 0 --> (2757) -5:PENB, PEGB2, +, PEGB0
			10'd71 : rdata = 48'b000011101111111011100000100000000000000010000000;
			// PEs: 56, 60 -> 56
			// srcs: (528, 67)(2762) -6, (1983) 2 --> (2763) -4:PENB, PEGB4, +, PEGB0
			10'd72 : rdata = 48'b000011101111111011100001000000000000000010000000;
			// PEs: 56 -> 
			// srcs: (530, 68)(2001) 0 --> (2001) 0:PENB, pass, 
			10'd73 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 56, 57 -> 56
			// srcs: (536, 69)(2779) 8, (2001) 0 --> (2780) 8:PENB, ALU, +, PEGB0
			10'd74 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 57, 56 -> 56
			// srcs: (537, 71)(2822) 5, (2044) 0 --> (2823) 5:NI8, PENB, +, PEGB0
			10'd75 : rdata = 48'b000011010000100011011111110000000000000010000000;
			// PEs: 59, 56 -> 57
			// srcs: (538, 72)(2825) -6, (2047) -4 --> (2826) -10:PEGB3, PENB, +, NI4
			10'd76 : rdata = 48'b000011110000011011011111110100100000000000000000;
			// PEs: 56 -> 
			// srcs: (540, 73)(2056) 0 --> (2056) 0:PENB, pass, 
			10'd77 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 56, 57 -> 56
			// srcs: (546, 74)(2833) -6, (2056) 0 --> (2834) -6:PENB, ALU, +, PEGB0
			10'd78 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 57, 56 -> 57
			// srcs: (547, 75)(2896) 0, (2118) -2 --> (2897) -2:NI9, PENB, +, NI5
			10'd79 : rdata = 48'b000011010000100111011111110100101000000000000000;
			// PEs: 57, 56 -> 56
			// srcs: (548, 76)(2899) 13, (2121) 0 --> (2900) 13:NI10, PENB, +, PEGB0
			10'd80 : rdata = 48'b000011010000101011011111110000000000000010000000;
			// PEs: 60, 56 -> 56
			// srcs: (549, 77)(2905) 2, (2127) -2 --> (2906) 0:PEGB4, PENB, +, PEGB0
			10'd81 : rdata = 48'b000011110000100011011111110000000000000010000000;
			// PEs: 56, 57 -> 57
			// srcs: (550, 78)(2930) 4, (2154) -4 --> (2931) 0:PENB, NI6, +, NI7
			10'd82 : rdata = 48'b000011101111111010100000110100111000000000000000;
			// PEs: 56, 62 -> 56
			// srcs: (558, 79)(2951) 4, (2173) 0 --> (2952) 4:PENB, PEGB6, +, PEGB0
			10'd83 : rdata = 48'b000011101111111011100001100000000000000010000000;
			// PEs: 56 -> 
			// srcs: (559, 80)(2185) -2 --> (2185) -2:PENB, pass, 
			10'd84 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 56, 57 -> 56
			// srcs: (564, 81)(2962) -5, (2185) -2 --> (2963) -7:PENB, ALU, +, PEGB0
			10'd85 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 56 -> 
			// srcs: (566, 82)(2188) 0 --> (2188) 0:PENB, pass, 
			10'd86 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 56, 57 -> 57
			// srcs: (572, 83)(2967) 5, (2188) 0 --> (2968) 5:PENB, ALU, +, NI6
			10'd87 : rdata = 48'b000011101111111000111111111100110000000000000000;
			// PEs: 56 -> 
			// srcs: (574, 86)(2280) 0 --> (2280) 0:PENB, pass, 
			10'd88 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 56, 57 -> 57
			// srcs: (580, 87)(3057) -5, (2280) 0 --> (3058) -5:PENB, ALU, +, NI8
			10'd89 : rdata = 48'b000011101111111000111111111101000000000000000000;
			// PEs: 57, 56 -> 56
			// srcs: (581, 88)(3066) -2, (2289) 0 --> (3067) -2:NI2, PENB, +, PEGB0
			10'd90 : rdata = 48'b000011010000001011011111110000000000000010000000;
			// PEs: 56 -> 
			// srcs: (583, 89)(2317) 0 --> (2317) 0:PENB, pass, 
			10'd91 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 56, 57 -> 56
			// srcs: (589, 90)(3094) -3, (2317) 0 --> (3095) -3:PENB, ALU, +, PEGB0
			10'd92 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 56 -> 
			// srcs: (591, 91)(2326) -2 --> (2326) -2:PENB, pass, 
			10'd93 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 56, 57 -> 57
			// srcs: (597, 92)(3102) 0, (2326) -2 --> (3103) -2:PENB, ALU, +, NI2
			10'd94 : rdata = 48'b000011101111111000111111111100010000000000000000;
			// PEs: 57, 56 -> 56
			// srcs: (598, 94)(2375) 5, (2377) -6 --> (2378) -1:NI1, PENB, +, PEGB0
			10'd95 : rdata = 48'b000011010000000111011111110000000000000010000000;
			// PEs: 56 -> 
			// srcs: (601, 96)(2463) 2 --> (2463) 2:PENB, pass, 
			10'd96 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 56, 57 -> 56
			// srcs: (607, 97)(2461) -2, (2463) 2 --> (2464) 0:PENB, ALU, +, PEGB0
			10'd97 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 56 -> 
			// srcs: (609, 98)(2511) -2 --> (2511) -2:PENB, pass, 
			10'd98 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 56, 57 -> 56
			// srcs: (615, 99)(2509) 3, (2511) -2 --> (2512) 1:PENB, ALU, +, PEGB0
			10'd99 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 57, 56 -> 57
			// srcs: (616, 100)(2570) 9, (2572) -1 --> (2573) 8:NI0, PENB, +, NI1
			10'd100 : rdata = 48'b000011010000000011011111110100001000000000000000;
			// PEs: 56 -> 
			// srcs: (618, 101)(2615) 4 --> (2615) 4:PENB, pass, 
			10'd101 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 56, 57 -> 57
			// srcs: (624, 102)(2613) 6, (2615) 4 --> (2616) 10:PENB, ALU, +, NI0
			10'd102 : rdata = 48'b000011101111111000111111111100000000000000000000;
			// PEs: 57, 56 -> 57
			// srcs: (625, 103)(2674) 6, (2676) -9 --> (2677) -3:NI3, PENB, +, NI9
			10'd103 : rdata = 48'b000011010000001111011111110101001000000000000000;
			// PEs: 56 -> 
			// srcs: (663, 104)(2786) 4 --> (2786) 4:PENB, pass, 
			10'd104 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 56, 57 -> 56
			// srcs: (669, 105)(2784) -4, (2786) 4 --> (2787) 0:PENB, ALU, +, PEGB0
			10'd105 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 57, 56 -> 56
			// srcs: (670, 106)(2826) -10, (2828) 1 --> (2829) -9:NI4, PENB, +, PEGB0
			10'd106 : rdata = 48'b000011010000010011011111110000000000000010000000;
			// PEs: 56, 57 -> 56
			// srcs: (671, 107)(2895) 13, (2897) -2 --> (2898) 11:PENB, NI5, +, PEGB0
			10'd107 : rdata = 48'b000011101111111010100000101000000000000010000000;
			// PEs: 56, 57 -> 57
			// srcs: (672, 108)(2929) 5, (2931) 0 --> (2932) 5:PENB, NI7, +, NI3
			10'd108 : rdata = 48'b000011101111111010100000111100011000000000000000;
			// PEs: 57, 56 -> 56
			// srcs: (673, 109)(2968) 5, (2970) 2 --> (2971) 7:NI6, PENB, +, PEGB0
			10'd109 : rdata = 48'b000011010000011011011111110000000000000010000000;
			// PEs: 57, 56 -> 56
			// srcs: (687, 110)(3058) -5, (3060) -10 --> (3061) -15:NI8, PENB, +, PEGB0
			10'd110 : rdata = 48'b000011010000100011011111110000000000000010000000;
			// PEs: 56, 57 -> 57
			// srcs: (688, 111)(3101) 4, (3103) -2 --> (3104) 2:PENB, NI2, +, NI4
			10'd111 : rdata = 48'b000011101111111010100000010100100000000000000000;
			// PEs: 56 -> 
			// srcs: (689, 112)(3108) -9 --> (3108) -9:PENB, pass, 
			10'd112 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 56, 57 -> 58
			// srcs: (695, 113)(3106) -5, (3108) -9 --> (3109) -14:PENB, ALU, +, PENB
			10'd113 : rdata = 48'b000011101111111000111111111000000000000100000000;
			// PEs: 56 -> 57
			// srcs: (697, 114)(2426) -8 --> (2426) -8:PENB, pass, NI2
			10'd114 : rdata = 48'b110001101111111000000000000100010000000000000000;
			// PEs: 57 -> 58
			// srcs: (702, 122)(3104) 2 --> (3104) 2:NI4, pass, PENB
			10'd115 : rdata = 48'b110001010000010000000000000000000000000100000000;
			// PEs: 56, 57 -> 56
			// srcs: (703, 115)(2421) 1, (2426) -8 --> (2427) -7:PENB, NI2, +, PEGB0
			10'd116 : rdata = 48'b000011101111111010100000010000000000000010000000;
			// PEs: 56, 57 -> 60
			// srcs: (1147, 116)(2568) 8, (2573) 8 --> (2574) 16:PENB, NI1, +, PEGB4
			10'd117 : rdata = 48'b000011101111111010100000001000000000000011000000;
			// PEs: 57, 56 -> 56
			// srcs: (1148, 117)(2616) 10, (2621) -1 --> (2622) 9:NI0, PENB, +, PEGB0
			10'd118 : rdata = 48'b000011010000000011011111110000000000000010000000;
			// PEs: 57, 56 -> 56
			// srcs: (1149, 118)(2677) -3, (2682) -1 --> (2683) -4:NI9, PENB, +, PEGB0
			10'd119 : rdata = 48'b000011010000100111011111110000000000000010000000;
			// PEs: 56 -> 
			// srcs: (1151, 119)(2840) -8 --> (2840) -8:PENB, pass, 
			10'd120 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 56, 57 -> 56
			// srcs: (1157, 120)(2835) -6, (2840) -8 --> (2841) -14:PENB, ALU, +, PEGB0
			10'd121 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 57, 56 -> 57
			// srcs: (1158, 121)(2932) 5, (2937) 9 --> (2938) 14:NI3, PENB, +, NI0
			10'd122 : rdata = 48'b000011010000001111011111110100000000000000000000;
			// PEs: 56 -> 
			// srcs: (1160, 123)(2476) 7 --> (2476) 7:PENB, pass, 
			10'd123 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 56, 57 -> 56
			// srcs: (1166, 124)(2465) 1, (2476) 7 --> (2477) 8:PENB, ALU, +, PEGB0
			10'd124 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 56, 61 -> 57
			// srcs: (1396, 125)(2731) 18, (2742) 20 --> (2743) 38:PENB, PEGB5, +, NI1
			10'd125 : rdata = 48'b000011101111111011100001010100001000000000000000;
			// PEs: 56, 57 -> 56
			// srcs: (1397, 126)(2927) -3, (2938) 14 --> (2939) 11:PENB, NI0, +, PEGB0
			10'd126 : rdata = 48'b000011101111111010100000000000000000000010000000;
			// PEs: 56 -> 
			// srcs: (1401, 127)(3062) -19 --> (3062) -19:PENB, pass, 
			10'd127 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 56, 57 -> 56
			// srcs: (1408, 128)(3051) -9, (3062) -19 --> (3063) -28:PENB, ALU, +, PEGB0
			10'd128 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 56, 57 -> 57
			// srcs: (1409, 129)(2720) -2, (2743) 38 --> (2744) 36:PENB, NI1, +, NI0
			10'd129 : rdata = 48'b000011101111111010100000001100000000000000000000;
			// PEs: 56 -> 
			// srcs: (1411, 130)(2989) -10 --> (2989) -10:PENB, pass, 
			10'd130 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 56, 57 -> 56
			// srcs: (1417, 131)(2966) 9, (2989) -10 --> (2990) -1:PENB, ALU, +, PEGB0
			10'd131 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 56, 57 -> 
			// srcs: (1424, 132)(2696) -14, (2744) 36 --> (2745) 22:PENB, NI0, +, 
			10'd132 : rdata = 48'b000011101111111010100000000000000000000000000000;
			// PEs: 56, 57 -> 56
			// srcs: (1437, 133)(2648) 52, (2745) 22 --> (2746) 74:PENB, ALU, +, PEGB0
			10'd133 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 56, 57 -> 58
			// srcs: (1544, 134)(3140) 47, (37) -2 --> (3174) -94:PENB, ND9, *, PENB
			10'd134 : rdata = 48'b000111101111111001100001001000000000000100000000;
			// PEs: 57, 58 -> 57
			// srcs: (1553, 148)(822) -3, (3958) -94 --> (4742) 91:NW9, PEGB2, -, NW9
			10'd135 : rdata = 48'b000100100000100111100000100000000110010000000000;
			// PEs: 56, 57 -> 58
			// srcs: (1580, 135)(3140) 47, (73) 1 --> (3210) 47:PENB, ND0, *, PENB
			10'd136 : rdata = 48'b000111101111111001100000000000000000000100000000;
			// PEs: 57, 58 -> 57
			// srcs: (1589, 149)(858) 1, (3994) 47 --> (4778) -46:NW0, PEGB2, -, NW0
			10'd137 : rdata = 48'b000100100000000011100000100000000100000000000000;
			// PEs: 56, 57 -> 58
			// srcs: (1661, 136)(3140) 47, (154) 0 --> (3291) 0:PENB, ND1, *, PENB
			10'd138 : rdata = 48'b000111101111111001100000001000000000000100000000;
			// PEs: 57, 58 -> 57
			// srcs: (1670, 150)(939) 2, (4075) 0 --> (4859) 2:NW1, PEGB2, -, NW1
			10'd139 : rdata = 48'b000100100000000111100000100000000100010000000000;
			// PEs: 56, 57 -> 58
			// srcs: (1728, 137)(3140) 47, (221) 1 --> (3358) 47:PENB, ND10, *, PENB
			10'd140 : rdata = 48'b000111101111111001100001010000000000000100000000;
			// PEs: 57, 58 -> 57
			// srcs: (1737, 151)(1006) 2, (4142) 47 --> (4926) -45:NW10, PEGB2, -, NW10
			10'd141 : rdata = 48'b000100100000101011100000100000000110100000000000;
			// PEs: 56, 57 -> 58
			// srcs: (1742, 138)(3140) 47, (235) -2 --> (3372) -94:PENB, ND2, *, PENB
			10'd142 : rdata = 48'b000111101111111001100000010000000000000100000000;
			// PEs: 57, 58 -> 57
			// srcs: (1751, 152)(1020) 2, (4156) -94 --> (4940) 96:NW2, PEGB2, -, NW2
			10'd143 : rdata = 48'b000100100000001011100000100000000100100000000000;
			// PEs: 56, 57 -> 58
			// srcs: (1822, 139)(3140) 47, (315) 1 --> (3452) 47:PENB, ND3, *, PENB
			10'd144 : rdata = 48'b000111101111111001100000011000000000000100000000;
			// PEs: 57, 58 -> 57
			// srcs: (1831, 153)(1100) -1, (4236) 47 --> (5020) -48:NW3, PEGB2, -, NW3
			10'd145 : rdata = 48'b000100100000001111100000100000000100110000000000;
			// PEs: 56, 57 -> 58
			// srcs: (1904, 140)(3140) 47, (397) -2 --> (3534) -94:PENB, ND4, *, PENB
			10'd146 : rdata = 48'b000111101111111001100000100000000000000100000000;
			// PEs: 56, 57 -> 58
			// srcs: (1912, 141)(3140) 47, (405) -3 --> (3542) -141:PENB, ND11, *, PENB
			10'd147 : rdata = 48'b000111101111111001100001011000000000000100000000;
			// PEs: 57, 58 -> 57
			// srcs: (1913, 154)(1182) -1, (4318) -94 --> (5102) 93:NW4, PEGB2, -, NW4
			10'd148 : rdata = 48'b000100100000010011100000100000000101000000000000;
			// PEs: 57, 58 -> 57
			// srcs: (1921, 155)(1190) -2, (4326) -141 --> (5110) 139:NW11, PEGB2, -, NW11
			10'd149 : rdata = 48'b000100100000101111100000100000000110110000000000;
			// PEs: 56, 57 -> 58
			// srcs: (1984, 142)(3140) 47, (477) -2 --> (3614) -94:PENB, ND5, *, PENB
			10'd150 : rdata = 48'b000111101111111001100000101000000000000100000000;
			// PEs: 57, 58 -> 57
			// srcs: (1993, 156)(1262) 2, (4398) -94 --> (5182) 96:NW5, PEGB2, -, NW5
			10'd151 : rdata = 48'b000100100000010111100000100000000101010000000000;
			// PEs: 56, 57 -> 58
			// srcs: (2064, 143)(3140) 47, (557) -2 --> (3694) -94:PENB, ND6, *, PENB
			10'd152 : rdata = 48'b000111101111111001100000110000000000000100000000;
			// PEs: 57, 58 -> 57
			// srcs: (2073, 157)(1342) -2, (4478) -94 --> (5262) 92:NW6, PEGB2, -, NW6
			10'd153 : rdata = 48'b000100100000011011100000100000000101100000000000;
			// PEs: 56, 57 -> 58
			// srcs: (2092, 144)(3140) 47, (585) -2 --> (3722) -94:PENB, ND12, *, PENB
			10'd154 : rdata = 48'b000111101111111001100001100000000000000100000000;
			// PEs: 57, 58 -> 57
			// srcs: (2101, 158)(1370) 2, (4506) -94 --> (5290) 96:NW12, PEGB2, -, NW12
			10'd155 : rdata = 48'b000100100000110011100000100000000111000000000000;
			// PEs: 56, 57 -> 58
			// srcs: (2146, 145)(3140) 47, (639) -1 --> (3776) -47:PENB, ND7, *, PENB
			10'd156 : rdata = 48'b000111101111111001100000111000000000000100000000;
			// PEs: 57, 58 -> 57
			// srcs: (2155, 159)(1424) -2, (4560) -47 --> (5344) 45:NW7, PEGB2, -, NW7
			10'd157 : rdata = 48'b000100100000011111100000100000000101110000000000;
			// PEs: 56, 57 -> 58
			// srcs: (2226, 146)(3140) 47, (719) -1 --> (3856) -47:PENB, ND8, *, PENB
			10'd158 : rdata = 48'b000111101111111001100001000000000000000100000000;
			// PEs: 57, 58 -> 57
			// srcs: (2235, 160)(1504) 2, (4640) -47 --> (5424) 49:NW8, PEGB2, -, NW8
			10'd159 : rdata = 48'b000100100000100011100000100000000110000000000000;
			// PEs: 56, 57 -> 58
			// srcs: (2276, 147)(3140) 47, (769) 0 --> (3906) 0:PENB, ND13, *, PENB
			10'd160 : rdata = 48'b000111101111111001100001101000000000000100000000;
			// PEs: 57, 58 -> 57
			// srcs: (2285, 161)(1554) -2, (4690) 0 --> (5474) -2:NW13, PEGB2, -, NW13
			10'd161 : rdata = 48'b000100100000110111100000100000000111010000000000;
			default : rdata = 48'b000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 58) begin
	always @(*) begin
		case(address)
			// PEs: 58, 58 -> 56
			// srcs: (1, 0)(75) -1, (860) 1 --> (1644) -1:ND0, NW0, *, PEGB0
			10'd0 : rdata = 48'b000110110000000001000000000000000000000010000000;
			// PEs: 58, 58 -> 56
			// srcs: (2, 1)(155) -2, (940) -1 --> (1724) 2:ND1, NW1, *, PEGB0
			10'd1 : rdata = 48'b000110110000000101000000001000000000000010000000;
			// PEs: 58, 58 -> 56
			// srcs: (3, 2)(237) 2, (1022) 2 --> (1806) 4:ND2, NW2, *, PEGB0
			10'd2 : rdata = 48'b000110110000001001000000010000000000000010000000;
			// PEs: 58, 58 -> 56
			// srcs: (4, 3)(317) -3, (1102) 2 --> (1886) -6:ND3, NW3, *, PEGB0
			10'd3 : rdata = 48'b000110110000001101000000011000000000000010000000;
			// PEs: 58, 58 -> 58
			// srcs: (5, 4)(398) 0, (1183) 2 --> (1967) 0:ND4, NW4, *, NI0
			10'd4 : rdata = 48'b000110110000010001000000100100000000000000000000;
			// PEs: 58, 58 -> 56
			// srcs: (6, 5)(479) 1, (1264) 1 --> (2048) 1:ND5, NW5, *, PEGB0
			10'd5 : rdata = 48'b000110110000010101000000101000000000000010000000;
			// PEs: 58, 58 -> 56
			// srcs: (7, 6)(559) -2, (1344) 2 --> (2128) -4:ND6, NW6, *, PEGB0
			10'd6 : rdata = 48'b000110110000011001000000110000000000000010000000;
			// PEs: 58, 58 -> 58
			// srcs: (8, 7)(641) 1, (1426) -1 --> (2210) -1:ND7, NW7, *, NI1
			10'd7 : rdata = 48'b000110110000011101000000111100001000000000000000;
			// PEs: 58, 58 -> 61
			// srcs: (9, 8)(721) 1, (1506) 2 --> (2290) 2:ND8, NW8, *, PEGB5
			10'd8 : rdata = 48'b000110110000100001000001000000000000000011010000;
			// PEs: 58, 58 -> 56
			// srcs: (10, 9)(40) -2, (825) -3 --> (1609) 6:ND9, NW9, *, PEGB0
			10'd9 : rdata = 48'b000110110000100101000001001000000000000010000000;
			// PEs: 58, 58 -> 56
			// srcs: (11, 10)(224) 1, (1009) -1 --> (1793) -1:ND10, NW10, *, PEGB0
			10'd10 : rdata = 48'b000110110000101001000001010000000000000010000000;
			// PEs: 58, 58 -> 57
			// srcs: (12, 11)(408) 0, (1193) 2 --> (1977) 0:ND11, NW11, *, PEGB1
			10'd11 : rdata = 48'b000110110000101101000001011000000000000010010000;
			// PEs: 58, 58 -> 58
			// srcs: (13, 12)(588) -2, (1373) -2 --> (2157) 4:ND12, NW12, *, NI2
			10'd12 : rdata = 48'b000110110000110001000001100100010000000000000000;
			// PEs: 58, 58 -> 58
			// srcs: (14, 13)(772) 2, (1557) -2 --> (2341) -4:ND13, NW13, *, NI3
			10'd13 : rdata = 48'b000110110000110101000001101100011000000000000000;
			// PEs: 63 -> 
			// srcs: (15, 18)(2297) 0 --> (2297) 0:PEGB7, pass, 
			10'd14 : rdata = 48'b110001110000111000000000000000000000000000000000;
			// PEs: 62, 58 -> 58
			// srcs: (17, 19)(2296) 4, (2297) 0 --> (3075) 4:PEGB6, ALU, +, NI4
			10'd15 : rdata = 48'b000011110000110000111111111100100000000000000000;
			// PEs: 56 -> 
			// srcs: (26, 14)(1715) -2 --> (1715) -2:PEGB0, pass, 
			10'd16 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 56, 58 -> 58
			// srcs: (35, 15)(1714) 9, (1715) -2 --> (2494) 7:PEGB0, ALU, +, NI5
			10'd17 : rdata = 48'b000011110000000000111111111100101000000000000000;
			// PEs: 56 -> 
			// srcs: (58, 16)(1881) 1 --> (1881) 1:PEGB0, pass, 
			10'd18 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 56, 58 -> 56
			// srcs: (67, 17)(1880) -1, (1881) 1 --> (2661) 0:PEGB0, ALU, +, PEGB0
			10'd19 : rdata = 48'b000011110000000000111111111000000000000010000000;
			// PEs: 58 -> 56
			// srcs: (97, 20)(1967) 0 --> (1967) 0:NI0, pass, PEGB0
			10'd20 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 58 -> 56
			// srcs: (99, 23)(2157) 4 --> (2157) 4:NI2, pass, PEGB0
			10'd21 : rdata = 48'b110001010000001000000000000000000000000010000000;
			// PEs: 58 -> 56
			// srcs: (114, 21)(2210) -1 --> (2210) -1:NI1, pass, PEGB0
			10'd22 : rdata = 48'b110001010000000100000000000000000000000010000000;
			// PEs: 58 -> 56
			// srcs: (140, 22)(2494) 7 --> (2494) 7:NI5, pass, PEGB0
			10'd23 : rdata = 48'b110001010000010100000000000000000000000010000000;
			// PEs: 58 -> 56
			// srcs: (153, 24)(3075) 4 --> (3075) 4:NI4, pass, PEGB0
			10'd24 : rdata = 48'b110001010000010000000000000000000000000010000000;
			// PEs: 58 -> 56
			// srcs: (291, 25)(2341) -4 --> (2341) -4:NI3, pass, PEGB0
			10'd25 : rdata = 48'b110001010000001100000000000000000000000010000000;
			// PEs: 57 -> 
			// srcs: (697, 26)(3109) -14 --> (3109) -14:PENB, pass, 
			10'd26 : rdata = 48'b110001101111111000000000000000000000000000000000;
			// PEs: 57, 58 -> 56
			// srcs: (704, 27)(3104) 2, (3109) -14 --> (3110) -12:PENB, ALU, +, PEGB0
			10'd27 : rdata = 48'b000011101111111000111111111000000000000010000000;
			// PEs: 58, 57 -> 57
			// srcs: (1547, 42)(3) 1, (3174) -94 --> (3958) -94:NM0, PENB, *, PEGB1
			10'd28 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 56, 58 -> 
			// srcs: (1550, 28)(3140) 47, (40) -2 --> (3177) -94:PEGB0, ND9, *, 
			10'd29 : rdata = 48'b000111110000000001100001001000000000000000000000;
			// PEs: 58, 58 -> 
			// srcs: (1553, 43)(3) 1, (3177) -94 --> (3961) -94:NM0, ALU, *, 
			10'd30 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 58, 58 -> 58
			// srcs: (1556, 61)(825) -3, (3961) -94 --> (4745) 91:NW9, ALU, -, NW9
			10'd31 : rdata = 48'b000100100000100100111111111000000110010000000000;
			// PEs: 58, 57 -> 57
			// srcs: (1583, 44)(3) 1, (3210) 47 --> (3994) 47:NM0, PENB, *, PEGB1
			10'd32 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 56, 58 -> 59
			// srcs: (1585, 29)(3140) 47, (75) -1 --> (3212) -47:PEGB0, ND0, *, PENB
			10'd33 : rdata = 48'b000111110000000001100000000000000000000100000000;
			// PEs: 58, 59 -> 58
			// srcs: (1594, 62)(860) 1, (3996) -47 --> (4780) 48:NW0, PEGB3, -, NW0
			10'd34 : rdata = 48'b000100100000000011100000110000000100000000000000;
			// PEs: 58, 57 -> 57
			// srcs: (1664, 45)(3) 1, (3291) 0 --> (4075) 0:NM0, PENB, *, PEGB1
			10'd35 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 56, 58 -> 59
			// srcs: (1665, 30)(3140) 47, (155) -2 --> (3292) -94:PEGB0, ND1, *, PENB
			10'd36 : rdata = 48'b000111110000000001100000001000000000000100000000;
			// PEs: 58, 59 -> 58
			// srcs: (1674, 63)(940) -1, (4076) -94 --> (4860) 93:NW1, PEGB3, -, NW1
			10'd37 : rdata = 48'b000100100000000111100000110000000100010000000000;
			// PEs: 58, 57 -> 57
			// srcs: (1731, 46)(3) 1, (3358) 47 --> (4142) 47:NM0, PENB, *, PEGB1
			10'd38 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 56, 58 -> 
			// srcs: (1734, 31)(3140) 47, (224) 1 --> (3361) 47:PEGB0, ND10, *, 
			10'd39 : rdata = 48'b000111110000000001100001010000000000000000000000;
			// PEs: 58, 58 -> 
			// srcs: (1737, 47)(3) 1, (3361) 47 --> (4145) 47:NM0, ALU, *, 
			10'd40 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 58, 58 -> 58
			// srcs: (1740, 64)(1009) -1, (4145) 47 --> (4929) -48:NW10, ALU, -, NW10
			10'd41 : rdata = 48'b000100100000101000111111111000000110100000000000;
			// PEs: 58, 57 -> 57
			// srcs: (1745, 48)(3) 1, (3372) -94 --> (4156) -94:NM0, PENB, *, PEGB1
			10'd42 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 56, 58 -> 59
			// srcs: (1747, 32)(3140) 47, (237) 2 --> (3374) 94:PEGB0, ND2, *, PENB
			10'd43 : rdata = 48'b000111110000000001100000010000000000000100000000;
			// PEs: 58, 59 -> 58
			// srcs: (1756, 65)(1022) 2, (4158) 94 --> (4942) -92:NW2, PEGB3, -, NW2
			10'd44 : rdata = 48'b000100100000001011100000110000000100100000000000;
			// PEs: 58, 57 -> 57
			// srcs: (1825, 49)(3) 1, (3452) 47 --> (4236) 47:NM0, PENB, *, PEGB1
			10'd45 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 56, 58 -> 59
			// srcs: (1827, 33)(3140) 47, (317) -3 --> (3454) -141:PEGB0, ND3, *, PENB
			10'd46 : rdata = 48'b000111110000000001100000011000000000000100000000;
			// PEs: 58, 59 -> 58
			// srcs: (1836, 66)(1102) 2, (4238) -141 --> (5022) 143:NW3, PEGB3, -, NW3
			10'd47 : rdata = 48'b000100100000001111100000110000000100110000000000;
			// PEs: 58, 57 -> 57
			// srcs: (1907, 50)(3) 1, (3534) -94 --> (4318) -94:NM0, PENB, *, PEGB1
			10'd48 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 56, 58 -> 59
			// srcs: (1908, 34)(3140) 47, (398) 0 --> (3535) 0:PEGB0, ND4, *, PENB
			10'd49 : rdata = 48'b000111110000000001100000100000000000000100000000;
			// PEs: 58, 57 -> 57
			// srcs: (1915, 51)(3) 1, (3542) -141 --> (4326) -141:NM0, PENB, *, PEGB1
			10'd50 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 58, 59 -> 58
			// srcs: (1917, 67)(1183) 2, (4319) 0 --> (5103) 2:NW4, PEGB3, -, NW4
			10'd51 : rdata = 48'b000100100000010011100000110000000101000000000000;
			// PEs: 56, 58 -> 
			// srcs: (1918, 35)(3140) 47, (408) 0 --> (3545) 0:PEGB0, ND11, *, 
			10'd52 : rdata = 48'b000111110000000001100001011000000000000000000000;
			// PEs: 58, 58 -> 
			// srcs: (1921, 52)(3) 1, (3545) 0 --> (4329) 0:NM0, ALU, *, 
			10'd53 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 58, 58 -> 58
			// srcs: (1924, 68)(1193) 2, (4329) 0 --> (5113) 2:NW11, ALU, -, NW11
			10'd54 : rdata = 48'b000100100000101100111111111000000110110000000000;
			// PEs: 58, 57 -> 57
			// srcs: (1987, 53)(3) 1, (3614) -94 --> (4398) -94:NM0, PENB, *, PEGB1
			10'd55 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 56, 58 -> 59
			// srcs: (1989, 36)(3140) 47, (479) 1 --> (3616) 47:PEGB0, ND5, *, PENB
			10'd56 : rdata = 48'b000111110000000001100000101000000000000100000000;
			// PEs: 58, 59 -> 58
			// srcs: (1998, 69)(1264) 1, (4400) 47 --> (5184) -46:NW5, PEGB3, -, NW5
			10'd57 : rdata = 48'b000100100000010111100000110000000101010000000000;
			// PEs: 58, 57 -> 57
			// srcs: (2067, 54)(3) 1, (3694) -94 --> (4478) -94:NM0, PENB, *, PEGB1
			10'd58 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 56, 58 -> 59
			// srcs: (2069, 37)(3140) 47, (559) -2 --> (3696) -94:PEGB0, ND6, *, PENB
			10'd59 : rdata = 48'b000111110000000001100000110000000000000100000000;
			// PEs: 58, 59 -> 58
			// srcs: (2078, 70)(1344) 2, (4480) -94 --> (5264) 96:NW6, PEGB3, -, NW6
			10'd60 : rdata = 48'b000100100000011011100000110000000101100000000000;
			// PEs: 58, 57 -> 57
			// srcs: (2095, 55)(3) 1, (3722) -94 --> (4506) -94:NM0, PENB, *, PEGB1
			10'd61 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 56, 58 -> 
			// srcs: (2098, 38)(3140) 47, (588) -2 --> (3725) -94:PEGB0, ND12, *, 
			10'd62 : rdata = 48'b000111110000000001100001100000000000000000000000;
			// PEs: 58, 58 -> 
			// srcs: (2101, 56)(3) 1, (3725) -94 --> (4509) -94:NM0, ALU, *, 
			10'd63 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 58, 58 -> 58
			// srcs: (2104, 71)(1373) -2, (4509) -94 --> (5293) 92:NW12, ALU, -, NW12
			10'd64 : rdata = 48'b000100100000110000111111111000000111000000000000;
			// PEs: 58, 57 -> 57
			// srcs: (2149, 57)(3) 1, (3776) -47 --> (4560) -47:NM0, PENB, *, PEGB1
			10'd65 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 56, 58 -> 59
			// srcs: (2151, 39)(3140) 47, (641) 1 --> (3778) 47:PEGB0, ND7, *, PENB
			10'd66 : rdata = 48'b000111110000000001100000111000000000000100000000;
			// PEs: 58, 59 -> 58
			// srcs: (2160, 72)(1426) -1, (4562) 47 --> (5346) -48:NW7, PEGB3, -, NW7
			10'd67 : rdata = 48'b000100100000011111100000110000000101110000000000;
			// PEs: 58, 57 -> 57
			// srcs: (2229, 58)(3) 1, (3856) -47 --> (4640) -47:NM0, PENB, *, PEGB1
			10'd68 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 56, 58 -> 59
			// srcs: (2231, 40)(3140) 47, (721) 1 --> (3858) 47:PEGB0, ND8, *, PENB
			10'd69 : rdata = 48'b000111110000000001100001000000000000000100000000;
			// PEs: 58, 59 -> 58
			// srcs: (2240, 73)(1506) 2, (4642) 47 --> (5426) -45:NW8, PEGB3, -, NW8
			10'd70 : rdata = 48'b000100100000100011100000110000000110000000000000;
			// PEs: 58, 57 -> 57
			// srcs: (2279, 59)(3) 1, (3906) 0 --> (4690) 0:NM0, PENB, *, PEGB1
			10'd71 : rdata = 48'b000111000000000011011111110000000000000010010000;
			// PEs: 56, 58 -> 
			// srcs: (2282, 41)(3140) 47, (772) 2 --> (3909) 94:PEGB0, ND13, *, 
			10'd72 : rdata = 48'b000111110000000001100001101000000000000000000000;
			// PEs: 58, 58 -> 
			// srcs: (2285, 60)(3) 1, (3909) 94 --> (4693) 94:NM0, ALU, *, 
			10'd73 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 58, 58 -> 58
			// srcs: (2288, 74)(1557) -2, (4693) 94 --> (5477) -96:NW13, ALU, -, NW13
			10'd74 : rdata = 48'b000100100000110100111111111000000111010000000000;
			default : rdata = 48'b000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 59) begin
	always @(*) begin
		case(address)
			// PEs: 59, 59 -> 56
			// srcs: (1, 0)(76) 2, (861) -2 --> (1645) -4:ND0, NW0, *, PEGB0
			10'd0 : rdata = 48'b000110110000000001000000000000000000000010000000;
			// PEs: 59, 59 -> 56
			// srcs: (2, 1)(156) -2, (941) -3 --> (1725) 6:ND1, NW1, *, PEGB0
			10'd1 : rdata = 48'b000110110000000101000000001000000000000010000000;
			// PEs: 59, 59 -> 56
			// srcs: (3, 2)(238) 2, (1023) 2 --> (1807) 4:ND2, NW2, *, PEGB0
			10'd2 : rdata = 48'b000110110000001001000000010000000000000010000000;
			// PEs: 59, 59 -> 56
			// srcs: (4, 3)(318) -2, (1103) 1 --> (1887) -2:ND3, NW3, *, PEGB0
			10'd3 : rdata = 48'b000110110000001101000000011000000000000010000000;
			// PEs: 59, 59 -> 59
			// srcs: (5, 4)(399) 0, (1184) 2 --> (1968) 0:ND4, NW4, *, NI0
			10'd4 : rdata = 48'b000110110000010001000000100100000000000000000000;
			// PEs: 59, 59 -> 56
			// srcs: (6, 5)(480) 0, (1265) 0 --> (2049) 0:ND5, NW5, *, PEGB0
			10'd5 : rdata = 48'b000110110000010101000000101000000000000010000000;
			// PEs: 59, 59 -> 56
			// srcs: (7, 6)(560) -3, (1345) -2 --> (2129) 6:ND6, NW6, *, PEGB0
			10'd6 : rdata = 48'b000110110000011001000000110000000000000010000000;
			// PEs: 59, 59 -> 59
			// srcs: (8, 7)(642) -1, (1427) 1 --> (2211) -1:ND7, NW7, *, NI1
			10'd7 : rdata = 48'b000110110000011101000000111100001000000000000000;
			// PEs: 59, 59 -> 61
			// srcs: (9, 8)(722) -2, (1507) -2 --> (2291) 4:ND8, NW8, *, PEGB5
			10'd8 : rdata = 48'b000110110000100001000001000000000000000011010000;
			// PEs: 59, 59 -> 59
			// srcs: (10, 9)(43) 0, (828) 2 --> (1612) 0:ND9, NW9, *, NI2
			10'd9 : rdata = 48'b000110110000100101000001001100010000000000000000;
			// PEs: 59, 59 -> 60
			// srcs: (11, 10)(227) 2, (1012) -3 --> (1796) -6:ND10, NW10, *, PENB
			10'd10 : rdata = 48'b000110110000101001000001010000000000000100000000;
			// PEs: 59, 59 -> 59
			// srcs: (12, 11)(411) 2, (1196) 0 --> (1980) 0:ND11, NW11, *, NI3
			10'd11 : rdata = 48'b000110110000101101000001011100011000000000000000;
			// PEs: 59, 59 -> 59
			// srcs: (13, 12)(591) 2, (1376) 2 --> (2160) 4:ND12, NW12, *, NI4
			10'd12 : rdata = 48'b000110110000110001000001100100100000000000000000;
			// PEs: 59, 59 -> 59
			// srcs: (14, 13)(775) 0, (1560) 1 --> (2344) 0:ND13, NW13, *, NI5
			10'd13 : rdata = 48'b000110110000110101000001101100101000000000000000;
			// PEs: 56 -> 
			// srcs: (28, 14)(1718) 2 --> (1718) 2:PEGB0, pass, 
			10'd14 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 56, 59 -> 56
			// srcs: (37, 15)(1717) 0, (1718) 2 --> (2496) 2:PEGB0, ALU, +, PEGB0
			10'd15 : rdata = 48'b000011110000000000111111111000000000000010000000;
			// PEs: 59 -> 56
			// srcs: (99, 23)(1980) 0 --> (1980) 0:NI3, pass, PEGB0
			10'd16 : rdata = 48'b110001010000001100000000000000000000000010000000;
			// PEs: 59 -> 56
			// srcs: (106, 20)(1968) 0 --> (1968) 0:NI0, pass, PEGB0
			10'd17 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 56 -> 
			// srcs: (107, 16)(2045) -2 --> (2045) -2:PEGB0, pass, 
			10'd18 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 59, 57 -> 57
			// srcs: (109, 17)(2045) -2, (2046) -4 --> (2825) -6:ALU, PEGB1, +, PEGB1
			10'd19 : rdata = 48'b000010011111111111100000010000000000000010010000;
			// PEs: 59 -> 56
			// srcs: (122, 21)(2211) -1 --> (2211) -1:NI1, pass, PEGB0
			10'd20 : rdata = 48'b110001010000000100000000000000000000000010000000;
			// PEs: 59 -> 56
			// srcs: (132, 22)(1612) 0 --> (1612) 0:NI2, pass, PEGB0
			10'd21 : rdata = 48'b110001010000001000000000000000000000000010000000;
			// PEs: 56 -> 
			// srcs: (234, 18)(1721) 1 --> (1721) 1:PEGB0, pass, 
			10'd22 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 56, 59 -> 56
			// srcs: (243, 19)(1720) 6, (1721) 1 --> (2502) 7:PEGB0, ALU, +, PEGB0
			10'd23 : rdata = 48'b000011110000000000111111111000000000000010000000;
			// PEs: 59 -> 56
			// srcs: (268, 24)(2160) 4 --> (2160) 4:NI4, pass, PEGB0
			10'd24 : rdata = 48'b110001010000010000000000000000000000000010000000;
			// PEs: 59 -> 56
			// srcs: (300, 25)(2344) 0 --> (2344) 0:NI5, pass, PEGB0
			10'd25 : rdata = 48'b110001010000010100000000000000000000000010000000;
			// PEs: 56, 59 -> 
			// srcs: (1553, 26)(3140) 47, (43) 0 --> (3180) 0:PEGB0, ND9, *, 
			10'd26 : rdata = 48'b000111110000000001100001001000000000000000000000;
			// PEs: 59, 59 -> 
			// srcs: (1556, 40)(3) 1, (3180) 0 --> (3964) 0:NM0, ALU, *, 
			10'd27 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 59, 59 -> 59
			// srcs: (1559, 55)(828) 2, (3964) 0 --> (4748) 2:NW9, ALU, -, NW9
			10'd28 : rdata = 48'b000100100000100100111111111000000110010000000000;
			// PEs: 56, 59 -> 59
			// srcs: (1586, 27)(3140) 47, (76) 2 --> (3213) 94:PEGB0, ND0, *, NI0
			10'd29 : rdata = 48'b000111110000000001100000000100000000000000000000;
			// PEs: 59, 58 -> 58
			// srcs: (1588, 41)(3) 1, (3212) -47 --> (3996) -47:NM0, PENB, *, PEGB2
			10'd30 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 59, 59 -> 
			// srcs: (1589, 42)(3) 1, (3213) 94 --> (3997) 94:NM0, NI0, *, 
			10'd31 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 59, 59 -> 59
			// srcs: (1592, 56)(861) -2, (3997) 94 --> (4781) -96:NW0, ALU, -, NW0
			10'd32 : rdata = 48'b000100100000000000111111111000000100000000000000;
			// PEs: 56, 59 -> 60
			// srcs: (1666, 28)(3140) 47, (156) -2 --> (3293) -94:PEGB0, ND1, *, PENB
			10'd33 : rdata = 48'b000111110000000001100000001000000000000100000000;
			// PEs: 59, 58 -> 58
			// srcs: (1668, 43)(3) 1, (3292) -94 --> (4076) -94:NM0, PENB, *, PEGB2
			10'd34 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 59, 60 -> 59
			// srcs: (1675, 57)(941) -3, (4077) -94 --> (4861) 91:NW1, PEGB4, -, NW1
			10'd35 : rdata = 48'b000100100000000111100001000000000100010000000000;
			// PEs: 56, 59 -> 
			// srcs: (1737, 29)(3140) 47, (227) 2 --> (3364) 94:PEGB0, ND10, *, 
			10'd36 : rdata = 48'b000111110000000001100001010000000000000000000000;
			// PEs: 59, 59 -> 
			// srcs: (1740, 44)(3) 1, (3364) 94 --> (4148) 94:NM0, ALU, *, 
			10'd37 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 59, 59 -> 59
			// srcs: (1743, 58)(1012) -3, (4148) 94 --> (4932) -97:NW10, ALU, -, NW10
			10'd38 : rdata = 48'b000100100000101000111111111000000110100000000000;
			// PEs: 56, 59 -> 60
			// srcs: (1748, 30)(3140) 47, (238) 2 --> (3375) 94:PEGB0, ND2, *, PENB
			10'd39 : rdata = 48'b000111110000000001100000010000000000000100000000;
			// PEs: 59, 58 -> 58
			// srcs: (1750, 45)(3) 1, (3374) 94 --> (4158) 94:NM0, PENB, *, PEGB2
			10'd40 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 59, 60 -> 59
			// srcs: (1757, 59)(1023) 2, (4159) 94 --> (4943) -92:NW2, PEGB4, -, NW2
			10'd41 : rdata = 48'b000100100000001011100001000000000100100000000000;
			// PEs: 56, 59 -> 60
			// srcs: (1828, 31)(3140) 47, (318) -2 --> (3455) -94:PEGB0, ND3, *, PENB
			10'd42 : rdata = 48'b000111110000000001100000011000000000000100000000;
			// PEs: 59, 58 -> 58
			// srcs: (1830, 46)(3) 1, (3454) -141 --> (4238) -141:NM0, PENB, *, PEGB2
			10'd43 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 59, 60 -> 59
			// srcs: (1837, 60)(1103) 1, (4239) -94 --> (5023) 95:NW3, PEGB4, -, NW3
			10'd44 : rdata = 48'b000100100000001111100001000000000100110000000000;
			// PEs: 56, 59 -> 60
			// srcs: (1909, 32)(3140) 47, (399) 0 --> (3536) 0:PEGB0, ND4, *, PENB
			10'd45 : rdata = 48'b000111110000000001100000100000000000000100000000;
			// PEs: 59, 58 -> 58
			// srcs: (1911, 47)(3) 1, (3535) 0 --> (4319) 0:NM0, PENB, *, PEGB2
			10'd46 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 59, 60 -> 59
			// srcs: (1918, 61)(1184) 2, (4320) 0 --> (5104) 2:NW4, PEGB4, -, NW4
			10'd47 : rdata = 48'b000100100000010011100001000000000101000000000000;
			// PEs: 56, 59 -> 
			// srcs: (1921, 33)(3140) 47, (411) 2 --> (3548) 94:PEGB0, ND11, *, 
			10'd48 : rdata = 48'b000111110000000001100001011000000000000000000000;
			// PEs: 59, 59 -> 
			// srcs: (1924, 48)(3) 1, (3548) 94 --> (4332) 94:NM0, ALU, *, 
			10'd49 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 59, 59 -> 59
			// srcs: (1927, 62)(1196) 0, (4332) 94 --> (5116) -94:NW11, ALU, -, NW11
			10'd50 : rdata = 48'b000100100000101100111111111000000110110000000000;
			// PEs: 56, 59 -> 60
			// srcs: (1990, 34)(3140) 47, (480) 0 --> (3617) 0:PEGB0, ND5, *, PENB
			10'd51 : rdata = 48'b000111110000000001100000101000000000000100000000;
			// PEs: 59, 58 -> 58
			// srcs: (1992, 49)(3) 1, (3616) 47 --> (4400) 47:NM0, PENB, *, PEGB2
			10'd52 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 59, 60 -> 59
			// srcs: (1999, 63)(1265) 0, (4401) 0 --> (5185) 0:NW5, PEGB4, -, NW5
			10'd53 : rdata = 48'b000100100000010111100001000000000101010000000000;
			// PEs: 56, 59 -> 60
			// srcs: (2070, 35)(3140) 47, (560) -3 --> (3697) -141:PEGB0, ND6, *, PENB
			10'd54 : rdata = 48'b000111110000000001100000110000000000000100000000;
			// PEs: 59, 58 -> 58
			// srcs: (2072, 50)(3) 1, (3696) -94 --> (4480) -94:NM0, PENB, *, PEGB2
			10'd55 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 59, 60 -> 59
			// srcs: (2079, 64)(1345) -2, (4481) -141 --> (5265) 139:NW6, PEGB4, -, NW6
			10'd56 : rdata = 48'b000100100000011011100001000000000101100000000000;
			// PEs: 56, 59 -> 
			// srcs: (2101, 36)(3140) 47, (591) 2 --> (3728) 94:PEGB0, ND12, *, 
			10'd57 : rdata = 48'b000111110000000001100001100000000000000000000000;
			// PEs: 59, 59 -> 
			// srcs: (2104, 51)(3) 1, (3728) 94 --> (4512) 94:NM0, ALU, *, 
			10'd58 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 59, 59 -> 59
			// srcs: (2107, 65)(1376) 2, (4512) 94 --> (5296) -92:NW12, ALU, -, NW12
			10'd59 : rdata = 48'b000100100000110000111111111000000111000000000000;
			// PEs: 56, 59 -> 60
			// srcs: (2152, 37)(3140) 47, (642) -1 --> (3779) -47:PEGB0, ND7, *, PENB
			10'd60 : rdata = 48'b000111110000000001100000111000000000000100000000;
			// PEs: 59, 58 -> 58
			// srcs: (2154, 52)(3) 1, (3778) 47 --> (4562) 47:NM0, PENB, *, PEGB2
			10'd61 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 59, 60 -> 59
			// srcs: (2161, 66)(1427) 1, (4563) -47 --> (5347) 48:NW7, PEGB4, -, NW7
			10'd62 : rdata = 48'b000100100000011111100001000000000101110000000000;
			// PEs: 56, 59 -> 60
			// srcs: (2232, 38)(3140) 47, (722) -2 --> (3859) -94:PEGB0, ND8, *, PENB
			10'd63 : rdata = 48'b000111110000000001100001000000000000000100000000;
			// PEs: 59, 58 -> 58
			// srcs: (2234, 53)(3) 1, (3858) 47 --> (4642) 47:NM0, PENB, *, PEGB2
			10'd64 : rdata = 48'b000111000000000011011111110000000000000010100000;
			// PEs: 59, 60 -> 59
			// srcs: (2241, 67)(1507) -2, (4643) -94 --> (5427) 92:NW8, PEGB4, -, NW8
			10'd65 : rdata = 48'b000100100000100011100001000000000110000000000000;
			// PEs: 56, 59 -> 
			// srcs: (2285, 39)(3140) 47, (775) 0 --> (3912) 0:PEGB0, ND13, *, 
			10'd66 : rdata = 48'b000111110000000001100001101000000000000000000000;
			// PEs: 59, 59 -> 
			// srcs: (2288, 54)(3) 1, (3912) 0 --> (4696) 0:NM0, ALU, *, 
			10'd67 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 59, 59 -> 59
			// srcs: (2291, 68)(1560) 1, (4696) 0 --> (5480) 1:NW13, ALU, -, NW13
			10'd68 : rdata = 48'b000100100000110100111111111000000111010000000000;
			default : rdata = 48'b000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 60) begin
	always @(*) begin
		case(address)
			// PEs: 60, 60 -> 56
			// srcs: (1, 0)(78) -2, (863) -1 --> (1647) 2:ND0, NW0, *, PEGB0
			10'd0 : rdata = 48'b000110110000000001000000000000000000000010000000;
			// PEs: 60, 60 -> 56
			// srcs: (2, 1)(158) 2, (943) 0 --> (1727) 0:ND1, NW1, *, PEGB0
			10'd1 : rdata = 48'b000110110000000101000000001000000000000010000000;
			// PEs: 60, 60 -> 56
			// srcs: (3, 2)(240) -3, (1025) -1 --> (1809) 3:ND2, NW2, *, PEGB0
			10'd2 : rdata = 48'b000110110000001001000000010000000000000010000000;
			// PEs: 60, 60 -> 56
			// srcs: (4, 3)(320) -3, (1105) 0 --> (1889) 0:ND3, NW3, *, PEGB0
			10'd3 : rdata = 48'b000110110000001101000000011000000000000010000000;
			// PEs: 60, 60 -> 56
			// srcs: (5, 4)(400) 2, (1185) -3 --> (1969) -6:ND4, NW4, *, PEGB0
			10'd4 : rdata = 48'b000110110000010001000000100000000000000010000000;
			// PEs: 60, 60 -> 56
			// srcs: (6, 5)(482) 2, (1267) -2 --> (2051) -4:ND5, NW5, *, PEGB0
			10'd5 : rdata = 48'b000110110000010101000000101000000000000010000000;
			// PEs: 60, 60 -> 56
			// srcs: (7, 6)(562) 1, (1347) 2 --> (2131) 2:ND6, NW6, *, PEGB0
			10'd6 : rdata = 48'b000110110000011001000000110000000000000010000000;
			// PEs: 60, 60 -> 56
			// srcs: (8, 7)(643) -3, (1428) 0 --> (2212) 0:ND7, NW7, *, PEGB0
			10'd7 : rdata = 48'b000110110000011101000000111000000000000010000000;
			// PEs: 60, 60 -> 62
			// srcs: (9, 8)(724) -3, (1509) 1 --> (2293) -3:ND8, NW8, *, PEGB6
			10'd8 : rdata = 48'b000110110000100001000001000000000000000011100000;
			// PEs: 60, 60 -> 57
			// srcs: (10, 9)(46) -1, (831) 0 --> (1615) 0:ND9, NW9, *, PEGB1
			10'd9 : rdata = 48'b000110110000100101000001001000000000000010010000;
			// PEs: 60, 60 -> 61
			// srcs: (11, 10)(230) 2, (1015) -2 --> (1799) -4:ND10, NW10, *, PENB
			10'd10 : rdata = 48'b000110110000101001000001010000000000000100000000;
			// PEs: 60, 60 -> 57
			// srcs: (12, 11)(414) 1, (1199) 2 --> (1983) 2:ND11, NW11, *, PEGB1
			10'd11 : rdata = 48'b000110110000101101000001011000000000000010010000;
			// PEs: 60, 60 -> 56
			// srcs: (13, 12)(598) -1, (1383) 1 --> (2167) -1:ND12, NW12, *, PEGB0
			10'd12 : rdata = 48'b000110110000110001000001100000000000000010000000;
			// PEs: 60, 60 -> 56
			// srcs: (14, 13)(778) 1, (1563) 2 --> (2347) 2:ND13, NW13, *, PEGB0
			10'd13 : rdata = 48'b000110110000110101000001101000000000000010000000;
			// PEs: 56 -> 
			// srcs: (38, 14)(1795) -4 --> (1795) -4:PEGB0, pass, 
			10'd14 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 56, 60 -> 
			// srcs: (48, 15)(1794) 0, (1795) -4 --> (2576) -4:PEGB0, ALU, +, 
			10'd15 : rdata = 48'b000011110000000000111111111000000000000000000000;
			// PEs: 60, 59 -> 61
			// srcs: (51, 20)(2576) -4, (1796) -6 --> (2577) -10:ALU, PENB, +, PENB
			10'd16 : rdata = 48'b000010011111111111011111110000000000000100000000;
			// PEs: 56 -> 
			// srcs: (131, 16)(2125) -2 --> (2125) -2:PEGB0, pass, 
			10'd17 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 60, 57 -> 57
			// srcs: (133, 17)(2125) -2, (2126) 4 --> (2905) 2:ALU, PEGB1, +, PEGB1
			10'd18 : rdata = 48'b000010011111111111100000010000000000000010010000;
			// PEs: 56 -> 
			// srcs: (244, 18)(1965) -3 --> (1965) -3:PEGB0, pass, 
			10'd19 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 60, 57 -> 56
			// srcs: (253, 19)(1965) -3, (1966) 2 --> (2748) -1:ALU, PEGB1, +, PEGB0
			10'd20 : rdata = 48'b000010011111111111100000010000000000000010000000;
			// PEs: 56 -> 
			// srcs: (602, 21)(2448) 3 --> (2448) 3:PEGB0, pass, 
			10'd21 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 57, 60 -> 56
			// srcs: (604, 22)(2446) 3, (2448) 3 --> (2449) 6:PEGB1, ALU, +, PEGB0
			10'd22 : rdata = 48'b000011110000001000111111111000000000000010000000;
			// PEs: 56 -> 
			// srcs: (665, 23)(2733) 0 --> (2733) 0:PEGB0, pass, 
			10'd23 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 60, 61 -> 61
			// srcs: (667, 24)(2733) 0, (2735) 2 --> (2736) 2:ALU, PEGB5, +, PENB
			10'd24 : rdata = 48'b000010011111111111100001010000000000000100000000;
			// PEs: 56 -> 
			// srcs: (1164, 25)(2563) 3 --> (2563) 3:PEGB0, pass, 
			10'd25 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 60, 57 -> 56
			// srcs: (1166, 26)(2563) 3, (2574) 16 --> (2575) 19:ALU, PEGB1, +, PEGB0
			10'd26 : rdata = 48'b000010011111111111100000010000000000000010000000;
			// PEs: 56, 60 -> 
			// srcs: (1556, 27)(3140) 47, (46) -1 --> (3183) -47:PEGB0, ND9, *, 
			10'd27 : rdata = 48'b000111110000000001100001001000000000000000000000;
			// PEs: 60, 60 -> 
			// srcs: (1559, 41)(3) 1, (3183) -47 --> (3967) -47:NM0, ALU, *, 
			10'd28 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 60, 60 -> 60
			// srcs: (1562, 55)(831) 0, (3967) -47 --> (4751) 47:NW9, ALU, -, NW9
			10'd29 : rdata = 48'b000100100000100100111111111000000110010000000000;
			// PEs: 56, 60 -> 61
			// srcs: (1588, 28)(3140) 47, (78) -2 --> (3215) -94:PEGB0, ND0, *, PENB
			10'd30 : rdata = 48'b000111110000000001100000000000000000000100000000;
			// PEs: 60, 61 -> 60
			// srcs: (1597, 56)(863) -1, (3999) -94 --> (4783) 93:NW0, PEGB5, -, NW0
			10'd31 : rdata = 48'b000100100000000011100001010000000100000000000000;
			// PEs: 56, 60 -> 61
			// srcs: (1668, 29)(3140) 47, (158) 2 --> (3295) 94:PEGB0, ND1, *, PENB
			10'd32 : rdata = 48'b000111110000000001100000001000000000000100000000;
			// PEs: 60, 59 -> 59
			// srcs: (1669, 42)(3) 1, (3293) -94 --> (4077) -94:NM0, PENB, *, PEGB3
			10'd33 : rdata = 48'b000111000000000011011111110000000000000010110000;
			// PEs: 60, 61 -> 60
			// srcs: (1677, 57)(943) 0, (4079) 94 --> (4863) -94:NW1, PEGB5, -, NW1
			10'd34 : rdata = 48'b000100100000000111100001010000000100010000000000;
			// PEs: 56, 60 -> 
			// srcs: (1740, 30)(3140) 47, (230) 2 --> (3367) 94:PEGB0, ND10, *, 
			10'd35 : rdata = 48'b000111110000000001100001010000000000000000000000;
			// PEs: 60, 60 -> 
			// srcs: (1743, 43)(3) 1, (3367) 94 --> (4151) 94:NM0, ALU, *, 
			10'd36 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 60, 60 -> 60
			// srcs: (1746, 58)(1015) -2, (4151) 94 --> (4935) -96:NW10, ALU, -, NW10
			10'd37 : rdata = 48'b000100100000101000111111111000000110100000000000;
			// PEs: 56, 60 -> 61
			// srcs: (1750, 31)(3140) 47, (240) -3 --> (3377) -141:PEGB0, ND2, *, PENB
			10'd38 : rdata = 48'b000111110000000001100000010000000000000100000000;
			// PEs: 60, 59 -> 59
			// srcs: (1751, 44)(3) 1, (3375) 94 --> (4159) 94:NM0, PENB, *, PEGB3
			10'd39 : rdata = 48'b000111000000000011011111110000000000000010110000;
			// PEs: 60, 61 -> 60
			// srcs: (1759, 59)(1025) -1, (4161) -141 --> (4945) 140:NW2, PEGB5, -, NW2
			10'd40 : rdata = 48'b000100100000001011100001010000000100100000000000;
			// PEs: 56, 60 -> 61
			// srcs: (1830, 32)(3140) 47, (320) -3 --> (3457) -141:PEGB0, ND3, *, PENB
			10'd41 : rdata = 48'b000111110000000001100000011000000000000100000000;
			// PEs: 60, 59 -> 59
			// srcs: (1831, 45)(3) 1, (3455) -94 --> (4239) -94:NM0, PENB, *, PEGB3
			10'd42 : rdata = 48'b000111000000000011011111110000000000000010110000;
			// PEs: 60, 61 -> 60
			// srcs: (1839, 60)(1105) 0, (4241) -141 --> (5025) 141:NW3, PEGB5, -, NW3
			10'd43 : rdata = 48'b000100100000001111100001010000000100110000000000;
			// PEs: 56, 60 -> 61
			// srcs: (1910, 33)(3140) 47, (400) 2 --> (3537) 94:PEGB0, ND4, *, PENB
			10'd44 : rdata = 48'b000111110000000001100000100000000000000100000000;
			// PEs: 60, 59 -> 59
			// srcs: (1912, 46)(3) 1, (3536) 0 --> (4320) 0:NM0, PENB, *, PEGB3
			10'd45 : rdata = 48'b000111000000000011011111110000000000000010110000;
			// PEs: 60, 61 -> 60
			// srcs: (1919, 61)(1185) -3, (4321) 94 --> (5105) -97:NW4, PEGB5, -, NW4
			10'd46 : rdata = 48'b000100100000010011100001010000000101000000000000;
			// PEs: 56, 60 -> 
			// srcs: (1924, 34)(3140) 47, (414) 1 --> (3551) 47:PEGB0, ND11, *, 
			10'd47 : rdata = 48'b000111110000000001100001011000000000000000000000;
			// PEs: 60, 60 -> 
			// srcs: (1927, 47)(3) 1, (3551) 47 --> (4335) 47:NM0, ALU, *, 
			10'd48 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 60, 60 -> 60
			// srcs: (1930, 62)(1199) 2, (4335) 47 --> (5119) -45:NW11, ALU, -, NW11
			10'd49 : rdata = 48'b000100100000101100111111111000000110110000000000;
			// PEs: 56, 60 -> 61
			// srcs: (1992, 35)(3140) 47, (482) 2 --> (3619) 94:PEGB0, ND5, *, PENB
			10'd50 : rdata = 48'b000111110000000001100000101000000000000100000000;
			// PEs: 60, 59 -> 59
			// srcs: (1993, 48)(3) 1, (3617) 0 --> (4401) 0:NM0, PENB, *, PEGB3
			10'd51 : rdata = 48'b000111000000000011011111110000000000000010110000;
			// PEs: 60, 61 -> 60
			// srcs: (2001, 63)(1267) -2, (4403) 94 --> (5187) -96:NW5, PEGB5, -, NW5
			10'd52 : rdata = 48'b000100100000010111100001010000000101010000000000;
			// PEs: 56, 60 -> 60
			// srcs: (2072, 36)(3140) 47, (562) 1 --> (3699) 47:PEGB0, ND6, *, NI0
			10'd53 : rdata = 48'b000111110000000001100000110100000000000000000000;
			// PEs: 60, 59 -> 59
			// srcs: (2073, 49)(3) 1, (3697) -141 --> (4481) -141:NM0, PENB, *, PEGB3
			10'd54 : rdata = 48'b000111000000000011011111110000000000000010110000;
			// PEs: 60, 60 -> 
			// srcs: (2075, 50)(3) 1, (3699) 47 --> (4483) 47:NM0, NI0, *, 
			10'd55 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 60, 60 -> 60
			// srcs: (2078, 64)(1347) 2, (4483) 47 --> (5267) -45:NW6, ALU, -, NW6
			10'd56 : rdata = 48'b000100100000011000111111111000000101100000000000;
			// PEs: 56, 60 -> 
			// srcs: (2108, 37)(3140) 47, (598) -1 --> (3735) -47:PEGB0, ND12, *, 
			10'd57 : rdata = 48'b000111110000000001100001100000000000000000000000;
			// PEs: 60, 60 -> 
			// srcs: (2111, 51)(3) 1, (3735) -47 --> (4519) -47:NM0, ALU, *, 
			10'd58 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 60, 60 -> 60
			// srcs: (2114, 65)(1383) 1, (4519) -47 --> (5303) 48:NW12, ALU, -, NW12
			10'd59 : rdata = 48'b000100100000110000111111111000000111000000000000;
			// PEs: 56, 60 -> 61
			// srcs: (2153, 38)(3140) 47, (643) -3 --> (3780) -141:PEGB0, ND7, *, PENB
			10'd60 : rdata = 48'b000111110000000001100000111000000000000100000000;
			// PEs: 60, 59 -> 59
			// srcs: (2155, 52)(3) 1, (3779) -47 --> (4563) -47:NM0, PENB, *, PEGB3
			10'd61 : rdata = 48'b000111000000000011011111110000000000000010110000;
			// PEs: 60, 61 -> 60
			// srcs: (2162, 66)(1428) 0, (4564) -141 --> (5348) 141:NW7, PEGB5, -, NW7
			10'd62 : rdata = 48'b000100100000011111100001010000000101110000000000;
			// PEs: 56, 60 -> 61
			// srcs: (2234, 39)(3140) 47, (724) -3 --> (3861) -141:PEGB0, ND8, *, PENB
			10'd63 : rdata = 48'b000111110000000001100001000000000000000100000000;
			// PEs: 60, 59 -> 59
			// srcs: (2235, 53)(3) 1, (3859) -94 --> (4643) -94:NM0, PENB, *, PEGB3
			10'd64 : rdata = 48'b000111000000000011011111110000000000000010110000;
			// PEs: 60, 61 -> 60
			// srcs: (2243, 67)(1509) 1, (4645) -141 --> (5429) 142:NW8, PEGB5, -, NW8
			10'd65 : rdata = 48'b000100100000100011100001010000000110000000000000;
			// PEs: 56, 60 -> 
			// srcs: (2288, 40)(3140) 47, (778) 1 --> (3915) 47:PEGB0, ND13, *, 
			10'd66 : rdata = 48'b000111110000000001100001101000000000000000000000;
			// PEs: 60, 60 -> 
			// srcs: (2291, 54)(3) 1, (3915) 47 --> (4699) 47:NM0, ALU, *, 
			10'd67 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 60, 60 -> 60
			// srcs: (2294, 68)(1563) 2, (4699) 47 --> (5483) -45:NW13, ALU, -, NW13
			10'd68 : rdata = 48'b000100100000110100111111111000000111010000000000;
			default : rdata = 48'b000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 61) begin
	always @(*) begin
		case(address)
			// PEs: 61, 61 -> 56
			// srcs: (1, 0)(79) -3, (864) 2 --> (1648) -6:ND0, NW0, *, PEGB0
			10'd0 : rdata = 48'b000110110000000001000000000000000000000010000000;
			// PEs: 61, 61 -> 56
			// srcs: (2, 1)(159) -2, (944) -3 --> (1728) 6:ND1, NW1, *, PEGB0
			10'd1 : rdata = 48'b000110110000000101000000001000000000000010000000;
			// PEs: 61, 61 -> 56
			// srcs: (3, 2)(241) -3, (1026) -1 --> (1810) 3:ND2, NW2, *, PEGB0
			10'd2 : rdata = 48'b000110110000001001000000010000000000000010000000;
			// PEs: 61, 61 -> 56
			// srcs: (4, 3)(321) 2, (1106) -1 --> (1890) -2:ND3, NW3, *, PEGB0
			10'd3 : rdata = 48'b000110110000001101000000011000000000000010000000;
			// PEs: 61, 61 -> 56
			// srcs: (5, 4)(401) 1, (1186) 2 --> (1970) 2:ND4, NW4, *, PEGB0
			10'd4 : rdata = 48'b000110110000010001000000100000000000000010000000;
			// PEs: 61, 61 -> 56
			// srcs: (6, 5)(483) 0, (1268) 2 --> (2052) 0:ND5, NW5, *, PEGB0
			10'd5 : rdata = 48'b000110110000010101000000101000000000000010000000;
			// PEs: 61, 61 -> 56
			// srcs: (7, 6)(563) 1, (1348) -2 --> (2132) -2:ND6, NW6, *, PEGB0
			10'd6 : rdata = 48'b000110110000011001000000110000000000000010000000;
			// PEs: 61, 61 -> 56
			// srcs: (8, 7)(644) 1, (1429) 0 --> (2213) 0:ND7, NW7, *, PEGB0
			10'd7 : rdata = 48'b000110110000011101000000111000000000000010000000;
			// PEs: 61, 61 -> 62
			// srcs: (9, 8)(725) -1, (1510) -2 --> (2294) 2:ND8, NW8, *, PENB
			10'd8 : rdata = 48'b000110110000100001000001000000000000000100000000;
			// PEs: 61, 61 -> 56
			// srcs: (10, 9)(49) -3, (834) 2 --> (1618) -6:ND9, NW9, *, PEGB0
			10'd9 : rdata = 48'b000110110000100101000001001000000000000010000000;
			// PEs: 61, 61 -> 62
			// srcs: (11, 10)(233) -1, (1018) -3 --> (1802) 3:ND10, NW10, *, PENB
			10'd10 : rdata = 48'b000110110000101001000001010000000000000100000000;
			// PEs: 61, 61 -> 56
			// srcs: (12, 11)(417) 0, (1202) 2 --> (1986) 0:ND11, NW11, *, PEGB0
			10'd11 : rdata = 48'b000110110000101101000001011000000000000010000000;
			// PEs: 61, 61 -> 56
			// srcs: (13, 12)(601) 2, (1386) -3 --> (2170) -6:ND12, NW12, *, PEGB0
			10'd12 : rdata = 48'b000110110000110001000001100000000000000010000000;
			// PEs: 61, 61 -> 61
			// srcs: (14, 13)(781) 1, (1566) -3 --> (2350) -3:ND13, NW13, *, NI0
			10'd13 : rdata = 48'b000110110000110101000001101100000000000000000000;
			// PEs: 59 -> 
			// srcs: (15, 16)(2291) 4 --> (2291) 4:PEGB3, pass, 
			10'd14 : rdata = 48'b110001110000011000000000000000000000000000000000;
			// PEs: 58, 61 -> 56
			// srcs: (17, 17)(2290) 2, (2291) 4 --> (3069) 6:PEGB2, ALU, +, PEGB0
			10'd15 : rdata = 48'b000011110000010000111111111000000000000010000000;
			// PEs: 56 -> 
			// srcs: (40, 14)(1798) -3 --> (1798) -3:PEGB0, pass, 
			10'd16 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 56, 61 -> 
			// srcs: (49, 15)(1797) -4, (1798) -3 --> (2578) -7:PEGB0, ALU, +, 
			10'd17 : rdata = 48'b000011110000000000111111111000000000000000000000;
			// PEs: 61, 60 -> 
			// srcs: (52, 18)(2578) -7, (1799) -4 --> (2579) -11:ALU, PENB, +, 
			10'd18 : rdata = 48'b000010011111111111011111110000000000000000000000;
			// PEs: 60, 61 -> 61
			// srcs: (55, 22)(2577) -10, (2579) -11 --> (2580) -21:PENB, ALU, +, NI1
			10'd19 : rdata = 48'b000011101111111000111111111100001000000000000000;
			// PEs: 61 -> 56
			// srcs: (284, 21)(2350) -3 --> (2350) -3:NI0, pass, PEGB0
			10'd20 : rdata = 48'b110001010000000000000000000000000000000010000000;
			// PEs: 56 -> 
			// srcs: (516, 19)(1958) 4 --> (1958) 4:PEGB0, pass, 
			10'd21 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 57, 61 -> 60
			// srcs: (518, 20)(2734) -2, (1958) 4 --> (2735) 2:PEGB1, ALU, +, PEGB4
			10'd22 : rdata = 48'b000011110000001000111111111000000000000011000000;
			// PEs: 61 -> 56
			// srcs: (606, 23)(2580) -21 --> (2580) -21:NI1, pass, PEGB0
			10'd23 : rdata = 48'b110001010000000100000000000000000000000010000000;
			// PEs: 60, 63 -> 57
			// srcs: (673, 24)(2736) 2, (2741) 18 --> (2742) 20:PENB, PEGB7, +, PEGB1
			10'd24 : rdata = 48'b000011101111111011100001110000000000000010010000;
			// PEs: 56, 61 -> 
			// srcs: (1559, 25)(3140) 47, (49) -3 --> (3186) -141:PEGB0, ND9, *, 
			10'd25 : rdata = 48'b000111110000000001100001001000000000000000000000;
			// PEs: 61, 61 -> 
			// srcs: (1562, 39)(3) 1, (3186) -141 --> (3970) -141:NM0, ALU, *, 
			10'd26 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 61, 61 -> 61
			// srcs: (1565, 55)(834) 2, (3970) -141 --> (4754) 143:NW9, ALU, -, NW9
			10'd27 : rdata = 48'b000100100000100100111111111000000110010000000000;
			// PEs: 56, 61 -> 62
			// srcs: (1589, 26)(3140) 47, (79) -3 --> (3216) -141:PEGB0, ND0, *, PENB
			10'd28 : rdata = 48'b000111110000000001100000000000000000000100000000;
			// PEs: 61, 60 -> 60
			// srcs: (1591, 40)(3) 1, (3215) -94 --> (3999) -94:NM0, PENB, *, PEGB4
			10'd29 : rdata = 48'b000111000000000011011111110000000000000011000000;
			// PEs: 61, 62 -> 61
			// srcs: (1598, 56)(864) 2, (4000) -141 --> (4784) 143:NW0, PEGB6, -, NW0
			10'd30 : rdata = 48'b000100100000000011100001100000000100000000000000;
			// PEs: 56, 61 -> 62
			// srcs: (1669, 27)(3140) 47, (159) -2 --> (3296) -94:PEGB0, ND1, *, PENB
			10'd31 : rdata = 48'b000111110000000001100000001000000000000100000000;
			// PEs: 61, 60 -> 60
			// srcs: (1671, 41)(3) 1, (3295) 94 --> (4079) 94:NM0, PENB, *, PEGB4
			10'd32 : rdata = 48'b000111000000000011011111110000000000000011000000;
			// PEs: 61, 62 -> 61
			// srcs: (1678, 57)(944) -3, (4080) -94 --> (4864) 91:NW1, PEGB6, -, NW1
			10'd33 : rdata = 48'b000100100000000111100001100000000100010000000000;
			// PEs: 56, 61 -> 
			// srcs: (1743, 28)(3140) 47, (233) -1 --> (3370) -47:PEGB0, ND10, *, 
			10'd34 : rdata = 48'b000111110000000001100001010000000000000000000000;
			// PEs: 61, 61 -> 
			// srcs: (1746, 42)(3) 1, (3370) -47 --> (4154) -47:NM0, ALU, *, 
			10'd35 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 61, 61 -> 61
			// srcs: (1749, 58)(1018) -3, (4154) -47 --> (4938) 44:NW10, ALU, -, NW10
			10'd36 : rdata = 48'b000100100000101000111111111000000110100000000000;
			// PEs: 56, 61 -> 61
			// srcs: (1751, 29)(3140) 47, (241) -3 --> (3378) -141:PEGB0, ND2, *, NI0
			10'd37 : rdata = 48'b000111110000000001100000010100000000000000000000;
			// PEs: 61, 60 -> 60
			// srcs: (1753, 43)(3) 1, (3377) -141 --> (4161) -141:NM0, PENB, *, PEGB4
			10'd38 : rdata = 48'b000111000000000011011111110000000000000011000000;
			// PEs: 61, 61 -> 
			// srcs: (1754, 44)(3) 1, (3378) -141 --> (4162) -141:NM0, NI0, *, 
			10'd39 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 61, 61 -> 61
			// srcs: (1757, 59)(1026) -1, (4162) -141 --> (4946) 140:NW2, ALU, -, NW2
			10'd40 : rdata = 48'b000100100000001000111111111000000100100000000000;
			// PEs: 56, 61 -> 62
			// srcs: (1831, 30)(3140) 47, (321) 2 --> (3458) 94:PEGB0, ND3, *, PENB
			10'd41 : rdata = 48'b000111110000000001100000011000000000000100000000;
			// PEs: 61, 60 -> 60
			// srcs: (1833, 45)(3) 1, (3457) -141 --> (4241) -141:NM0, PENB, *, PEGB4
			10'd42 : rdata = 48'b000111000000000011011111110000000000000011000000;
			// PEs: 61, 62 -> 61
			// srcs: (1840, 60)(1106) -1, (4242) 94 --> (5026) -95:NW3, PEGB6, -, NW3
			10'd43 : rdata = 48'b000100100000001111100001100000000100110000000000;
			// PEs: 56, 61 -> 62
			// srcs: (1911, 31)(3140) 47, (401) 1 --> (3538) 47:PEGB0, ND4, *, PENB
			10'd44 : rdata = 48'b000111110000000001100000100000000000000100000000;
			// PEs: 61, 60 -> 60
			// srcs: (1913, 46)(3) 1, (3537) 94 --> (4321) 94:NM0, PENB, *, PEGB4
			10'd45 : rdata = 48'b000111000000000011011111110000000000000011000000;
			// PEs: 61, 62 -> 61
			// srcs: (1920, 61)(1186) 2, (4322) 47 --> (5106) -45:NW4, PEGB6, -, NW4
			10'd46 : rdata = 48'b000100100000010011100001100000000101000000000000;
			// PEs: 56, 61 -> 
			// srcs: (1927, 32)(3140) 47, (417) 0 --> (3554) 0:PEGB0, ND11, *, 
			10'd47 : rdata = 48'b000111110000000001100001011000000000000000000000;
			// PEs: 61, 61 -> 
			// srcs: (1930, 47)(3) 1, (3554) 0 --> (4338) 0:NM0, ALU, *, 
			10'd48 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 61, 61 -> 61
			// srcs: (1933, 62)(1202) 2, (4338) 0 --> (5122) 2:NW11, ALU, -, NW11
			10'd49 : rdata = 48'b000100100000101100111111111000000110110000000000;
			// PEs: 56, 61 -> 61
			// srcs: (1993, 33)(3140) 47, (483) 0 --> (3620) 0:PEGB0, ND5, *, NI0
			10'd50 : rdata = 48'b000111110000000001100000101100000000000000000000;
			// PEs: 61, 60 -> 60
			// srcs: (1995, 48)(3) 1, (3619) 94 --> (4403) 94:NM0, PENB, *, PEGB4
			10'd51 : rdata = 48'b000111000000000011011111110000000000000011000000;
			// PEs: 61, 61 -> 
			// srcs: (1996, 49)(3) 1, (3620) 0 --> (4404) 0:NM0, NI0, *, 
			10'd52 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 61, 61 -> 61
			// srcs: (1999, 63)(1268) 2, (4404) 0 --> (5188) 2:NW5, ALU, -, NW5
			10'd53 : rdata = 48'b000100100000010100111111111000000101010000000000;
			// PEs: 56, 61 -> 
			// srcs: (2073, 34)(3140) 47, (563) 1 --> (3700) 47:PEGB0, ND6, *, 
			10'd54 : rdata = 48'b000111110000000001100000110000000000000000000000;
			// PEs: 61, 61 -> 
			// srcs: (2076, 50)(3) 1, (3700) 47 --> (4484) 47:NM0, ALU, *, 
			10'd55 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 61, 61 -> 61
			// srcs: (2079, 64)(1348) -2, (4484) 47 --> (5268) -49:NW6, ALU, -, NW6
			10'd56 : rdata = 48'b000100100000011000111111111000000101100000000000;
			// PEs: 56, 61 -> 
			// srcs: (2111, 35)(3140) 47, (601) 2 --> (3738) 94:PEGB0, ND12, *, 
			10'd57 : rdata = 48'b000111110000000001100001100000000000000000000000;
			// PEs: 61, 61 -> 
			// srcs: (2114, 51)(3) 1, (3738) 94 --> (4522) 94:NM0, ALU, *, 
			10'd58 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 61, 61 -> 61
			// srcs: (2117, 65)(1386) -3, (4522) 94 --> (5306) -97:NW12, ALU, -, NW12
			10'd59 : rdata = 48'b000100100000110000111111111000000111000000000000;
			// PEs: 56, 61 -> 62
			// srcs: (2154, 36)(3140) 47, (644) 1 --> (3781) 47:PEGB0, ND7, *, PENB
			10'd60 : rdata = 48'b000111110000000001100000111000000000000100000000;
			// PEs: 61, 60 -> 60
			// srcs: (2156, 52)(3) 1, (3780) -141 --> (4564) -141:NM0, PENB, *, PEGB4
			10'd61 : rdata = 48'b000111000000000011011111110000000000000011000000;
			// PEs: 61, 62 -> 61
			// srcs: (2163, 66)(1429) 0, (4565) 47 --> (5349) -47:NW7, PEGB6, -, NW7
			10'd62 : rdata = 48'b000100100000011111100001100000000101110000000000;
			// PEs: 56, 61 -> 62
			// srcs: (2235, 37)(3140) 47, (725) -1 --> (3862) -47:PEGB0, ND8, *, PENB
			10'd63 : rdata = 48'b000111110000000001100001000000000000000100000000;
			// PEs: 61, 60 -> 60
			// srcs: (2237, 53)(3) 1, (3861) -141 --> (4645) -141:NM0, PENB, *, PEGB4
			10'd64 : rdata = 48'b000111000000000011011111110000000000000011000000;
			// PEs: 61, 62 -> 61
			// srcs: (2244, 67)(1510) -2, (4646) -47 --> (5430) 45:NW8, PEGB6, -, NW8
			10'd65 : rdata = 48'b000100100000100011100001100000000110000000000000;
			// PEs: 56, 61 -> 
			// srcs: (2291, 38)(3140) 47, (781) 1 --> (3918) 47:PEGB0, ND13, *, 
			10'd66 : rdata = 48'b000111110000000001100001101000000000000000000000;
			// PEs: 61, 61 -> 
			// srcs: (2294, 54)(3) 1, (3918) 47 --> (4702) 47:NM0, ALU, *, 
			10'd67 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 61, 61 -> 61
			// srcs: (2297, 68)(1566) -3, (4702) 47 --> (5486) -50:NW13, ALU, -, NW13
			10'd68 : rdata = 48'b000100100000110100111111111000000111010000000000;
			default : rdata = 48'b000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 62) begin
	always @(*) begin
		case(address)
			// PEs: 62, 62 -> 56
			// srcs: (1, 0)(81) -3, (866) -3 --> (1650) 9:ND0, NW0, *, PEGB0
			10'd0 : rdata = 48'b000110110000000001000000000000000000000010000000;
			// PEs: 62, 62 -> 56
			// srcs: (2, 1)(161) -1, (946) 0 --> (1730) 0:ND1, NW1, *, PEGB0
			10'd1 : rdata = 48'b000110110000000101000000001000000000000010000000;
			// PEs: 62, 62 -> 56
			// srcs: (3, 2)(243) -3, (1028) -1 --> (1812) 3:ND2, NW2, *, PEGB0
			10'd2 : rdata = 48'b000110110000001001000000010000000000000010000000;
			// PEs: 62, 62 -> 56
			// srcs: (4, 3)(323) 2, (1108) 1 --> (1892) 2:ND3, NW3, *, PEGB0
			10'd3 : rdata = 48'b000110110000001101000000011000000000000010000000;
			// PEs: 62, 62 -> 56
			// srcs: (5, 4)(403) 2, (1188) -1 --> (1972) -2:ND4, NW4, *, PEGB0
			10'd4 : rdata = 48'b000110110000010001000000100000000000000010000000;
			// PEs: 62, 62 -> 56
			// srcs: (6, 5)(485) -3, (1270) 2 --> (2054) -6:ND5, NW5, *, PEGB0
			10'd5 : rdata = 48'b000110110000010101000000101000000000000010000000;
			// PEs: 62, 62 -> 56
			// srcs: (7, 6)(565) -2, (1350) -1 --> (2134) 2:ND6, NW6, *, PEGB0
			10'd6 : rdata = 48'b000110110000011001000000110000000000000010000000;
			// PEs: 62, 62 -> 56
			// srcs: (8, 7)(645) 1, (1430) -3 --> (2214) -3:ND7, NW7, *, PEGB0
			10'd7 : rdata = 48'b000110110000011101000000111000000000000010000000;
			// PEs: 62, 62 -> 58
			// srcs: (9, 8)(727) 2, (1512) 2 --> (2296) 4:ND8, NW8, *, PEGB2
			10'd8 : rdata = 48'b000110110000100001000001000000000000000010100000;
			// PEs: 62, 62 -> 56
			// srcs: (10, 9)(52) 2, (837) 1 --> (1621) 2:ND9, NW9, *, PEGB0
			10'd9 : rdata = 48'b000110110000100101000001001000000000000010000000;
			// PEs: 62, 62 -> 56
			// srcs: (11, 10)(236) 0, (1021) 2 --> (1805) 0:ND10, NW10, *, PEGB0
			10'd10 : rdata = 48'b000110110000101001000001010000000000000010000000;
			// PEs: 62, 62 -> 56
			// srcs: (12, 11)(420) -2, (1205) -2 --> (1989) 4:ND11, NW11, *, PEGB0
			10'd11 : rdata = 48'b000110110000101101000001011000000000000010000000;
			// PEs: 62, 62 -> 62
			// srcs: (13, 12)(604) 0, (1389) 0 --> (2173) 0:ND12, NW12, *, NI0
			10'd12 : rdata = 48'b000110110000110001000001100100000000000000000000;
			// PEs: 62, 62 -> 62
			// srcs: (14, 13)(784) -1, (1569) -1 --> (2353) 1:ND13, NW13, *, NI1
			10'd13 : rdata = 48'b000110110000110101000001101100001000000000000000;
			// PEs: 60, 61 -> 56
			// srcs: (15, 16)(2293) -3, (2294) 2 --> (3071) -1:PEGB4, PENB, +, PEGB0
			10'd14 : rdata = 48'b000011110000100011011111110000000000000010000000;
			// PEs: 56 -> 
			// srcs: (45, 14)(1801) 0 --> (1801) 0:PEGB0, pass, 
			10'd15 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 56, 62 -> 
			// srcs: (54, 15)(1800) -2, (1801) 0 --> (2581) -2:PEGB0, ALU, +, 
			10'd16 : rdata = 48'b000011110000000000111111111000000000000000000000;
			// PEs: 62, 61 -> 62
			// srcs: (57, 19)(2581) -2, (1802) 3 --> (2582) 1:ALU, PENB, +, NI2
			10'd17 : rdata = 48'b000010011111111111011111110100010000000000000000;
			// PEs: 56 -> 
			// srcs: (200, 17)(1623) 0 --> (1623) 0:PEGB0, pass, 
			10'd18 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 56, 62 -> 57
			// srcs: (209, 18)(1622) -6, (1623) 0 --> (2405) -6:PEGB0, ALU, +, PEGB1
			10'd19 : rdata = 48'b000011110000000000111111111000000000000010010000;
			// PEs: 62 -> 56
			// srcs: (277, 23)(2353) 1 --> (2353) 1:NI1, pass, PEGB0
			10'd20 : rdata = 48'b110001010000000100000000000000000000000010000000;
			// PEs: 62 -> 56
			// srcs: (501, 24)(2582) 1 --> (2582) 1:NI2, pass, PEGB0
			10'd21 : rdata = 48'b110001010000001000000000000000000000000010000000;
			// PEs: 56 -> 
			// srcs: (518, 20)(1964) 9 --> (1964) 9:PEGB0, pass, 
			10'd22 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 57, 62 -> 63
			// srcs: (520, 21)(2739) 6, (1964) 9 --> (2740) 15:PEGB1, ALU, +, PENB
			10'd23 : rdata = 48'b000011110000001000111111111000000000000100000000;
			// PEs: 62 -> 57
			// srcs: (553, 22)(2173) 0 --> (2173) 0:NI0, pass, PEGB1
			10'd24 : rdata = 48'b110001010000000000000000000000000000000010010000;
			// PEs: 56, 62 -> 
			// srcs: (1562, 25)(3140) 47, (52) 2 --> (3189) 94:PEGB0, ND9, *, 
			10'd25 : rdata = 48'b000111110000000001100001001000000000000000000000;
			// PEs: 62, 62 -> 
			// srcs: (1565, 39)(3) 1, (3189) 94 --> (3973) 94:NM0, ALU, *, 
			10'd26 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 62, 62 -> 62
			// srcs: (1568, 56)(837) 1, (3973) 94 --> (4757) -93:NW9, ALU, -, NW9
			10'd27 : rdata = 48'b000100100000100100111111111000000110010000000000;
			// PEs: 56, 62 -> 63
			// srcs: (1591, 26)(3140) 47, (81) -3 --> (3218) -141:PEGB0, ND0, *, PENB
			10'd28 : rdata = 48'b000111110000000001100000000000000000000100000000;
			// PEs: 62, 61 -> 61
			// srcs: (1592, 40)(3) 1, (3216) -141 --> (4000) -141:NM0, PENB, *, PEGB5
			10'd29 : rdata = 48'b000111000000000011011111110000000000000011010000;
			// PEs: 62, 63 -> 62
			// srcs: (1600, 57)(866) -3, (4002) -141 --> (4786) 138:NW0, PEGB7, -, NW0
			10'd30 : rdata = 48'b000100100000000011100001110000000100000000000000;
			// PEs: 56, 62 -> 62
			// srcs: (1671, 27)(3140) 47, (161) -1 --> (3298) -47:PEGB0, ND1, *, NI0
			10'd31 : rdata = 48'b000111110000000001100000001100000000000000000000;
			// PEs: 62, 61 -> 61
			// srcs: (1672, 41)(3) 1, (3296) -94 --> (4080) -94:NM0, PENB, *, PEGB5
			10'd32 : rdata = 48'b000111000000000011011111110000000000000011010000;
			// PEs: 62, 62 -> 
			// srcs: (1674, 42)(3) 1, (3298) -47 --> (4082) -47:NM0, NI0, *, 
			10'd33 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 62, 62 -> 62
			// srcs: (1677, 58)(946) 0, (4082) -47 --> (4866) 47:NW1, ALU, -, NW1
			10'd34 : rdata = 48'b000100100000000100111111111000000100010000000000;
			// PEs: 56, 62 -> 
			// srcs: (1746, 28)(3140) 47, (236) 0 --> (3373) 0:PEGB0, ND10, *, 
			10'd35 : rdata = 48'b000111110000000001100001010000000000000000000000;
			// PEs: 62, 62 -> 
			// srcs: (1749, 43)(3) 1, (3373) 0 --> (4157) 0:NM0, ALU, *, 
			10'd36 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 62, 62 -> 62
			// srcs: (1752, 59)(1021) 2, (4157) 0 --> (4941) 2:NW10, ALU, -, NW10
			10'd37 : rdata = 48'b000100100000101000111111111000000110100000000000;
			// PEs: 56, 62 -> 
			// srcs: (1753, 29)(3140) 47, (243) -3 --> (3380) -141:PEGB0, ND2, *, 
			10'd38 : rdata = 48'b000111110000000001100000010000000000000000000000;
			// PEs: 62, 62 -> 
			// srcs: (1756, 44)(3) 1, (3380) -141 --> (4164) -141:NM0, ALU, *, 
			10'd39 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 62, 62 -> 62
			// srcs: (1759, 60)(1028) -1, (4164) -141 --> (4948) 140:NW2, ALU, -, NW2
			10'd40 : rdata = 48'b000100100000001000111111111000000100100000000000;
			// PEs: 56, 62 -> 63
			// srcs: (1833, 30)(3140) 47, (323) 2 --> (3460) 94:PEGB0, ND3, *, PENB
			10'd41 : rdata = 48'b000111110000000001100000011000000000000100000000;
			// PEs: 62, 61 -> 61
			// srcs: (1834, 45)(3) 1, (3458) 94 --> (4242) 94:NM0, PENB, *, PEGB5
			10'd42 : rdata = 48'b000111000000000011011111110000000000000011010000;
			// PEs: 62, 63 -> 62
			// srcs: (1842, 61)(1108) 1, (4244) 94 --> (5028) -93:NW3, PEGB7, -, NW3
			10'd43 : rdata = 48'b000100100000001111100001110000000100110000000000;
			// PEs: 56, 62 -> 62
			// srcs: (1913, 31)(3140) 47, (403) 2 --> (3540) 94:PEGB0, ND4, *, NI0
			10'd44 : rdata = 48'b000111110000000001100000100100000000000000000000;
			// PEs: 62, 61 -> 61
			// srcs: (1914, 46)(3) 1, (3538) 47 --> (4322) 47:NM0, PENB, *, PEGB5
			10'd45 : rdata = 48'b000111000000000011011111110000000000000011010000;
			// PEs: 62, 62 -> 
			// srcs: (1916, 47)(3) 1, (3540) 94 --> (4324) 94:NM0, NI0, *, 
			10'd46 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 62, 62 -> 62
			// srcs: (1919, 62)(1188) -1, (4324) 94 --> (5108) -95:NW4, ALU, -, NW4
			10'd47 : rdata = 48'b000100100000010000111111111000000101000000000000;
			// PEs: 56, 62 -> 
			// srcs: (1930, 32)(3140) 47, (420) -2 --> (3557) -94:PEGB0, ND11, *, 
			10'd48 : rdata = 48'b000111110000000001100001011000000000000000000000;
			// PEs: 62, 62 -> 
			// srcs: (1933, 48)(3) 1, (3557) -94 --> (4341) -94:NM0, ALU, *, 
			10'd49 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 62, 62 -> 62
			// srcs: (1936, 63)(1205) -2, (4341) -94 --> (5125) 92:NW11, ALU, -, NW11
			10'd50 : rdata = 48'b000100100000101100111111111000000110110000000000;
			// PEs: 56, 62 -> 
			// srcs: (1995, 33)(3140) 47, (485) -3 --> (3622) -141:PEGB0, ND5, *, 
			10'd51 : rdata = 48'b000111110000000001100000101000000000000000000000;
			// PEs: 62, 62 -> 
			// srcs: (1998, 49)(3) 1, (3622) -141 --> (4406) -141:NM0, ALU, *, 
			10'd52 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 62, 62 -> 62
			// srcs: (2001, 64)(1270) 2, (4406) -141 --> (5190) 143:NW5, ALU, -, NW5
			10'd53 : rdata = 48'b000100100000010100111111111000000101010000000000;
			// PEs: 56, 62 -> 
			// srcs: (2075, 34)(3140) 47, (565) -2 --> (3702) -94:PEGB0, ND6, *, 
			10'd54 : rdata = 48'b000111110000000001100000110000000000000000000000;
			// PEs: 62, 62 -> 
			// srcs: (2078, 50)(3) 1, (3702) -94 --> (4486) -94:NM0, ALU, *, 
			10'd55 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 62, 62 -> 62
			// srcs: (2081, 65)(1350) -1, (4486) -94 --> (5270) 93:NW6, ALU, -, NW6
			10'd56 : rdata = 48'b000100100000011000111111111000000101100000000000;
			// PEs: 56, 62 -> 
			// srcs: (2114, 35)(3140) 47, (604) 0 --> (3741) 0:PEGB0, ND12, *, 
			10'd57 : rdata = 48'b000111110000000001100001100000000000000000000000;
			// PEs: 62, 62 -> 
			// srcs: (2117, 51)(3) 1, (3741) 0 --> (4525) 0:NM0, ALU, *, 
			10'd58 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 62, 62 -> 62
			// srcs: (2120, 66)(1389) 0, (4525) 0 --> (5309) 0:NW12, ALU, -, NW12
			10'd59 : rdata = 48'b000100100000110000111111111000000111000000000000;
			// PEs: 56, 62 -> 63
			// srcs: (2155, 36)(3140) 47, (645) 1 --> (3782) 47:PEGB0, ND7, *, PENB
			10'd60 : rdata = 48'b000111110000000001100000111000000000000100000000;
			// PEs: 62, 61 -> 61
			// srcs: (2157, 52)(3) 1, (3781) 47 --> (4565) 47:NM0, PENB, *, PEGB5
			10'd61 : rdata = 48'b000111000000000011011111110000000000000011010000;
			// PEs: 62, 63 -> 62
			// srcs: (2164, 67)(1430) -3, (4566) 47 --> (5350) -50:NW7, PEGB7, -, NW7
			10'd62 : rdata = 48'b000100100000011111100001110000000101110000000000;
			// PEs: 56, 62 -> 62
			// srcs: (2237, 37)(3140) 47, (727) 2 --> (3864) 94:PEGB0, ND8, *, NI0
			10'd63 : rdata = 48'b000111110000000001100001000100000000000000000000;
			// PEs: 62, 61 -> 61
			// srcs: (2238, 53)(3) 1, (3862) -47 --> (4646) -47:NM0, PENB, *, PEGB5
			10'd64 : rdata = 48'b000111000000000011011111110000000000000011010000;
			// PEs: 62, 62 -> 
			// srcs: (2240, 54)(3) 1, (3864) 94 --> (4648) 94:NM0, NI0, *, 
			10'd65 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 62, 62 -> 62
			// srcs: (2243, 68)(1512) 2, (4648) 94 --> (5432) -92:NW8, ALU, -, NW8
			10'd66 : rdata = 48'b000100100000100000111111111000000110000000000000;
			// PEs: 56, 62 -> 
			// srcs: (2294, 38)(3140) 47, (784) -1 --> (3921) -47:PEGB0, ND13, *, 
			10'd67 : rdata = 48'b000111110000000001100001101000000000000000000000;
			// PEs: 62, 62 -> 
			// srcs: (2297, 55)(3) 1, (3921) -47 --> (4705) -47:NM0, ALU, *, 
			10'd68 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 62, 62 -> 62
			// srcs: (2300, 69)(1569) -1, (4705) -47 --> (5489) 46:NW13, ALU, -, NW13
			10'd69 : rdata = 48'b000100100000110100111111111000000111010000000000;
			default : rdata = 48'b000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 63) begin
	always @(*) begin
		case(address)
			// PEs: 63, 63 -> 56
			// srcs: (1, 0)(82) -1, (867) 2 --> (1651) -2:ND0, NW0, *, PENB
			10'd0 : rdata = 48'b000110110000000001000000000000000000000100000000;
			// PEs: 63, 63 -> 56
			// srcs: (2, 1)(162) -2, (947) 1 --> (1731) -2:ND1, NW1, *, PENB
			10'd1 : rdata = 48'b000110110000000101000000001000000000000100000000;
			// PEs: 63, 63 -> 56
			// srcs: (3, 2)(244) 1, (1029) 2 --> (1813) 2:ND2, NW2, *, PENB
			10'd2 : rdata = 48'b000110110000001001000000010000000000000100000000;
			// PEs: 63, 63 -> 56
			// srcs: (4, 3)(324) -3, (1109) 0 --> (1893) 0:ND3, NW3, *, PENB
			10'd3 : rdata = 48'b000110110000001101000000011000000000000100000000;
			// PEs: 63, 63 -> 56
			// srcs: (5, 4)(404) -3, (1189) 2 --> (1973) -6:ND4, NW4, *, PENB
			10'd4 : rdata = 48'b000110110000010001000000100000000000000100000000;
			// PEs: 63, 63 -> 56
			// srcs: (6, 5)(486) 0, (1271) 0 --> (2055) 0:ND5, NW5, *, PENB
			10'd5 : rdata = 48'b000110110000010101000000101000000000000100000000;
			// PEs: 63, 63 -> 56
			// srcs: (7, 6)(566) 1, (1351) -3 --> (2135) -3:ND6, NW6, *, PENB
			10'd6 : rdata = 48'b000110110000011001000000110000000000000100000000;
			// PEs: 63, 63 -> 56
			// srcs: (8, 7)(646) -2, (1431) -1 --> (2215) 2:ND7, NW7, *, PENB
			10'd7 : rdata = 48'b000110110000011101000000111000000000000100000000;
			// PEs: 63, 63 -> 58
			// srcs: (9, 8)(728) 0, (1513) 1 --> (2297) 0:ND8, NW8, *, PEGB2
			10'd8 : rdata = 48'b000110110000100001000001000000000000000010100000;
			// PEs: 63, 63 -> 56
			// srcs: (10, 9)(59) -2, (844) -1 --> (1628) 2:ND9, NW9, *, PENB
			10'd9 : rdata = 48'b000110110000100101000001001000000000000100000000;
			// PEs: 63, 63 -> 63
			// srcs: (11, 10)(239) 0, (1024) -3 --> (1808) 0:ND10, NW10, *, NI0
			10'd10 : rdata = 48'b000110110000101001000001010100000000000000000000;
			// PEs: 63, 63 -> 63
			// srcs: (12, 11)(423) -2, (1208) -2 --> (1992) 4:ND11, NW11, *, NI1
			10'd11 : rdata = 48'b000110110000101101000001011100001000000000000000;
			// PEs: 63, 63 -> 63
			// srcs: (13, 12)(607) -1, (1392) -2 --> (2176) 2:ND12, NW12, *, NI2
			10'd12 : rdata = 48'b000110110000110001000001100100010000000000000000;
			// PEs: 63, 63 -> 63
			// srcs: (14, 13)(787) 0, (1572) -1 --> (2356) 0:ND13, NW13, *, NI3
			10'd13 : rdata = 48'b000110110000110101000001101100011000000000000000;
			// PEs: 56 -> 
			// srcs: (52, 14)(1875) 0 --> (1875) 0:PEGB0, pass, 
			10'd14 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 56, 63 -> 56
			// srcs: (61, 15)(1874) -2, (1875) 0 --> (2655) -2:PEGB0, ALU, +, PENB
			10'd15 : rdata = 48'b000011110000000000111111111000000000000100000000;
			// PEs: 63 -> 56
			// srcs: (138, 21)(1992) 4 --> (1992) 4:NI1, pass, PENB
			10'd16 : rdata = 48'b110001010000000100000000000000000000000100000000;
			// PEs: 63 -> 56
			// srcs: (140, 22)(2176) 2 --> (2176) 2:NI2, pass, PENB
			10'd17 : rdata = 48'b110001010000001000000000000000000000000100000000;
			// PEs: 56 -> 
			// srcs: (251, 16)(1576) 0 --> (1576) 0:PEGB0, pass, 
			10'd18 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 56, 63 -> 56
			// srcs: (260, 17)(1575) 0, (1576) 0 --> (2358) 0:PEGB0, ALU, +, PENB
			10'd19 : rdata = 48'b000011110000000000111111111000000000000100000000;
			// PEs: 63 -> 56
			// srcs: (267, 18)(1808) 0 --> (1808) 0:NI0, pass, PENB
			10'd20 : rdata = 48'b110001010000000000000000000000000000000100000000;
			// PEs: 63 -> 56
			// srcs: (300, 23)(2356) 0 --> (2356) 0:NI3, pass, PENB
			10'd21 : rdata = 48'b110001010000001100000000000000000000000100000000;
			// PEs: 56 -> 
			// srcs: (517, 19)(1961) 3 --> (1961) 3:PEGB0, pass, 
			10'd22 : rdata = 48'b110001110000000000000000000000000000000000000000;
			// PEs: 57, 63 -> 
			// srcs: (519, 20)(2737) 0, (1961) 3 --> (2738) 3:PEGB1, ALU, +, 
			10'd23 : rdata = 48'b000011110000001000111111111000000000000000000000;
			// PEs: 63, 62 -> 61
			// srcs: (523, 24)(2738) 3, (2740) 15 --> (2741) 18:ALU, PENB, +, PEGB5
			10'd24 : rdata = 48'b000010011111111111011111110000000000000011010000;
			// PEs: 56, 63 -> 
			// srcs: (1569, 25)(3140) 47, (59) -2 --> (3196) -94:PEGB0, ND9, *, 
			10'd25 : rdata = 48'b000111110000000001100001001000000000000000000000;
			// PEs: 63, 63 -> 
			// srcs: (1572, 39)(3) 1, (3196) -94 --> (3980) -94:NM0, ALU, *, 
			10'd26 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 63, 63 -> 63
			// srcs: (1575, 56)(844) -1, (3980) -94 --> (4764) 93:NW9, ALU, -, NW9
			10'd27 : rdata = 48'b000100100000100100111111111000000110010000000000;
			// PEs: 56, 63 -> 63
			// srcs: (1592, 26)(3140) 47, (82) -1 --> (3219) -47:PEGB0, ND0, *, NI0
			10'd28 : rdata = 48'b000111110000000001100000000100000000000000000000;
			// PEs: 63, 62 -> 62
			// srcs: (1594, 40)(3) 1, (3218) -141 --> (4002) -141:NM0, PENB, *, PEGB6
			10'd29 : rdata = 48'b000111000000000011011111110000000000000011100000;
			// PEs: 63, 63 -> 
			// srcs: (1595, 41)(3) 1, (3219) -47 --> (4003) -47:NM0, NI0, *, 
			10'd30 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 63, 63 -> 63
			// srcs: (1598, 57)(867) 2, (4003) -47 --> (4787) 49:NW0, ALU, -, NW0
			10'd31 : rdata = 48'b000100100000000000111111111000000100000000000000;
			// PEs: 56, 63 -> 
			// srcs: (1672, 27)(3140) 47, (162) -2 --> (3299) -94:PEGB0, ND1, *, 
			10'd32 : rdata = 48'b000111110000000001100000001000000000000000000000;
			// PEs: 63, 63 -> 
			// srcs: (1675, 42)(3) 1, (3299) -94 --> (4083) -94:NM0, ALU, *, 
			10'd33 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 63, 63 -> 63
			// srcs: (1678, 58)(947) 1, (4083) -94 --> (4867) 95:NW1, ALU, -, NW1
			10'd34 : rdata = 48'b000100100000000100111111111000000100010000000000;
			// PEs: 56, 63 -> 
			// srcs: (1749, 28)(3140) 47, (239) 0 --> (3376) 0:PEGB0, ND10, *, 
			10'd35 : rdata = 48'b000111110000000001100001010000000000000000000000;
			// PEs: 63, 63 -> 63
			// srcs: (1752, 43)(3) 1, (3376) 0 --> (4160) 0:NM0, ALU, *, NI0
			10'd36 : rdata = 48'b000111000000000000111111111100000000000000000000;
			// PEs: 56, 63 -> 63
			// srcs: (1754, 29)(3140) 47, (244) 1 --> (3381) 47:PEGB0, ND2, *, NI1
			10'd37 : rdata = 48'b000111110000000001100000010100001000000000000000;
			// PEs: 63, 63 -> 63
			// srcs: (1755, 59)(1024) -3, (4160) 0 --> (4944) -3:NW10, NI0, -, NW10
			10'd38 : rdata = 48'b000100100000101010100000000000000110100000000000;
			// PEs: 63, 63 -> 
			// srcs: (1757, 44)(3) 1, (3381) 47 --> (4165) 47:NM0, NI1, *, 
			10'd39 : rdata = 48'b000111000000000010100000001000000000000000000000;
			// PEs: 63, 63 -> 63
			// srcs: (1760, 60)(1029) 2, (4165) 47 --> (4949) -45:NW2, ALU, -, NW2
			10'd40 : rdata = 48'b000100100000001000111111111000000100100000000000;
			// PEs: 56, 63 -> 63
			// srcs: (1834, 30)(3140) 47, (324) -3 --> (3461) -141:PEGB0, ND3, *, NI0
			10'd41 : rdata = 48'b000111110000000001100000011100000000000000000000;
			// PEs: 63, 62 -> 62
			// srcs: (1836, 45)(3) 1, (3460) 94 --> (4244) 94:NM0, PENB, *, PEGB6
			10'd42 : rdata = 48'b000111000000000011011111110000000000000011100000;
			// PEs: 63, 63 -> 
			// srcs: (1837, 46)(3) 1, (3461) -141 --> (4245) -141:NM0, NI0, *, 
			10'd43 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 63, 63 -> 63
			// srcs: (1840, 61)(1109) 0, (4245) -141 --> (5029) 141:NW3, ALU, -, NW3
			10'd44 : rdata = 48'b000100100000001100111111111000000100110000000000;
			// PEs: 56, 63 -> 
			// srcs: (1914, 31)(3140) 47, (404) -3 --> (3541) -141:PEGB0, ND4, *, 
			10'd45 : rdata = 48'b000111110000000001100000100000000000000000000000;
			// PEs: 63, 63 -> 
			// srcs: (1917, 47)(3) 1, (3541) -141 --> (4325) -141:NM0, ALU, *, 
			10'd46 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 63, 63 -> 63
			// srcs: (1920, 62)(1189) 2, (4325) -141 --> (5109) 143:NW4, ALU, -, NW4
			10'd47 : rdata = 48'b000100100000010000111111111000000101000000000000;
			// PEs: 56, 63 -> 
			// srcs: (1933, 32)(3140) 47, (423) -2 --> (3560) -94:PEGB0, ND11, *, 
			10'd48 : rdata = 48'b000111110000000001100001011000000000000000000000;
			// PEs: 63, 63 -> 
			// srcs: (1936, 48)(3) 1, (3560) -94 --> (4344) -94:NM0, ALU, *, 
			10'd49 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 63, 63 -> 63
			// srcs: (1939, 63)(1208) -2, (4344) -94 --> (5128) 92:NW11, ALU, -, NW11
			10'd50 : rdata = 48'b000100100000101100111111111000000110110000000000;
			// PEs: 56, 63 -> 
			// srcs: (1996, 33)(3140) 47, (486) 0 --> (3623) 0:PEGB0, ND5, *, 
			10'd51 : rdata = 48'b000111110000000001100000101000000000000000000000;
			// PEs: 63, 63 -> 
			// srcs: (1999, 49)(3) 1, (3623) 0 --> (4407) 0:NM0, ALU, *, 
			10'd52 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 63, 63 -> 63
			// srcs: (2002, 64)(1271) 0, (4407) 0 --> (5191) 0:NW5, ALU, -, NW5
			10'd53 : rdata = 48'b000100100000010100111111111000000101010000000000;
			// PEs: 56, 63 -> 
			// srcs: (2076, 34)(3140) 47, (566) 1 --> (3703) 47:PEGB0, ND6, *, 
			10'd54 : rdata = 48'b000111110000000001100000110000000000000000000000;
			// PEs: 63, 63 -> 
			// srcs: (2079, 50)(3) 1, (3703) 47 --> (4487) 47:NM0, ALU, *, 
			10'd55 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 63, 63 -> 63
			// srcs: (2082, 65)(1351) -3, (4487) 47 --> (5271) -50:NW6, ALU, -, NW6
			10'd56 : rdata = 48'b000100100000011000111111111000000101100000000000;
			// PEs: 56, 63 -> 
			// srcs: (2117, 35)(3140) 47, (607) -1 --> (3744) -47:PEGB0, ND12, *, 
			10'd57 : rdata = 48'b000111110000000001100001100000000000000000000000;
			// PEs: 63, 63 -> 
			// srcs: (2120, 51)(3) 1, (3744) -47 --> (4528) -47:NM0, ALU, *, 
			10'd58 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 63, 63 -> 63
			// srcs: (2123, 66)(1392) -2, (4528) -47 --> (5312) 45:NW12, ALU, -, NW12
			10'd59 : rdata = 48'b000100100000110000111111111000000111000000000000;
			// PEs: 56, 63 -> 63
			// srcs: (2156, 36)(3140) 47, (646) -2 --> (3783) -94:PEGB0, ND7, *, NI0
			10'd60 : rdata = 48'b000111110000000001100000111100000000000000000000;
			// PEs: 63, 62 -> 62
			// srcs: (2158, 52)(3) 1, (3782) 47 --> (4566) 47:NM0, PENB, *, PEGB6
			10'd61 : rdata = 48'b000111000000000011011111110000000000000011100000;
			// PEs: 63, 63 -> 
			// srcs: (2159, 53)(3) 1, (3783) -94 --> (4567) -94:NM0, NI0, *, 
			10'd62 : rdata = 48'b000111000000000010100000000000000000000000000000;
			// PEs: 63, 63 -> 63
			// srcs: (2162, 67)(1431) -1, (4567) -94 --> (5351) 93:NW7, ALU, -, NW7
			10'd63 : rdata = 48'b000100100000011100111111111000000101110000000000;
			// PEs: 56, 63 -> 
			// srcs: (2238, 37)(3140) 47, (728) 0 --> (3865) 0:PEGB0, ND8, *, 
			10'd64 : rdata = 48'b000111110000000001100001000000000000000000000000;
			// PEs: 63, 63 -> 
			// srcs: (2241, 54)(3) 1, (3865) 0 --> (4649) 0:NM0, ALU, *, 
			10'd65 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 63, 63 -> 63
			// srcs: (2244, 68)(1513) 1, (4649) 0 --> (5433) 1:NW8, ALU, -, NW8
			10'd66 : rdata = 48'b000100100000100000111111111000000110000000000000;
			// PEs: 56, 63 -> 
			// srcs: (2297, 38)(3140) 47, (787) 0 --> (3924) 0:PEGB0, ND13, *, 
			10'd67 : rdata = 48'b000111110000000001100001101000000000000000000000;
			// PEs: 63, 63 -> 
			// srcs: (2300, 55)(3) 1, (3924) 0 --> (4708) 0:NM0, ALU, *, 
			10'd68 : rdata = 48'b000111000000000000111111111000000000000000000000;
			// PEs: 63, 63 -> 63
			// srcs: (2303, 69)(1572) -1, (4708) 0 --> (5492) -1:NW13, ALU, -, NW13
			10'd69 : rdata = 48'b000100100000110100111111111000000111010000000000;
			default : rdata = 48'b000000000000000000000000000000000000000000000000;
		endcase
	end
end

endgenerate
/*****************************************************************************/
endmodule
