`timescale 1ns/1ps
module sigmoid#(
    parameter dataLen = 32,
	parameter indexLen =9,
	parameter fracLen = 7
)(
	input[dataLen-1:0]in,
	output[dataLen-1:0]out
);

	wire signed [dataLen - 1 : 0] in;
	reg signed [dataLen - 1 : 0] out;
	reg [indexLen - 1 :0] index;

	always @(in)
	begin
		out = 0;

		if (in < -(8 << 7)) begin
			out = 0;
		end else if (in > (8 << 7)) begin
			out = 1<<7;
		end else begin
		index[indexLen-1]	= in[dataLen-1];
		index[indexLen-2:0]	= in[fracLen+indexLen-5:fracLen-5];
		case(index)
            //
            9'd0: out = 32'b00000000000000000000000001000000;
            9'd1: out = 32'b00000000000000000000000001000000;
            9'd2: out = 32'b00000000000000000000000001000001;
            9'd3: out = 32'b00000000000000000000000001000010;
            9'd4: out = 32'b00000000000000000000000001000011;
            9'd5: out = 32'b00000000000000000000000001000100;
            9'd6: out = 32'b00000000000000000000000001000101;
            9'd7: out = 32'b00000000000000000000000001000110;
            9'd8: out = 32'b00000000000000000000000001000111;
            9'd9: out = 32'b00000000000000000000000001001000;
            9'd10: out = 32'b00000000000000000000000001001001;
            9'd11: out = 32'b00000000000000000000000001001010;
            9'd12: out = 32'b00000000000000000000000001001011;
            9'd13: out = 32'b00000000000000000000000001001100;
            9'd14: out = 32'b00000000000000000000000001001101;
            9'd15: out = 32'b00000000000000000000000001001110;
            9'd16: out = 32'b00000000000000000000000001001111;
            9'd17: out = 32'b00000000000000000000000001010000;
            9'd18: out = 32'b00000000000000000000000001010001;
            9'd19: out = 32'b00000000000000000000000001010010;
            9'd20: out = 32'b00000000000000000000000001010011;
            9'd21: out = 32'b00000000000000000000000001010100;
            9'd22: out = 32'b00000000000000000000000001010101;
            9'd23: out = 32'b00000000000000000000000001010110;
            9'd24: out = 32'b00000000000000000000000001010110;
            9'd25: out = 32'b00000000000000000000000001010111;
            9'd26: out = 32'b00000000000000000000000001011000;
            9'd27: out = 32'b00000000000000000000000001011001;
            9'd28: out = 32'b00000000000000000000000001011010;
            9'd29: out = 32'b00000000000000000000000001011011;
            9'd30: out = 32'b00000000000000000000000001011011;
            9'd31: out = 32'b00000000000000000000000001011100;
            9'd32: out = 32'b00000000000000000000000001011101;
            9'd33: out = 32'b00000000000000000000000001011110;
            9'd34: out = 32'b00000000000000000000000001011111;
            9'd35: out = 32'b00000000000000000000000001011111;
            9'd36: out = 32'b00000000000000000000000001100000;
            9'd37: out = 32'b00000000000000000000000001100001;
            9'd38: out = 32'b00000000000000000000000001100010;
            9'd39: out = 32'b00000000000000000000000001100010;
            9'd40: out = 32'b00000000000000000000000001100011;
            9'd41: out = 32'b00000000000000000000000001100100;
            9'd42: out = 32'b00000000000000000000000001100100;
            9'd43: out = 32'b00000000000000000000000001100101;
            9'd44: out = 32'b00000000000000000000000001100110;
            9'd45: out = 32'b00000000000000000000000001100110;
            9'd46: out = 32'b00000000000000000000000001100111;
            9'd47: out = 32'b00000000000000000000000001101000;
            9'd48: out = 32'b00000000000000000000000001101000;
            9'd49: out = 32'b00000000000000000000000001101001;
            9'd50: out = 32'b00000000000000000000000001101001;
            9'd51: out = 32'b00000000000000000000000001101010;
            9'd52: out = 32'b00000000000000000000000001101010;
            9'd53: out = 32'b00000000000000000000000001101011;
            9'd54: out = 32'b00000000000000000000000001101100;
            9'd55: out = 32'b00000000000000000000000001101100;
            9'd56: out = 32'b00000000000000000000000001101101;
            9'd57: out = 32'b00000000000000000000000001101101;
            9'd58: out = 32'b00000000000000000000000001101110;
            9'd59: out = 32'b00000000000000000000000001101110;
            9'd60: out = 32'b00000000000000000000000001101110;
            9'd61: out = 32'b00000000000000000000000001101111;
            9'd62: out = 32'b00000000000000000000000001101111;
            9'd63: out = 32'b00000000000000000000000001110000;
            9'd64: out = 32'b00000000000000000000000001110000;
            9'd65: out = 32'b00000000000000000000000001110001;
            9'd66: out = 32'b00000000000000000000000001110001;
            9'd67: out = 32'b00000000000000000000000001110001;
            9'd68: out = 32'b00000000000000000000000001110010;
            9'd69: out = 32'b00000000000000000000000001110010;
            9'd70: out = 32'b00000000000000000000000001110011;
            9'd71: out = 32'b00000000000000000000000001110011;
            9'd72: out = 32'b00000000000000000000000001110011;
            9'd73: out = 32'b00000000000000000000000001110100;
            9'd74: out = 32'b00000000000000000000000001110100;
            9'd75: out = 32'b00000000000000000000000001110100;
            9'd76: out = 32'b00000000000000000000000001110101;
            9'd77: out = 32'b00000000000000000000000001110101;
            9'd78: out = 32'b00000000000000000000000001110101;
            9'd79: out = 32'b00000000000000000000000001110110;
            9'd80: out = 32'b00000000000000000000000001110110;
            9'd81: out = 32'b00000000000000000000000001110110;
            9'd82: out = 32'b00000000000000000000000001110110;
            9'd83: out = 32'b00000000000000000000000001110111;
            9'd84: out = 32'b00000000000000000000000001110111;
            9'd85: out = 32'b00000000000000000000000001110111;
            9'd86: out = 32'b00000000000000000000000001110111;
            9'd87: out = 32'b00000000000000000000000001111000;
            9'd88: out = 32'b00000000000000000000000001111000;
            9'd89: out = 32'b00000000000000000000000001111000;
            9'd90: out = 32'b00000000000000000000000001111000;
            9'd91: out = 32'b00000000000000000000000001111000;
            9'd92: out = 32'b00000000000000000000000001111001;
            9'd93: out = 32'b00000000000000000000000001111001;
            9'd94: out = 32'b00000000000000000000000001111001;
            9'd95: out = 32'b00000000000000000000000001111001;
            9'd96: out = 32'b00000000000000000000000001111001;
            9'd97: out = 32'b00000000000000000000000001111010;
            9'd98: out = 32'b00000000000000000000000001111010;
            9'd99: out = 32'b00000000000000000000000001111010;
            9'd100: out = 32'b00000000000000000000000001111010;
            9'd101: out = 32'b00000000000000000000000001111010;
            9'd102: out = 32'b00000000000000000000000001111010;
            9'd103: out = 32'b00000000000000000000000001111011;
            9'd104: out = 32'b00000000000000000000000001111011;
            9'd105: out = 32'b00000000000000000000000001111011;
            9'd106: out = 32'b00000000000000000000000001111011;
            9'd107: out = 32'b00000000000000000000000001111011;
            9'd108: out = 32'b00000000000000000000000001111011;
            9'd109: out = 32'b00000000000000000000000001111011;
            9'd110: out = 32'b00000000000000000000000001111100;
            9'd111: out = 32'b00000000000000000000000001111100;
            9'd112: out = 32'b00000000000000000000000001111100;
            9'd113: out = 32'b00000000000000000000000001111100;
            9'd114: out = 32'b00000000000000000000000001111100;
            9'd115: out = 32'b00000000000000000000000001111100;
            9'd116: out = 32'b00000000000000000000000001111100;
            9'd117: out = 32'b00000000000000000000000001111100;
            9'd118: out = 32'b00000000000000000000000001111100;
            9'd119: out = 32'b00000000000000000000000001111100;
            9'd120: out = 32'b00000000000000000000000001111101;
            9'd121: out = 32'b00000000000000000000000001111101;
            9'd122: out = 32'b00000000000000000000000001111101;
            9'd123: out = 32'b00000000000000000000000001111101;
            9'd124: out = 32'b00000000000000000000000001111101;
            9'd125: out = 32'b00000000000000000000000001111101;
            9'd126: out = 32'b00000000000000000000000001111101;
            9'd127: out = 32'b00000000000000000000000001111101;
            9'd128: out = 32'b00000000000000000000000001111101;
            9'd129: out = 32'b00000000000000000000000001111101;
            9'd130: out = 32'b00000000000000000000000001111101;
            9'd131: out = 32'b00000000000000000000000001111101;
            9'd132: out = 32'b00000000000000000000000001111101;
            9'd133: out = 32'b00000000000000000000000001111110;
            9'd134: out = 32'b00000000000000000000000001111110;
            9'd135: out = 32'b00000000000000000000000001111110;
            9'd136: out = 32'b00000000000000000000000001111110;
            9'd137: out = 32'b00000000000000000000000001111110;
            9'd138: out = 32'b00000000000000000000000001111110;
            9'd139: out = 32'b00000000000000000000000001111110;
            9'd140: out = 32'b00000000000000000000000001111110;
            9'd141: out = 32'b00000000000000000000000001111110;
            9'd142: out = 32'b00000000000000000000000001111110;
            9'd143: out = 32'b00000000000000000000000001111110;
            9'd144: out = 32'b00000000000000000000000001111110;
            9'd145: out = 32'b00000000000000000000000001111110;
            9'd146: out = 32'b00000000000000000000000001111110;
            9'd147: out = 32'b00000000000000000000000001111110;
            9'd148: out = 32'b00000000000000000000000001111110;
            9'd149: out = 32'b00000000000000000000000001111110;
            9'd150: out = 32'b00000000000000000000000001111110;
            9'd151: out = 32'b00000000000000000000000001111110;
            9'd152: out = 32'b00000000000000000000000001111110;
            9'd153: out = 32'b00000000000000000000000001111110;
            9'd154: out = 32'b00000000000000000000000001111110;
            9'd155: out = 32'b00000000000000000000000001111110;
            9'd156: out = 32'b00000000000000000000000001111111;
            9'd157: out = 32'b00000000000000000000000001111111;
            9'd158: out = 32'b00000000000000000000000001111111;
            9'd159: out = 32'b00000000000000000000000001111111;
            9'd160: out = 32'b00000000000000000000000001111111;
            9'd161: out = 32'b00000000000000000000000001111111;
            9'd162: out = 32'b00000000000000000000000001111111;
            9'd163: out = 32'b00000000000000000000000001111111;
            9'd164: out = 32'b00000000000000000000000001111111;
            9'd165: out = 32'b00000000000000000000000001111111;
            9'd166: out = 32'b00000000000000000000000001111111;
            9'd167: out = 32'b00000000000000000000000001111111;
            9'd168: out = 32'b00000000000000000000000001111111;
            9'd169: out = 32'b00000000000000000000000001111111;
            9'd170: out = 32'b00000000000000000000000001111111;
            9'd171: out = 32'b00000000000000000000000001111111;
            9'd172: out = 32'b00000000000000000000000001111111;
            9'd173: out = 32'b00000000000000000000000001111111;
            9'd174: out = 32'b00000000000000000000000001111111;
            9'd175: out = 32'b00000000000000000000000001111111;
            9'd176: out = 32'b00000000000000000000000001111111;
            9'd177: out = 32'b00000000000000000000000001111111;
            9'd178: out = 32'b00000000000000000000000001111111;
            9'd179: out = 32'b00000000000000000000000001111111;
            9'd180: out = 32'b00000000000000000000000001111111;
            9'd181: out = 32'b00000000000000000000000001111111;
            9'd182: out = 32'b00000000000000000000000001111111;
            9'd183: out = 32'b00000000000000000000000001111111;
            9'd184: out = 32'b00000000000000000000000001111111;
            9'd185: out = 32'b00000000000000000000000001111111;
            9'd186: out = 32'b00000000000000000000000001111111;
            9'd187: out = 32'b00000000000000000000000001111111;
            9'd188: out = 32'b00000000000000000000000001111111;
            9'd189: out = 32'b00000000000000000000000001111111;
            9'd190: out = 32'b00000000000000000000000001111111;
            9'd191: out = 32'b00000000000000000000000001111111;
            9'd192: out = 32'b00000000000000000000000001111111;
            9'd193: out = 32'b00000000000000000000000001111111;
            9'd194: out = 32'b00000000000000000000000001111111;
            9'd195: out = 32'b00000000000000000000000001111111;
            9'd196: out = 32'b00000000000000000000000001111111;
            9'd197: out = 32'b00000000000000000000000001111111;
            9'd198: out = 32'b00000000000000000000000001111111;
            9'd199: out = 32'b00000000000000000000000001111111;
            9'd200: out = 32'b00000000000000000000000001111111;
            9'd201: out = 32'b00000000000000000000000001111111;
            9'd202: out = 32'b00000000000000000000000001111111;
            9'd203: out = 32'b00000000000000000000000001111111;
            9'd204: out = 32'b00000000000000000000000001111111;
            9'd205: out = 32'b00000000000000000000000001111111;
            9'd206: out = 32'b00000000000000000000000001111111;
            9'd207: out = 32'b00000000000000000000000001111111;
            9'd208: out = 32'b00000000000000000000000001111111;
            9'd209: out = 32'b00000000000000000000000001111111;
            9'd210: out = 32'b00000000000000000000000001111111;
            9'd211: out = 32'b00000000000000000000000001111111;
            9'd212: out = 32'b00000000000000000000000001111111;
            9'd213: out = 32'b00000000000000000000000001111111;
            9'd214: out = 32'b00000000000000000000000001111111;
            9'd215: out = 32'b00000000000000000000000001111111;
            9'd216: out = 32'b00000000000000000000000001111111;
            9'd217: out = 32'b00000000000000000000000001111111;
            9'd218: out = 32'b00000000000000000000000001111111;
            9'd219: out = 32'b00000000000000000000000001111111;
            9'd220: out = 32'b00000000000000000000000001111111;
            9'd221: out = 32'b00000000000000000000000001111111;
            9'd222: out = 32'b00000000000000000000000001111111;
            9'd223: out = 32'b00000000000000000000000001111111;
            9'd224: out = 32'b00000000000000000000000001111111;
            9'd225: out = 32'b00000000000000000000000001111111;
            9'd226: out = 32'b00000000000000000000000001111111;
            9'd227: out = 32'b00000000000000000000000001111111;
            9'd228: out = 32'b00000000000000000000000001111111;
            9'd229: out = 32'b00000000000000000000000001111111;
            9'd230: out = 32'b00000000000000000000000001111111;
            9'd231: out = 32'b00000000000000000000000001111111;
            9'd232: out = 32'b00000000000000000000000001111111;
            9'd233: out = 32'b00000000000000000000000001111111;
            9'd234: out = 32'b00000000000000000000000001111111;
            9'd235: out = 32'b00000000000000000000000001111111;
            9'd236: out = 32'b00000000000000000000000001111111;
            9'd237: out = 32'b00000000000000000000000001111111;
            9'd238: out = 32'b00000000000000000000000001111111;
            9'd239: out = 32'b00000000000000000000000001111111;
            9'd240: out = 32'b00000000000000000000000001111111;
            9'd241: out = 32'b00000000000000000000000001111111;
            9'd242: out = 32'b00000000000000000000000001111111;
            9'd243: out = 32'b00000000000000000000000001111111;
            9'd244: out = 32'b00000000000000000000000001111111;
            9'd245: out = 32'b00000000000000000000000001111111;
            9'd246: out = 32'b00000000000000000000000001111111;
            9'd247: out = 32'b00000000000000000000000001111111;
            9'd248: out = 32'b00000000000000000000000001111111;
            9'd249: out = 32'b00000000000000000000000001111111;
            9'd250: out = 32'b00000000000000000000000001111111;
            9'd251: out = 32'b00000000000000000000000001111111;
            9'd252: out = 32'b00000000000000000000000001111111;
            9'd253: out = 32'b00000000000000000000000001111111;
            9'd254: out = 32'b00000000000000000000000001111111;
            9'd255: out = 32'b00000000000000000000000001111111;
            9'd257: out = 32'b00000000000000000000000000000000;
            9'd258: out = 32'b00000000000000000000000000000000;
            9'd259: out = 32'b00000000000000000000000000000000;
            9'd260: out = 32'b00000000000000000000000000000000;
            9'd261: out = 32'b00000000000000000000000000000000;
            9'd262: out = 32'b00000000000000000000000000000000;
            9'd263: out = 32'b00000000000000000000000000000000;
            9'd264: out = 32'b00000000000000000000000000000000;
            9'd265: out = 32'b00000000000000000000000000000000;
            9'd266: out = 32'b00000000000000000000000000000000;
            9'd267: out = 32'b00000000000000000000000000000000;
            9'd268: out = 32'b00000000000000000000000000000000;
            9'd269: out = 32'b00000000000000000000000000000000;
            9'd270: out = 32'b00000000000000000000000000000000;
            9'd271: out = 32'b00000000000000000000000000000000;
            9'd272: out = 32'b00000000000000000000000000000000;
            9'd273: out = 32'b00000000000000000000000000000000;
            9'd274: out = 32'b00000000000000000000000000000000;
            9'd275: out = 32'b00000000000000000000000000000000;
            9'd276: out = 32'b00000000000000000000000000000000;
            9'd277: out = 32'b00000000000000000000000000000000;
            9'd278: out = 32'b00000000000000000000000000000000;
            9'd279: out = 32'b00000000000000000000000000000000;
            9'd280: out = 32'b00000000000000000000000000000000;
            9'd281: out = 32'b00000000000000000000000000000000;
            9'd282: out = 32'b00000000000000000000000000000000;
            9'd283: out = 32'b00000000000000000000000000000000;
            9'd284: out = 32'b00000000000000000000000000000000;
            9'd285: out = 32'b00000000000000000000000000000000;
            9'd286: out = 32'b00000000000000000000000000000000;
            9'd287: out = 32'b00000000000000000000000000000000;
            9'd288: out = 32'b00000000000000000000000000000000;
            9'd289: out = 32'b00000000000000000000000000000000;
            9'd290: out = 32'b00000000000000000000000000000000;
            9'd291: out = 32'b00000000000000000000000000000000;
            9'd292: out = 32'b00000000000000000000000000000000;
            9'd293: out = 32'b00000000000000000000000000000000;
            9'd294: out = 32'b00000000000000000000000000000000;
            9'd295: out = 32'b00000000000000000000000000000000;
            9'd296: out = 32'b00000000000000000000000000000000;
            9'd297: out = 32'b00000000000000000000000000000000;
            9'd298: out = 32'b00000000000000000000000000000000;
            9'd299: out = 32'b00000000000000000000000000000000;
            9'd300: out = 32'b00000000000000000000000000000000;
            9'd301: out = 32'b00000000000000000000000000000000;
            9'd302: out = 32'b00000000000000000000000000000000;
            9'd303: out = 32'b00000000000000000000000000000000;
            9'd304: out = 32'b00000000000000000000000000000000;
            9'd305: out = 32'b00000000000000000000000000000000;
            9'd306: out = 32'b00000000000000000000000000000000;
            9'd307: out = 32'b00000000000000000000000000000000;
            9'd308: out = 32'b00000000000000000000000000000000;
            9'd309: out = 32'b00000000000000000000000000000000;
            9'd310: out = 32'b00000000000000000000000000000000;
            9'd311: out = 32'b00000000000000000000000000000000;
            9'd312: out = 32'b00000000000000000000000000000000;
            9'd313: out = 32'b00000000000000000000000000000000;
            9'd314: out = 32'b00000000000000000000000000000000;
            9'd315: out = 32'b00000000000000000000000000000000;
            9'd316: out = 32'b00000000000000000000000000000000;
            9'd317: out = 32'b00000000000000000000000000000000;
            9'd318: out = 32'b00000000000000000000000000000000;
            9'd319: out = 32'b00000000000000000000000000000000;
            9'd320: out = 32'b00000000000000000000000000000000;
            9'd321: out = 32'b00000000000000000000000000000000;
            9'd322: out = 32'b00000000000000000000000000000000;
            9'd323: out = 32'b00000000000000000000000000000000;
            9'd324: out = 32'b00000000000000000000000000000000;
            9'd325: out = 32'b00000000000000000000000000000000;
            9'd326: out = 32'b00000000000000000000000000000000;
            9'd327: out = 32'b00000000000000000000000000000000;
            9'd328: out = 32'b00000000000000000000000000000000;
            9'd329: out = 32'b00000000000000000000000000000000;
            9'd330: out = 32'b00000000000000000000000000000000;
            9'd331: out = 32'b00000000000000000000000000000000;
            9'd332: out = 32'b00000000000000000000000000000000;
            9'd333: out = 32'b00000000000000000000000000000000;
            9'd334: out = 32'b00000000000000000000000000000000;
            9'd335: out = 32'b00000000000000000000000000000000;
            9'd336: out = 32'b00000000000000000000000000000000;
            9'd337: out = 32'b00000000000000000000000000000000;
            9'd338: out = 32'b00000000000000000000000000000000;
            9'd339: out = 32'b00000000000000000000000000000000;
            9'd340: out = 32'b00000000000000000000000000000000;
            9'd341: out = 32'b00000000000000000000000000000000;
            9'd342: out = 32'b00000000000000000000000000000000;
            9'd343: out = 32'b00000000000000000000000000000000;
            9'd344: out = 32'b00000000000000000000000000000000;
            9'd345: out = 32'b00000000000000000000000000000000;
            9'd346: out = 32'b00000000000000000000000000000000;
            9'd347: out = 32'b00000000000000000000000000000000;
            9'd348: out = 32'b00000000000000000000000000000000;
            9'd349: out = 32'b00000000000000000000000000000000;
            9'd350: out = 32'b00000000000000000000000000000000;
            9'd351: out = 32'b00000000000000000000000000000000;
            9'd352: out = 32'b00000000000000000000000000000000;
            9'd353: out = 32'b00000000000000000000000000000000;
            9'd354: out = 32'b00000000000000000000000000000000;
            9'd355: out = 32'b00000000000000000000000000000000;
            9'd356: out = 32'b00000000000000000000000000000000;
            9'd357: out = 32'b00000000000000000000000000000001;
            9'd358: out = 32'b00000000000000000000000000000001;
            9'd359: out = 32'b00000000000000000000000000000001;
            9'd360: out = 32'b00000000000000000000000000000001;
            9'd361: out = 32'b00000000000000000000000000000001;
            9'd362: out = 32'b00000000000000000000000000000001;
            9'd363: out = 32'b00000000000000000000000000000001;
            9'd364: out = 32'b00000000000000000000000000000001;
            9'd365: out = 32'b00000000000000000000000000000001;
            9'd366: out = 32'b00000000000000000000000000000001;
            9'd367: out = 32'b00000000000000000000000000000001;
            9'd368: out = 32'b00000000000000000000000000000001;
            9'd369: out = 32'b00000000000000000000000000000001;
            9'd370: out = 32'b00000000000000000000000000000001;
            9'd371: out = 32'b00000000000000000000000000000001;
            9'd372: out = 32'b00000000000000000000000000000001;
            9'd373: out = 32'b00000000000000000000000000000001;
            9'd374: out = 32'b00000000000000000000000000000001;
            9'd375: out = 32'b00000000000000000000000000000001;
            9'd376: out = 32'b00000000000000000000000000000001;
            9'd377: out = 32'b00000000000000000000000000000001;
            9'd378: out = 32'b00000000000000000000000000000001;
            9'd379: out = 32'b00000000000000000000000000000001;
            9'd380: out = 32'b00000000000000000000000000000010;
            9'd381: out = 32'b00000000000000000000000000000010;
            9'd382: out = 32'b00000000000000000000000000000010;
            9'd383: out = 32'b00000000000000000000000000000010;
            9'd384: out = 32'b00000000000000000000000000000010;
            9'd385: out = 32'b00000000000000000000000000000010;
            9'd386: out = 32'b00000000000000000000000000000010;
            9'd387: out = 32'b00000000000000000000000000000010;
            9'd388: out = 32'b00000000000000000000000000000010;
            9'd389: out = 32'b00000000000000000000000000000010;
            9'd390: out = 32'b00000000000000000000000000000010;
            9'd391: out = 32'b00000000000000000000000000000010;
            9'd392: out = 32'b00000000000000000000000000000010;
            9'd393: out = 32'b00000000000000000000000000000011;
            9'd394: out = 32'b00000000000000000000000000000011;
            9'd395: out = 32'b00000000000000000000000000000011;
            9'd396: out = 32'b00000000000000000000000000000011;
            9'd397: out = 32'b00000000000000000000000000000011;
            9'd398: out = 32'b00000000000000000000000000000011;
            9'd399: out = 32'b00000000000000000000000000000011;
            9'd400: out = 32'b00000000000000000000000000000011;
            9'd401: out = 32'b00000000000000000000000000000011;
            9'd402: out = 32'b00000000000000000000000000000011;
            9'd403: out = 32'b00000000000000000000000000000100;
            9'd404: out = 32'b00000000000000000000000000000100;
            9'd405: out = 32'b00000000000000000000000000000100;
            9'd406: out = 32'b00000000000000000000000000000100;
            9'd407: out = 32'b00000000000000000000000000000100;
            9'd408: out = 32'b00000000000000000000000000000100;
            9'd409: out = 32'b00000000000000000000000000000100;
            9'd410: out = 32'b00000000000000000000000000000101;
            9'd411: out = 32'b00000000000000000000000000000101;
            9'd412: out = 32'b00000000000000000000000000000101;
            9'd413: out = 32'b00000000000000000000000000000101;
            9'd414: out = 32'b00000000000000000000000000000101;
            9'd415: out = 32'b00000000000000000000000000000101;
            9'd416: out = 32'b00000000000000000000000000000110;
            9'd417: out = 32'b00000000000000000000000000000110;
            9'd418: out = 32'b00000000000000000000000000000110;
            9'd419: out = 32'b00000000000000000000000000000110;
            9'd420: out = 32'b00000000000000000000000000000110;
            9'd421: out = 32'b00000000000000000000000000000111;
            9'd422: out = 32'b00000000000000000000000000000111;
            9'd423: out = 32'b00000000000000000000000000000111;
            9'd424: out = 32'b00000000000000000000000000000111;
            9'd425: out = 32'b00000000000000000000000000000111;
            9'd426: out = 32'b00000000000000000000000000001000;
            9'd427: out = 32'b00000000000000000000000000001000;
            9'd428: out = 32'b00000000000000000000000000001000;
            9'd429: out = 32'b00000000000000000000000000001000;
            9'd430: out = 32'b00000000000000000000000000001001;
            9'd431: out = 32'b00000000000000000000000000001001;
            9'd432: out = 32'b00000000000000000000000000001001;
            9'd433: out = 32'b00000000000000000000000000001001;
            9'd434: out = 32'b00000000000000000000000000001010;
            9'd435: out = 32'b00000000000000000000000000001010;
            9'd436: out = 32'b00000000000000000000000000001010;
            9'd437: out = 32'b00000000000000000000000000001011;
            9'd438: out = 32'b00000000000000000000000000001011;
            9'd439: out = 32'b00000000000000000000000000001011;
            9'd440: out = 32'b00000000000000000000000000001100;
            9'd441: out = 32'b00000000000000000000000000001100;
            9'd442: out = 32'b00000000000000000000000000001100;
            9'd443: out = 32'b00000000000000000000000000001101;
            9'd444: out = 32'b00000000000000000000000000001101;
            9'd445: out = 32'b00000000000000000000000000001110;
            9'd446: out = 32'b00000000000000000000000000001110;
            9'd447: out = 32'b00000000000000000000000000001110;
            9'd448: out = 32'b00000000000000000000000000001111;
            9'd449: out = 32'b00000000000000000000000000001111;
            9'd450: out = 32'b00000000000000000000000000010000;
            9'd451: out = 32'b00000000000000000000000000010000;
            9'd452: out = 32'b00000000000000000000000000010001;
            9'd453: out = 32'b00000000000000000000000000010001;
            9'd454: out = 32'b00000000000000000000000000010001;
            9'd455: out = 32'b00000000000000000000000000010010;
            9'd456: out = 32'b00000000000000000000000000010010;
            9'd457: out = 32'b00000000000000000000000000010011;
            9'd458: out = 32'b00000000000000000000000000010011;
            9'd459: out = 32'b00000000000000000000000000010100;
            9'd460: out = 32'b00000000000000000000000000010101;
            9'd461: out = 32'b00000000000000000000000000010101;
            9'd462: out = 32'b00000000000000000000000000010110;
            9'd463: out = 32'b00000000000000000000000000010110;
            9'd464: out = 32'b00000000000000000000000000010111;
            9'd465: out = 32'b00000000000000000000000000010111;
            9'd466: out = 32'b00000000000000000000000000011000;
            9'd467: out = 32'b00000000000000000000000000011001;
            9'd468: out = 32'b00000000000000000000000000011001;
            9'd469: out = 32'b00000000000000000000000000011010;
            9'd470: out = 32'b00000000000000000000000000011011;
            9'd471: out = 32'b00000000000000000000000000011011;
            9'd472: out = 32'b00000000000000000000000000011100;
            9'd473: out = 32'b00000000000000000000000000011101;
            9'd474: out = 32'b00000000000000000000000000011101;
            9'd475: out = 32'b00000000000000000000000000011110;
            9'd476: out = 32'b00000000000000000000000000011111;
            9'd477: out = 32'b00000000000000000000000000100000;
            9'd478: out = 32'b00000000000000000000000000100000;
            9'd479: out = 32'b00000000000000000000000000100001;
            9'd480: out = 32'b00000000000000000000000000100010;
            9'd481: out = 32'b00000000000000000000000000100011;
            9'd482: out = 32'b00000000000000000000000000100100;
            9'd483: out = 32'b00000000000000000000000000100100;
            9'd484: out = 32'b00000000000000000000000000100101;
            9'd485: out = 32'b00000000000000000000000000100110;
            9'd486: out = 32'b00000000000000000000000000100111;
            9'd487: out = 32'b00000000000000000000000000101000;
            9'd488: out = 32'b00000000000000000000000000101001;
            9'd489: out = 32'b00000000000000000000000000101001;
            9'd490: out = 32'b00000000000000000000000000101010;
            9'd491: out = 32'b00000000000000000000000000101011;
            9'd492: out = 32'b00000000000000000000000000101100;
            9'd493: out = 32'b00000000000000000000000000101101;
            9'd494: out = 32'b00000000000000000000000000101110;
            9'd495: out = 32'b00000000000000000000000000101111;
            9'd496: out = 32'b00000000000000000000000000110000;
            9'd497: out = 32'b00000000000000000000000000110001;
            9'd498: out = 32'b00000000000000000000000000110010;
            9'd499: out = 32'b00000000000000000000000000110011;
            9'd500: out = 32'b00000000000000000000000000110100;
            9'd501: out = 32'b00000000000000000000000000110101;
            9'd502: out = 32'b00000000000000000000000000110110;
            9'd503: out = 32'b00000000000000000000000000110111;
            9'd504: out = 32'b00000000000000000000000000111000;
            9'd505: out = 32'b00000000000000000000000000111001;
            9'd506: out = 32'b00000000000000000000000000111010;
            9'd507: out = 32'b00000000000000000000000000111011;
            9'd508: out = 32'b00000000000000000000000000111100;
            9'd509: out = 32'b00000000000000000000000000111101;
            9'd510: out = 32'b00000000000000000000000000111110;
            9'd511: out = 32'b00000000000000000000000000111111;
		endcase
		end
	end

endmodule
  
