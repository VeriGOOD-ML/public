
`timescale 1ns/1ps
module instruction_memory #(
    parameter integer addrLen = 5,
    parameter integer dataLen = 32,
    parameter integer peId  = 1
)(
    input clk,
    input rstn,
    
    input stall,
    input start,
    input restart,
    
    output reg [dataLen - 1: 0] data_out
);
//--------------------------------------------------------------------------------------
//reg [dataLen - 1: 0] mem  [0: (1 << addrLen) - 1];
reg [addrLen-1:0]        address;
reg enable;
reg [dataLen - 1: 0] rdata;
wire end_of_instruction;
always @(posedge clk or negedge rstn)
    if(~rstn)
        enable <= 1'b0;
    else if(start)
        enable <= 1'b1;
    else if(end_of_instruction)
       enable <= 1'b0;
always @(posedge clk or negedge rstn) begin
    if(~rstn)
        address <= {addrLen{1'b0}};
    else begin
        if(end_of_instruction)
            address <= {addrLen{1'b0}};
        else if(~stall && enable )
            address <= address + {{addrLen-1{1'b0}},1'b1};   
    end     
end
always @(posedge clk or negedge rstn) begin
    if(~rstn)
        data_out <= {1'b1,{dataLen-1{1'b0}}};
    else if((~stall && enable && ~end_of_instruction)||(end_of_instruction && start))
       data_out <= rdata;
end
    
assign end_of_instruction = (data_out[dataLen-1:dataLen-5] == 5'b0);
/****************************************************************************/
generate
if(peId == 0) begin
	always @(*) begin
		case(address)
			// PEs: 7 -> 8
			// srcs: (3, 0)(120) 72 --> (120) 72:PENB, pass, PUNB
			6'd0 : rdata = 41'b11000110111111100000000000000001000000000;
			// PEs: 56 -> 0
			// srcs: (8, 3)(146) 48 --> (146) 48:PUNB, pass, NI0
			6'd1 : rdata = 41'b11000110111111110000000000010000000000000;
			// PEs: 6 -> 16
			// srcs: (9, 1)(170) 19 --> (170) 19:PEGB6, pass, PUGB2
			6'd2 : rdata = 41'b11000111000011000000000000000000000001010;
			// PEs: 24 -> 1
			// srcs: (11, 2)(196) 7 --> (196) 7:PUGB3, pass, PENB
			6'd3 : rdata = 41'b11000111000001110000000000000000100000000;
			// PEs: 1 -> 48
			// srcs: (17, 5)(169) 74 --> (169) 74:PEGB1, pass, PUGB6
			6'd4 : rdata = 41'b11000111000000100000000000000000000001110;
			// PEs: 0 -> 1
			// srcs: (18, 4)(146) 48 --> (146) 48:NI0, pass, PENB
			6'd5 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 1 -> 8
			// srcs: (25, 6)(197) 55 --> (197) 55:PEGB1, pass, PUNB
			6'd6 : rdata = 41'b11000111000000100000000000000001000000000;
			// PEs: 40 -> 0
			// srcs: (30, 7)(211) 82 --> (211) 82:PUGB5, pass, NI0
			6'd7 : rdata = 41'b11000111000010110000000000010000000000000;
			// PEs: 56 -> 1
			// srcs: (41, 8)(216) 112 --> (216) 112:PUNB, pass, PENB
			6'd8 : rdata = 41'b11000110111111110000000000000000100000000;
			// PEs: 0 -> 1
			// srcs: (51, 9)(211) 82 --> (211) 82:NI0, pass, PENB
			6'd9 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 1 -> 24
			// srcs: (58, 10)(217) 194 --> (217) 194:PEGB1, pass, PUGB3
			6'd10 : rdata = 41'b11000111000000100000000000000000000001011;
			// PEs: 32 -> 1
			// srcs: (105, 11)(221) -3 --> (221) -3:PUGB4, pass, PENB
			6'd11 : rdata = 41'b11000111000010010000000000000000100000000;
			// PEs: 32 -> 2
			// srcs: (109, 12)(221) -3 --> (221) -3:PUGB4, pass, PEGB2
			6'd12 : rdata = 41'b11000111000010010000000000000000010100000;
			// PEs: 32 -> 3
			// srcs: (110, 13)(221) -3 --> (221) -3:PUGB4, pass, PEGB3
			6'd13 : rdata = 41'b11000111000010010000000000000000010110000;
			// PEs: 32 -> 4
			// srcs: (111, 14)(221) -3 --> (221) -3:PUGB4, pass, PEGB4
			6'd14 : rdata = 41'b11000111000010010000000000000000011000000;
			// PEs: 32 -> 5
			// srcs: (112, 15)(221) -3 --> (221) -3:PUGB4, pass, PEGB5
			6'd15 : rdata = 41'b11000111000010010000000000000000011010000;
			// PEs: 32 -> 6
			// srcs: (113, 16)(221) -3 --> (221) -3:PUGB4, pass, PEGB6
			6'd16 : rdata = 41'b11000111000010010000000000000000011100000;
			// PEs: 32 -> 7
			// srcs: (115, 17)(221) -3 --> (221) -3:PUGB4, pass, PEGB7
			6'd17 : rdata = 41'b11000111000010010000000000000000011110000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 1) begin
	always @(*) begin
		case(address)
			// PEs: 1, 1 -> 2
			// srcs: (1, 0)(4) 2, (59) 4 --> (113) 8:ND0, NW0, *, PENB
			6'd0 : rdata = 41'b00011011000000000100000000000000100000000;
			// PEs: 4 -> 
			// srcs: (9, 1)(168) 21 --> (168) 21:PEGB4, pass, 
			6'd1 : rdata = 41'b11000111000010000000000000000000000000000;
			// PEs: 2, 1 -> 0
			// srcs: (12, 2)(167) 53, (168) 21 --> (169) 74:PEGB2, ALU, +, PEGB0
			6'd2 : rdata = 41'b00001111000001000011111111100000010000000;
			// PEs: 0 -> 
			// srcs: (13, 3)(196) 7 --> (196) 7:PENB, pass, 
			6'd3 : rdata = 41'b11000110111111100000000000000000000000000;
			// PEs: 1, 0 -> 0
			// srcs: (20, 4)(196) 7, (146) 48 --> (197) 55:ALU, PENB, +, PEGB0
			6'd4 : rdata = 41'b00001001111111111101111111000000010000000;
			// PEs: 0 -> 
			// srcs: (43, 5)(216) 112 --> (216) 112:PENB, pass, 
			6'd5 : rdata = 41'b11000110111111100000000000000000000000000;
			// PEs: 0, 1 -> 0
			// srcs: (53, 6)(211) 82, (216) 112 --> (217) 194:PENB, ALU, +, PEGB0
			6'd6 : rdata = 41'b00001110111111100011111111100000010000000;
			// PEs: 0, 1 -> 2
			// srcs: (108, 7)(221) -3, (4) 2 --> (222) -6:PENB, ND0, *, PENB
			6'd7 : rdata = 41'b00011110111111100110000000000000100000000;
			// PEs: 1, 2 -> 1
			// srcs: (117, 8)(59) 4, (276) -6 --> (330) 10:NW0, PEGB2, -, NW0
			6'd8 : rdata = 41'b00010010000000001110000010000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 2) begin
	always @(*) begin
		case(address)
			// PEs: 2, 2 -> 
			// srcs: (1, 0)(5) 9, (60) 5 --> (114) 45:ND0, NW0, *, 
			6'd0 : rdata = 41'b00011011000000000100000000000000000000000;
			// PEs: 1, 2 -> 1
			// srcs: (4, 1)(113) 8, (114) 45 --> (167) 53:PENB, ALU, +, PEGB1
			6'd1 : rdata = 41'b00001110111111100011111111100000010010000;
			// PEs: 2, 1 -> 1
			// srcs: (111, 3)(3) 1, (222) -6 --> (276) -6:NM0, PENB, *, PEGB1
			6'd2 : rdata = 41'b00011100000000001101111111000000010010000;
			// PEs: 0, 2 -> 3
			// srcs: (114, 2)(221) -3, (5) 9 --> (223) -27:PEGB0, ND0, *, PENB
			6'd3 : rdata = 41'b00011111000000000110000000000000100000000;
			// PEs: 2, 3 -> 2
			// srcs: (123, 4)(60) 5, (277) -27 --> (331) 32:NW0, PEGB3, -, NW0
			6'd4 : rdata = 41'b00010010000000001110000011000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 3) begin
	always @(*) begin
		case(address)
			// PEs: 3, 3 -> 4
			// srcs: (1, 0)(6) 6, (61) 1 --> (115) 6:ND0, NW0, *, PENB
			6'd0 : rdata = 41'b00011011000000000100000000000000100000000;
			// PEs: 0, 3 -> 3
			// srcs: (115, 1)(221) -3, (6) 6 --> (224) -18:PEGB0, ND0, *, NI0
			6'd1 : rdata = 41'b00011111000000000110000000010000000000000;
			// PEs: 3, 2 -> 2
			// srcs: (117, 2)(3) 1, (223) -27 --> (277) -27:NM0, PENB, *, PEGB2
			6'd2 : rdata = 41'b00011100000000001101111111000000010100000;
			// PEs: 3, 3 -> 
			// srcs: (118, 3)(3) 1, (224) -18 --> (278) -18:NM0, NI0, *, 
			6'd3 : rdata = 41'b00011100000000001010000000000000000000000;
			// PEs: 3, 3 -> 3
			// srcs: (121, 4)(61) 1, (278) -18 --> (332) 19:NW0, ALU, -, NW0
			6'd4 : rdata = 41'b00010010000000000011111111100100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 4) begin
	always @(*) begin
		case(address)
			// PEs: 4, 4 -> 
			// srcs: (1, 0)(7) 3, (62) 5 --> (116) 15:ND0, NW0, *, 
			6'd0 : rdata = 41'b00011011000000000100000000000000000000000;
			// PEs: 3, 4 -> 1
			// srcs: (4, 1)(115) 6, (116) 15 --> (168) 21:PENB, ALU, +, PEGB1
			6'd1 : rdata = 41'b00001110111111100011111111100000010010000;
			// PEs: 0, 4 -> 5
			// srcs: (116, 2)(221) -3, (7) 3 --> (225) -9:PEGB0, ND0, *, PENB
			6'd2 : rdata = 41'b00011111000000000110000000000000100000000;
			// PEs: 4, 5 -> 4
			// srcs: (125, 3)(62) 5, (279) -9 --> (333) 14:NW0, PEGB5, -, NW0
			6'd3 : rdata = 41'b00010010000000001110000101000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 5) begin
	always @(*) begin
		case(address)
			// PEs: 5, 5 -> 6
			// srcs: (1, 0)(8) 2, (63) 6 --> (117) 12:ND0, NW0, *, PENB
			6'd0 : rdata = 41'b00011011000000000100000000000000100000000;
			// PEs: 0, 5 -> 5
			// srcs: (117, 1)(221) -3, (8) 2 --> (226) -6:PEGB0, ND0, *, NI0
			6'd1 : rdata = 41'b00011111000000000110000000010000000000000;
			// PEs: 5, 4 -> 4
			// srcs: (119, 2)(3) 1, (225) -9 --> (279) -9:NM0, PENB, *, PEGB4
			6'd2 : rdata = 41'b00011100000000001101111111000000011000000;
			// PEs: 5, 5 -> 
			// srcs: (120, 3)(3) 1, (226) -6 --> (280) -6:NM0, NI0, *, 
			6'd3 : rdata = 41'b00011100000000001010000000000000000000000;
			// PEs: 5, 5 -> 5
			// srcs: (123, 4)(63) 6, (280) -6 --> (334) 12:NW0, ALU, -, NW0
			6'd4 : rdata = 41'b00010010000000000011111111100100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 6) begin
	always @(*) begin
		case(address)
			// PEs: 6, 6 -> 
			// srcs: (1, 0)(9) 1, (64) 7 --> (118) 7:ND0, NW0, *, 
			6'd0 : rdata = 41'b00011011000000000100000000000000000000000;
			// PEs: 5, 6 -> 0
			// srcs: (4, 1)(117) 12, (118) 7 --> (170) 19:PENB, ALU, +, PEGB0
			6'd1 : rdata = 41'b00001110111111100011111111100000010000000;
			// PEs: 0, 6 -> 7
			// srcs: (118, 2)(221) -3, (9) 1 --> (227) -3:PEGB0, ND0, *, PENB
			6'd2 : rdata = 41'b00011111000000000110000000000000100000000;
			// PEs: 6, 7 -> 6
			// srcs: (127, 3)(64) 7, (281) -3 --> (335) 10:NW0, PEGB7, -, NW0
			6'd3 : rdata = 41'b00010010000000001110000111000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 7) begin
	always @(*) begin
		case(address)
			// PEs: 7, 7 -> 0
			// srcs: (1, 0)(11) 8, (66) 9 --> (120) 72:ND0, NW0, *, PENB
			6'd0 : rdata = 41'b00011011000000000100000000000000100000000;
			// PEs: 0, 7 -> 7
			// srcs: (120, 1)(221) -3, (11) 8 --> (229) -24:PEGB0, ND0, *, NI0
			6'd1 : rdata = 41'b00011111000000000110000000010000000000000;
			// PEs: 7, 6 -> 6
			// srcs: (121, 2)(3) 1, (227) -3 --> (281) -3:NM0, PENB, *, PEGB6
			6'd2 : rdata = 41'b00011100000000001101111111000000011100000;
			// PEs: 7, 7 -> 
			// srcs: (123, 3)(3) 1, (229) -24 --> (283) -24:NM0, NI0, *, 
			6'd3 : rdata = 41'b00011100000000001010000000000000000000000;
			// PEs: 7, 7 -> 7
			// srcs: (126, 4)(66) 9, (283) -24 --> (337) 33:NW0, ALU, -, NW0
			6'd4 : rdata = 41'b00010010000000000011111111100100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 8) begin
	always @(*) begin
		case(address)
			// PEs: 0 -> 9
			// srcs: (5, 0)(120) 72 --> (120) 72:PUNB, pass, PENB
			6'd0 : rdata = 41'b11000110111111110000000000000000100000000;
			// PEs: 15 -> 16
			// srcs: (6, 2)(180) 78 --> (180) 78:PENB, pass, PUNB
			6'd1 : rdata = 41'b11000110111111100000000000000001000000000;
			// PEs: 13 -> 32
			// srcs: (9, 1)(176) 86 --> (176) 86:PEGB5, pass, PUGB4
			6'd2 : rdata = 41'b11000111000010100000000000000000000001100;
			// PEs: 32 -> 8
			// srcs: (14, 3)(202) 76 --> (202) 76:PUGB4, pass, NI0
			6'd3 : rdata = 41'b11000111000010010000000000010000000000000;
			// PEs: 56 -> 9
			// srcs: (15, 4)(153) 0 --> (153) 0:PUGB7, pass, PENB
			6'd4 : rdata = 41'b11000111000011110000000000000000100000000;
			// PEs: 10 -> 24
			// srcs: (19, 6)(175) 147 --> (175) 147:PEGB2, pass, PUGB3
			6'd5 : rdata = 41'b11000111000001000000000000000000000001011;
			// PEs: 8 -> 9
			// srcs: (21, 5)(202) 76 --> (202) 76:NI0, pass, PENB
			6'd6 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 24 -> 8
			// srcs: (22, 7)(195) 105 --> (195) 105:PUGB3, pass, NI0
			6'd7 : rdata = 41'b11000111000001110000000000010000000000000;
			// PEs: 0 -> 9
			// srcs: (27, 8)(197) 55 --> (197) 55:PUNB, pass, PENB
			6'd8 : rdata = 41'b11000110111111110000000000000000100000000;
			// PEs: 9 -> 16
			// srcs: (28, 10)(203) 76 --> (203) 76:PEGB1, pass, PUNB
			6'd9 : rdata = 41'b11000111000000100000000000000001000000000;
			// PEs: 8 -> 9
			// srcs: (37, 9)(195) 105 --> (195) 105:NI0, pass, PENB
			6'd10 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 9 -> 16
			// srcs: (44, 11)(198) 160 --> (198) 160:PEGB1, pass, PUNB
			6'd11 : rdata = 41'b11000111000000100000000000000001000000000;
			// PEs: 32 -> 9
			// srcs: (116, 12)(221) -3 --> (221) -3:PUGB4, pass, PENB
			6'd12 : rdata = 41'b11000111000010010000000000000000100000000;
			// PEs: 32 -> 10
			// srcs: (117, 13)(221) -3 --> (221) -3:PUGB4, pass, PEGB2
			6'd13 : rdata = 41'b11000111000010010000000000000000010100000;
			// PEs: 32 -> 11
			// srcs: (118, 14)(221) -3 --> (221) -3:PUGB4, pass, PEGB3
			6'd14 : rdata = 41'b11000111000010010000000000000000010110000;
			// PEs: 32 -> 12
			// srcs: (119, 15)(221) -3 --> (221) -3:PUGB4, pass, PEGB4
			6'd15 : rdata = 41'b11000111000010010000000000000000011000000;
			// PEs: 32 -> 13
			// srcs: (120, 16)(221) -3 --> (221) -3:PUGB4, pass, PEGB5
			6'd16 : rdata = 41'b11000111000010010000000000000000011010000;
			// PEs: 32 -> 14
			// srcs: (122, 17)(221) -3 --> (221) -3:PUGB4, pass, PEGB6
			6'd17 : rdata = 41'b11000111000010010000000000000000011100000;
			// PEs: 32 -> 15
			// srcs: (123, 18)(221) -3 --> (221) -3:PUGB4, pass, PEGB7
			6'd18 : rdata = 41'b11000111000010010000000000000000011110000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 9) begin
	always @(*) begin
		case(address)
			// PEs: 9, 9 -> 
			// srcs: (1, 0)(12) 6, (67) 4 --> (121) 24:ND0, NW0, *, 
			6'd0 : rdata = 41'b00011011000000000100000000000000000000000;
			// PEs: 8, 9 -> 10
			// srcs: (8, 1)(120) 72, (121) 24 --> (173) 96:PENB, ALU, +, PENB
			6'd1 : rdata = 41'b00001110111111100011111111100000100000000;
			// PEs: 8 -> 
			// srcs: (17, 2)(153) 0 --> (153) 0:PENB, pass, 
			6'd2 : rdata = 41'b11000110111111100000000000000000000000000;
			// PEs: 8, 9 -> 8
			// srcs: (23, 3)(202) 76, (153) 0 --> (203) 76:PENB, ALU, +, PEGB0
			6'd3 : rdata = 41'b00001110111111100011111111100000010000000;
			// PEs: 8 -> 
			// srcs: (29, 4)(197) 55 --> (197) 55:PENB, pass, 
			6'd4 : rdata = 41'b11000110111111100000000000000000000000000;
			// PEs: 8, 9 -> 8
			// srcs: (39, 5)(195) 105, (197) 55 --> (198) 160:PENB, ALU, +, PEGB0
			6'd5 : rdata = 41'b00001110111111100011111111100000010000000;
			// PEs: 8, 9 -> 10
			// srcs: (118, 6)(221) -3, (12) 6 --> (230) -18:PENB, ND0, *, PENB
			6'd6 : rdata = 41'b00011110111111100110000000000000100000000;
			// PEs: 9, 10 -> 9
			// srcs: (127, 7)(67) 4, (284) -18 --> (338) 22:NW0, PEGB2, -, NW0
			6'd7 : rdata = 41'b00010010000000001110000010000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 10) begin
	always @(*) begin
		case(address)
			// PEs: 10, 10 -> 11
			// srcs: (1, 0)(13) 3, (68) 5 --> (122) 15:ND0, NW0, *, PENB
			6'd0 : rdata = 41'b00011011000000000100000000000000100000000;
			// PEs: 9, 11 -> 8
			// srcs: (14, 1)(173) 96, (174) 51 --> (175) 147:PENB, PEGB3, +, PEGB0
			6'd1 : rdata = 41'b00001110111111101110000011000000010000000;
			// PEs: 10, 9 -> 9
			// srcs: (121, 3)(3) 1, (230) -18 --> (284) -18:NM0, PENB, *, PEGB1
			6'd2 : rdata = 41'b00011100000000001101111111000000010010000;
			// PEs: 8, 10 -> 11
			// srcs: (122, 2)(221) -3, (13) 3 --> (231) -9:PEGB0, ND0, *, PENB
			6'd3 : rdata = 41'b00011111000000000110000000000000100000000;
			// PEs: 10, 11 -> 10
			// srcs: (131, 4)(68) 5, (285) -9 --> (339) 14:NW0, PEGB3, -, NW0
			6'd4 : rdata = 41'b00010010000000001110000011000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 11) begin
	always @(*) begin
		case(address)
			// PEs: 11, 11 -> 
			// srcs: (1, 0)(14) 9, (69) 4 --> (123) 36:ND0, NW0, *, 
			6'd0 : rdata = 41'b00011011000000000100000000000000000000000;
			// PEs: 10, 11 -> 10
			// srcs: (4, 1)(122) 15, (123) 36 --> (174) 51:PENB, ALU, +, PEGB2
			6'd1 : rdata = 41'b00001110111111100011111111100000010100000;
			// PEs: 8, 11 -> 12
			// srcs: (123, 2)(221) -3, (14) 9 --> (232) -27:PEGB0, ND0, *, PENB
			6'd2 : rdata = 41'b00011111000000000110000000000000100000000;
			// PEs: 11, 10 -> 10
			// srcs: (125, 3)(3) 1, (231) -9 --> (285) -9:NM0, PENB, *, PEGB2
			6'd3 : rdata = 41'b00011100000000001101111111000000010100000;
			// PEs: 11, 12 -> 11
			// srcs: (132, 4)(69) 4, (286) -27 --> (340) 31:NW0, PEGB4, -, NW0
			6'd4 : rdata = 41'b00010010000000001110000100000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 12) begin
	always @(*) begin
		case(address)
			// PEs: 12, 12 -> 13
			// srcs: (1, 0)(15) 9, (70) 6 --> (124) 54:ND0, NW0, *, PENB
			6'd0 : rdata = 41'b00011011000000000100000000000000100000000;
			// PEs: 8, 12 -> 12
			// srcs: (124, 1)(221) -3, (15) 9 --> (233) -27:PEGB0, ND0, *, NI0
			6'd1 : rdata = 41'b00011111000000000110000000010000000000000;
			// PEs: 12, 11 -> 11
			// srcs: (126, 2)(3) 1, (232) -27 --> (286) -27:NM0, PENB, *, PEGB3
			6'd2 : rdata = 41'b00011100000000001101111111000000010110000;
			// PEs: 12, 12 -> 
			// srcs: (127, 3)(3) 1, (233) -27 --> (287) -27:NM0, NI0, *, 
			6'd3 : rdata = 41'b00011100000000001010000000000000000000000;
			// PEs: 12, 12 -> 12
			// srcs: (130, 4)(70) 6, (287) -27 --> (341) 33:NW0, ALU, -, NW0
			6'd4 : rdata = 41'b00010010000000000011111111100100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 13) begin
	always @(*) begin
		case(address)
			// PEs: 13, 13 -> 
			// srcs: (1, 0)(16) 4, (71) 8 --> (125) 32:ND0, NW0, *, 
			6'd0 : rdata = 41'b00011011000000000100000000000000000000000;
			// PEs: 12, 13 -> 8
			// srcs: (4, 1)(124) 54, (125) 32 --> (176) 86:PENB, ALU, +, PEGB0
			6'd1 : rdata = 41'b00001110111111100011111111100000010000000;
			// PEs: 8, 13 -> 14
			// srcs: (125, 2)(221) -3, (16) 4 --> (234) -12:PEGB0, ND0, *, PENB
			6'd2 : rdata = 41'b00011111000000000110000000000000100000000;
			// PEs: 13, 14 -> 13
			// srcs: (134, 3)(71) 8, (288) -12 --> (342) 20:NW0, PEGB6, -, NW0
			6'd3 : rdata = 41'b00010010000000001110000110000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 14) begin
	always @(*) begin
		case(address)
			// PEs: 14, 14 -> 15
			// srcs: (1, 0)(18) 9, (73) 7 --> (127) 63:ND0, NW0, *, PENB
			6'd0 : rdata = 41'b00011011000000000100000000000000100000000;
			// PEs: 8, 14 -> 14
			// srcs: (127, 1)(221) -3, (18) 9 --> (236) -27:PEGB0, ND0, *, NI0
			6'd1 : rdata = 41'b00011111000000000110000000010000000000000;
			// PEs: 14, 13 -> 13
			// srcs: (128, 2)(3) 1, (234) -12 --> (288) -12:NM0, PENB, *, PEGB5
			6'd2 : rdata = 41'b00011100000000001101111111000000011010000;
			// PEs: 14, 14 -> 
			// srcs: (130, 3)(3) 1, (236) -27 --> (290) -27:NM0, NI0, *, 
			6'd3 : rdata = 41'b00011100000000001010000000000000000000000;
			// PEs: 14, 14 -> 14
			// srcs: (133, 4)(73) 7, (290) -27 --> (344) 34:NW0, ALU, -, NW0
			6'd4 : rdata = 41'b00010010000000000011111111100100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 15) begin
	always @(*) begin
		case(address)
			// PEs: 15, 15 -> 
			// srcs: (1, 0)(19) 3, (74) 5 --> (128) 15:ND0, NW0, *, 
			6'd0 : rdata = 41'b00011011000000000100000000000000000000000;
			// PEs: 14, 15 -> 8
			// srcs: (4, 1)(127) 63, (128) 15 --> (180) 78:PENB, ALU, +, PENB
			6'd1 : rdata = 41'b00001110111111100011111111100000100000000;
			// PEs: 8, 15 -> 
			// srcs: (128, 2)(221) -3, (19) 3 --> (237) -9:PEGB0, ND0, *, 
			6'd2 : rdata = 41'b00011111000000000110000000000000000000000;
			// PEs: 15, 15 -> 
			// srcs: (131, 3)(3) 1, (237) -9 --> (291) -9:NM0, ALU, *, 
			6'd3 : rdata = 41'b00011100000000000011111111100000000000000;
			// PEs: 15, 15 -> 15
			// srcs: (134, 4)(74) 5, (291) -9 --> (345) 14:NW0, ALU, -, NW0
			6'd4 : rdata = 41'b00010010000000000011111111100100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 16) begin
	always @(*) begin
		case(address)
			// PEs: 23 -> 24
			// srcs: (3, 0)(137) 14 --> (137) 14:PENB, pass, PUNB
			6'd0 : rdata = 41'b11000110111111100000000000000001000000000;
			// PEs: 20 -> 48
			// srcs: (9, 5)(183) 3 --> (183) 3:PEGB4, pass, PUGB6
			6'd1 : rdata = 41'b11000111000010000000000000000000000001110;
			// PEs: 22 -> 56
			// srcs: (10, 6)(186) 87 --> (186) 87:PEGB6, pass, PUGB7
			6'd2 : rdata = 41'b11000111000011000000000000000000000001111;
			// PEs: 48 -> 16
			// srcs: (11, 2)(119) 18 --> (119) 18:PUGB6, pass, NI0
			6'd3 : rdata = 41'b11000111000011010000000000010000000000000;
			// PEs: 0 -> 17
			// srcs: (14, 1)(170) 19 --> (170) 19:PUGB0, pass, PENB
			6'd4 : rdata = 41'b11000111000000010000000000000000100000000;
			// PEs: 16 -> 17
			// srcs: (21, 3)(119) 18 --> (119) 18:NI0, pass, PENB
			6'd5 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 8 -> 17
			// srcs: (22, 4)(180) 78 --> (180) 78:PUNB, pass, PENB
			6'd6 : rdata = 41'b11000110111111110000000000000000100000000;
			// PEs: 32 -> 16
			// srcs: (23, 9)(201) 50 --> (201) 50:PUGB4, pass, NI0
			6'd7 : rdata = 41'b11000111000010010000000000010000000000000;
			// PEs: 17 -> 48
			// srcs: (28, 7)(171) 37 --> (171) 37:PEGB1, pass, PUGB6
			6'd8 : rdata = 41'b11000111000000100000000000000000000001110;
			// PEs: 17 -> 32
			// srcs: (29, 8)(182) 79 --> (182) 79:PEGB1, pass, PUGB4
			6'd9 : rdata = 41'b11000111000000100000000000000000000001100;
			// PEs: 8 -> 17
			// srcs: (30, 10)(203) 76 --> (203) 76:PUNB, pass, PENB
			6'd10 : rdata = 41'b11000110111111110000000000000000100000000;
			// PEs: 16 -> 17
			// srcs: (40, 11)(201) 50 --> (201) 50:NI0, pass, PENB
			6'd11 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 8 -> 17
			// srcs: (46, 12)(198) 160 --> (198) 160:PUNB, pass, PENB
			6'd12 : rdata = 41'b11000110111111110000000000000000100000000;
			// PEs: 17 -> 24
			// srcs: (57, 13)(205) 286 --> (205) 286:PEGB1, pass, PUNB
			6'd13 : rdata = 41'b11000111000000100000000000000001000000000;
			// PEs: 32 -> 17
			// srcs: (124, 14)(221) -3 --> (221) -3:PUGB4, pass, PENB
			6'd14 : rdata = 41'b11000111000010010000000000000000100000000;
			// PEs: 32 -> 18
			// srcs: (125, 15)(221) -3 --> (221) -3:PUGB4, pass, PEGB2
			6'd15 : rdata = 41'b11000111000010010000000000000000010100000;
			// PEs: 32 -> 19
			// srcs: (126, 16)(221) -3 --> (221) -3:PUGB4, pass, PEGB3
			6'd16 : rdata = 41'b11000111000010010000000000000000010110000;
			// PEs: 32 -> 20
			// srcs: (127, 17)(221) -3 --> (221) -3:PUGB4, pass, PEGB4
			6'd17 : rdata = 41'b11000111000010010000000000000000011000000;
			// PEs: 32 -> 21
			// srcs: (129, 18)(221) -3 --> (221) -3:PUGB4, pass, PEGB5
			6'd18 : rdata = 41'b11000111000010010000000000000000011010000;
			// PEs: 32 -> 22
			// srcs: (130, 19)(221) -3 --> (221) -3:PUGB4, pass, PEGB6
			6'd19 : rdata = 41'b11000111000010010000000000000000011100000;
			// PEs: 32 -> 23
			// srcs: (132, 20)(221) -3 --> (221) -3:PUGB4, pass, PEGB7
			6'd20 : rdata = 41'b11000111000010010000000000000000011110000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 17) begin
	always @(*) begin
		case(address)
			// PEs: 17, 17 -> 18
			// srcs: (1, 0)(20) 1, (75) 0 --> (129) 0:ND0, NW0, *, PENB
			6'd0 : rdata = 41'b00011011000000000100000000000000100000000;
			// PEs: 16 -> 
			// srcs: (16, 1)(170) 19 --> (170) 19:PENB, pass, 
			6'd1 : rdata = 41'b11000110111111100000000000000000000000000;
			// PEs: 17, 16 -> 16
			// srcs: (23, 2)(170) 19, (119) 18 --> (171) 37:ALU, PENB, +, PEGB0
			6'd2 : rdata = 41'b00001001111111111101111111000000010000000;
			// PEs: 16, 18 -> 16
			// srcs: (24, 3)(180) 78, (181) 1 --> (182) 79:PENB, PEGB2, +, PEGB0
			6'd3 : rdata = 41'b00001110111111101110000010000000010000000;
			// PEs: 16 -> 
			// srcs: (32, 4)(203) 76 --> (203) 76:PENB, pass, 
			6'd4 : rdata = 41'b11000110111111100000000000000000000000000;
			// PEs: 16, 17 -> 
			// srcs: (42, 5)(201) 50, (203) 76 --> (204) 126:PENB, ALU, +, 
			6'd5 : rdata = 41'b00001110111111100011111111100000000000000;
			// PEs: 16, 17 -> 16
			// srcs: (52, 6)(198) 160, (204) 126 --> (205) 286:PENB, ALU, +, PEGB0
			6'd6 : rdata = 41'b00001110111111100011111111100000010000000;
			// PEs: 16, 17 -> 18
			// srcs: (126, 7)(221) -3, (20) 1 --> (238) -3:PENB, ND0, *, PENB
			6'd7 : rdata = 41'b00011110111111100110000000000000100000000;
			// PEs: 17, 18 -> 17
			// srcs: (135, 8)(75) 0, (292) -3 --> (346) 3:NW0, PEGB2, -, NW0
			6'd8 : rdata = 41'b00010010000000001110000010000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 18) begin
	always @(*) begin
		case(address)
			// PEs: 18, 18 -> 
			// srcs: (1, 0)(21) 1, (76) 1 --> (130) 1:ND0, NW0, *, 
			6'd0 : rdata = 41'b00011011000000000100000000000000000000000;
			// PEs: 17, 18 -> 17
			// srcs: (4, 1)(129) 0, (130) 1 --> (181) 1:PENB, ALU, +, PEGB1
			6'd1 : rdata = 41'b00001110111111100011111111100000010010000;
			// PEs: 18, 17 -> 17
			// srcs: (129, 3)(3) 1, (238) -3 --> (292) -3:NM0, PENB, *, PEGB1
			6'd2 : rdata = 41'b00011100000000001101111111000000010010000;
			// PEs: 16, 18 -> 19
			// srcs: (130, 2)(221) -3, (21) 1 --> (239) -3:PEGB0, ND0, *, PENB
			6'd3 : rdata = 41'b00011111000000000110000000000000100000000;
			// PEs: 18, 19 -> 18
			// srcs: (139, 4)(76) 1, (293) -3 --> (347) 4:NW0, PEGB3, -, NW0
			6'd4 : rdata = 41'b00010010000000001110000011000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 19) begin
	always @(*) begin
		case(address)
			// PEs: 19, 19 -> 20
			// srcs: (1, 0)(22) 1, (77) 3 --> (131) 3:ND0, NW0, *, PENB
			6'd0 : rdata = 41'b00011011000000000100000000000000100000000;
			// PEs: 16, 19 -> 19
			// srcs: (131, 1)(221) -3, (22) 1 --> (240) -3:PEGB0, ND0, *, NI0
			6'd1 : rdata = 41'b00011111000000000110000000010000000000000;
			// PEs: 19, 18 -> 18
			// srcs: (133, 2)(3) 1, (239) -3 --> (293) -3:NM0, PENB, *, PEGB2
			6'd2 : rdata = 41'b00011100000000001101111111000000010100000;
			// PEs: 19, 19 -> 
			// srcs: (134, 3)(3) 1, (240) -3 --> (294) -3:NM0, NI0, *, 
			6'd3 : rdata = 41'b00011100000000001010000000000000000000000;
			// PEs: 19, 19 -> 19
			// srcs: (137, 4)(77) 3, (294) -3 --> (348) 6:NW0, ALU, -, NW0
			6'd4 : rdata = 41'b00010010000000000011111111100100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 20) begin
	always @(*) begin
		case(address)
			// PEs: 20, 20 -> 
			// srcs: (1, 0)(23) 0, (78) 9 --> (132) 0:ND0, NW0, *, 
			6'd0 : rdata = 41'b00011011000000000100000000000000000000000;
			// PEs: 19, 20 -> 16
			// srcs: (4, 1)(131) 3, (132) 0 --> (183) 3:PENB, ALU, +, PEGB0
			6'd1 : rdata = 41'b00001110111111100011111111100000010000000;
			// PEs: 16, 20 -> 21
			// srcs: (132, 2)(221) -3, (23) 0 --> (241) 0:PEGB0, ND0, *, PENB
			6'd2 : rdata = 41'b00011111000000000110000000000000100000000;
			// PEs: 20, 21 -> 20
			// srcs: (141, 3)(78) 9, (295) 0 --> (349) 9:NW0, PEGB5, -, NW0
			6'd3 : rdata = 41'b00010010000000001110000101000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 21) begin
	always @(*) begin
		case(address)
			// PEs: 21, 21 -> 22
			// srcs: (1, 0)(25) 3, (80) 2 --> (134) 6:ND0, NW0, *, PENB
			6'd0 : rdata = 41'b00011011000000000100000000000000100000000;
			// PEs: 16, 21 -> 21
			// srcs: (134, 1)(221) -3, (25) 3 --> (243) -9:PEGB0, ND0, *, NI0
			6'd1 : rdata = 41'b00011111000000000110000000010000000000000;
			// PEs: 21, 20 -> 20
			// srcs: (135, 2)(3) 1, (241) 0 --> (295) 0:NM0, PENB, *, PEGB4
			6'd2 : rdata = 41'b00011100000000001101111111000000011000000;
			// PEs: 21, 21 -> 
			// srcs: (137, 3)(3) 1, (243) -9 --> (297) -9:NM0, NI0, *, 
			6'd3 : rdata = 41'b00011100000000001010000000000000000000000;
			// PEs: 21, 21 -> 21
			// srcs: (140, 4)(80) 2, (297) -9 --> (351) 11:NW0, ALU, -, NW0
			6'd4 : rdata = 41'b00010010000000000011111111100100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 22) begin
	always @(*) begin
		case(address)
			// PEs: 22, 22 -> 
			// srcs: (1, 0)(26) 9, (81) 9 --> (135) 81:ND0, NW0, *, 
			6'd0 : rdata = 41'b00011011000000000100000000000000000000000;
			// PEs: 21, 22 -> 16
			// srcs: (4, 1)(134) 6, (135) 81 --> (186) 87:PENB, ALU, +, PEGB0
			6'd1 : rdata = 41'b00001110111111100011111111100000010000000;
			// PEs: 16, 22 -> 23
			// srcs: (135, 2)(221) -3, (26) 9 --> (244) -27:PEGB0, ND0, *, PENB
			6'd2 : rdata = 41'b00011111000000000110000000000000100000000;
			// PEs: 22, 23 -> 22
			// srcs: (144, 3)(81) 9, (298) -27 --> (352) 36:NW0, PEGB7, -, NW0
			6'd3 : rdata = 41'b00010010000000001110000111000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 23) begin
	always @(*) begin
		case(address)
			// PEs: 23, 23 -> 16
			// srcs: (1, 0)(28) 2, (83) 7 --> (137) 14:ND0, NW0, *, PENB
			6'd0 : rdata = 41'b00011011000000000100000000000000100000000;
			// PEs: 16, 23 -> 23
			// srcs: (137, 1)(221) -3, (28) 2 --> (246) -6:PEGB0, ND0, *, NI0
			6'd1 : rdata = 41'b00011111000000000110000000010000000000000;
			// PEs: 23, 22 -> 22
			// srcs: (138, 2)(3) 1, (244) -27 --> (298) -27:NM0, PENB, *, PEGB6
			6'd2 : rdata = 41'b00011100000000001101111111000000011100000;
			// PEs: 23, 23 -> 
			// srcs: (140, 3)(3) 1, (246) -6 --> (300) -6:NM0, NI0, *, 
			6'd3 : rdata = 41'b00011100000000001010000000000000000000000;
			// PEs: 23, 23 -> 23
			// srcs: (143, 4)(83) 7, (300) -6 --> (354) 13:NW0, ALU, -, NW0
			6'd4 : rdata = 41'b00010010000000000011111111100100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 24) begin
	always @(*) begin
		case(address)
			// PEs: 16 -> 25
			// srcs: (5, 0)(137) 14 --> (137) 14:PUNB, pass, PENB
			6'd0 : rdata = 41'b11000110111111110000000000000000100000000;
			// PEs: 31 -> 0
			// srcs: (6, 2)(196) 7 --> (196) 7:PENB, pass, PUGB0
			6'd1 : rdata = 41'b11000110111111100000000000000000000001000;
			// PEs: 48 -> 25
			// srcs: (8, 1)(139) 49 --> (139) 49:PUGB6, pass, PENB
			6'd2 : rdata = 41'b11000111000011010000000000000000100000000;
			// PEs: 26 -> 8
			// srcs: (17, 7)(195) 105 --> (195) 105:PEGB2, pass, PUGB1
			6'd3 : rdata = 41'b11000111000001000000000000000000000001001;
			// PEs: 25 -> 40
			// srcs: (23, 6)(189) 78 --> (189) 78:PEGB1, pass, PUGB5
			6'd4 : rdata = 41'b11000111000000100000000000000000000001101;
			// PEs: 8 -> 24
			// srcs: (24, 3)(175) 147 --> (175) 147:PUGB1, pass, NI0
			6'd5 : rdata = 41'b11000111000000110000000000010000000000000;
			// PEs: 32 -> 25
			// srcs: (33, 4)(177) 158 --> (177) 158:PUGB4, pass, PENB
			6'd6 : rdata = 41'b11000111000010010000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (40, 5)(175) 147 --> (175) 147:NI0, pass, PENB
			6'd7 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 25 -> 48
			// srcs: (47, 8)(178) 305 --> (178) 305:PEGB1, pass, PUGB6
			6'd8 : rdata = 41'b11000111000000100000000000000000000001110;
			// PEs: 16 -> 24
			// srcs: (59, 9)(205) 286 --> (205) 286:PUNB, pass, NI0
			6'd9 : rdata = 41'b11000110111111110000000000010000000000000;
			// PEs: 0 -> 25
			// srcs: (63, 10)(217) 194 --> (217) 194:PUGB0, pass, PENB
			6'd10 : rdata = 41'b11000111000000010000000000000000100000000;
			// PEs: 24 -> 25
			// srcs: (70, 11)(205) 286 --> (205) 286:NI0, pass, PENB
			6'd11 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 25 -> 32
			// srcs: (77, 12)(218) 480 --> (218) 480:PEGB1, pass, PUNB
			6'd12 : rdata = 41'b11000111000000100000000000000001000000000;
			// PEs: 32 -> 25
			// srcs: (133, 13)(221) -3 --> (221) -3:PUGB4, pass, PENB
			6'd13 : rdata = 41'b11000111000010010000000000000000100000000;
			// PEs: 32 -> 26
			// srcs: (135, 14)(221) -3 --> (221) -3:PUGB4, pass, PEGB2
			6'd14 : rdata = 41'b11000111000010010000000000000000010100000;
			// PEs: 32 -> 27
			// srcs: (136, 15)(221) -3 --> (221) -3:PUGB4, pass, PEGB3
			6'd15 : rdata = 41'b11000111000010010000000000000000010110000;
			// PEs: 32 -> 28
			// srcs: (137, 16)(221) -3 --> (221) -3:PUGB4, pass, PEGB4
			6'd16 : rdata = 41'b11000111000010010000000000000000011000000;
			// PEs: 32 -> 29
			// srcs: (138, 17)(221) -3 --> (221) -3:PUGB4, pass, PEGB5
			6'd17 : rdata = 41'b11000111000010010000000000000000011010000;
			// PEs: 32 -> 30
			// srcs: (139, 18)(221) -3 --> (221) -3:PUGB4, pass, PEGB6
			6'd18 : rdata = 41'b11000111000010010000000000000000011100000;
			// PEs: 32 -> 31
			// srcs: (140, 19)(221) -3 --> (221) -3:PUGB4, pass, PEGB7
			6'd19 : rdata = 41'b11000111000010010000000000000000011110000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 25) begin
	always @(*) begin
		case(address)
			// PEs: 25, 25 -> 
			// srcs: (1, 0)(29) 5, (84) 3 --> (138) 15:ND0, NW0, *, 
			6'd0 : rdata = 41'b00011011000000000100000000000000000000000;
			// PEs: 24, 25 -> 
			// srcs: (8, 1)(137) 14, (138) 15 --> (188) 29:PENB, ALU, +, 
			6'd1 : rdata = 41'b00001110111111100011111111100000000000000;
			// PEs: 25, 24 -> 24
			// srcs: (18, 2)(188) 29, (139) 49 --> (189) 78:ALU, PENB, +, PEGB0
			6'd2 : rdata = 41'b00001001111111111101111111000000010000000;
			// PEs: 24 -> 
			// srcs: (35, 3)(177) 158 --> (177) 158:PENB, pass, 
			6'd3 : rdata = 41'b11000110111111100000000000000000000000000;
			// PEs: 24, 25 -> 24
			// srcs: (42, 4)(175) 147, (177) 158 --> (178) 305:PENB, ALU, +, PEGB0
			6'd4 : rdata = 41'b00001110111111100011111111100000010000000;
			// PEs: 24 -> 
			// srcs: (65, 5)(217) 194 --> (217) 194:PENB, pass, 
			6'd5 : rdata = 41'b11000110111111100000000000000000000000000;
			// PEs: 24, 25 -> 24
			// srcs: (72, 6)(205) 286, (217) 194 --> (218) 480:PENB, ALU, +, PEGB0
			6'd6 : rdata = 41'b00001110111111100011111111100000010000000;
			// PEs: 24, 25 -> 26
			// srcs: (135, 7)(221) -3, (29) 5 --> (247) -15:PENB, ND0, *, PENB
			6'd7 : rdata = 41'b00011110111111100110000000000000100000000;
			// PEs: 25, 26 -> 25
			// srcs: (144, 8)(84) 3, (301) -15 --> (355) 18:NW0, PEGB2, -, NW0
			6'd8 : rdata = 41'b00010010000000001110000010000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 26) begin
	always @(*) begin
		case(address)
			// PEs: 26, 26 -> 27
			// srcs: (1, 0)(31) 9, (86) 5 --> (140) 45:ND0, NW0, *, PENB
			6'd0 : rdata = 41'b00011011000000000100000000000000100000000;
			// PEs: 29 -> 
			// srcs: (9, 1)(194) 45 --> (194) 45:PEGB5, pass, 
			6'd1 : rdata = 41'b11000111000010100000000000000000000000000;
			// PEs: 27, 26 -> 24
			// srcs: (12, 2)(193) 60, (194) 45 --> (195) 105:PEGB3, ALU, +, PEGB0
			6'd2 : rdata = 41'b00001111000001100011111111100000010000000;
			// PEs: 26, 25 -> 25
			// srcs: (138, 4)(3) 1, (247) -15 --> (301) -15:NM0, PENB, *, PEGB1
			6'd3 : rdata = 41'b00011100000000001101111111000000010010000;
			// PEs: 24, 26 -> 27
			// srcs: (140, 3)(221) -3, (31) 9 --> (249) -27:PEGB0, ND0, *, PENB
			6'd4 : rdata = 41'b00011111000000000110000000000000100000000;
			// PEs: 26, 27 -> 26
			// srcs: (149, 5)(86) 5, (303) -27 --> (357) 32:NW0, PEGB3, -, NW0
			6'd5 : rdata = 41'b00010010000000001110000011000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 27) begin
	always @(*) begin
		case(address)
			// PEs: 27, 27 -> 
			// srcs: (1, 0)(32) 3, (87) 5 --> (141) 15:ND0, NW0, *, 
			6'd0 : rdata = 41'b00011011000000000100000000000000000000000;
			// PEs: 26, 27 -> 26
			// srcs: (4, 1)(140) 45, (141) 15 --> (193) 60:PENB, ALU, +, PEGB2
			6'd1 : rdata = 41'b00001110111111100011111111100000010100000;
			// PEs: 24, 27 -> 28
			// srcs: (141, 2)(221) -3, (32) 3 --> (250) -9:PEGB0, ND0, *, PENB
			6'd2 : rdata = 41'b00011111000000000110000000000000100000000;
			// PEs: 27, 26 -> 26
			// srcs: (143, 3)(3) 1, (249) -27 --> (303) -27:NM0, PENB, *, PEGB2
			6'd3 : rdata = 41'b00011100000000001101111111000000010100000;
			// PEs: 27, 28 -> 27
			// srcs: (150, 4)(87) 5, (304) -9 --> (358) 14:NW0, PEGB4, -, NW0
			6'd4 : rdata = 41'b00010010000000001110000100000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 28) begin
	always @(*) begin
		case(address)
			// PEs: 28, 28 -> 29
			// srcs: (1, 0)(33) 0, (88) 0 --> (142) 0:ND0, NW0, *, PENB
			6'd0 : rdata = 41'b00011011000000000100000000000000100000000;
			// PEs: 24, 28 -> 28
			// srcs: (142, 1)(221) -3, (33) 0 --> (251) 0:PEGB0, ND0, *, NI0
			6'd1 : rdata = 41'b00011111000000000110000000010000000000000;
			// PEs: 28, 27 -> 27
			// srcs: (144, 2)(3) 1, (250) -9 --> (304) -9:NM0, PENB, *, PEGB3
			6'd2 : rdata = 41'b00011100000000001101111111000000010110000;
			// PEs: 28, 28 -> 
			// srcs: (145, 3)(3) 1, (251) 0 --> (305) 0:NM0, NI0, *, 
			6'd3 : rdata = 41'b00011100000000001010000000000000000000000;
			// PEs: 28, 28 -> 28
			// srcs: (148, 4)(88) 0, (305) 0 --> (359) 0:NW0, ALU, -, NW0
			6'd4 : rdata = 41'b00010010000000000011111111100100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 29) begin
	always @(*) begin
		case(address)
			// PEs: 29, 29 -> 
			// srcs: (1, 0)(34) 5, (89) 9 --> (143) 45:ND0, NW0, *, 
			6'd0 : rdata = 41'b00011011000000000100000000000000000000000;
			// PEs: 28, 29 -> 26
			// srcs: (4, 1)(142) 0, (143) 45 --> (194) 45:PENB, ALU, +, PEGB2
			6'd1 : rdata = 41'b00001110111111100011111111100000010100000;
			// PEs: 24, 29 -> 30
			// srcs: (143, 2)(221) -3, (34) 5 --> (252) -15:PEGB0, ND0, *, PENB
			6'd2 : rdata = 41'b00011111000000000110000000000000100000000;
			// PEs: 29, 30 -> 29
			// srcs: (152, 3)(89) 9, (306) -15 --> (360) 24:NW0, PEGB6, -, NW0
			6'd3 : rdata = 41'b00010010000000001110000110000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 30) begin
	always @(*) begin
		case(address)
			// PEs: 30, 30 -> 31
			// srcs: (1, 0)(35) 1, (90) 7 --> (144) 7:ND0, NW0, *, PENB
			6'd0 : rdata = 41'b00011011000000000100000000000000100000000;
			// PEs: 24, 30 -> 30
			// srcs: (144, 1)(221) -3, (35) 1 --> (253) -3:PEGB0, ND0, *, NI0
			6'd1 : rdata = 41'b00011111000000000110000000010000000000000;
			// PEs: 30, 29 -> 29
			// srcs: (146, 2)(3) 1, (252) -15 --> (306) -15:NM0, PENB, *, PEGB5
			6'd2 : rdata = 41'b00011100000000001101111111000000011010000;
			// PEs: 30, 30 -> 
			// srcs: (147, 3)(3) 1, (253) -3 --> (307) -3:NM0, NI0, *, 
			6'd3 : rdata = 41'b00011100000000001010000000000000000000000;
			// PEs: 30, 30 -> 30
			// srcs: (150, 4)(90) 7, (307) -3 --> (361) 10:NW0, ALU, -, NW0
			6'd4 : rdata = 41'b00010010000000000011111111100100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 31) begin
	always @(*) begin
		case(address)
			// PEs: 31, 31 -> 
			// srcs: (1, 0)(36) 0, (91) 3 --> (145) 0:ND0, NW0, *, 
			6'd0 : rdata = 41'b00011011000000000100000000000000000000000;
			// PEs: 30, 31 -> 24
			// srcs: (4, 1)(144) 7, (145) 0 --> (196) 7:PENB, ALU, +, PENB
			6'd1 : rdata = 41'b00001110111111100011111111100000100000000;
			// PEs: 24, 31 -> 
			// srcs: (145, 2)(221) -3, (36) 0 --> (254) 0:PEGB0, ND0, *, 
			6'd2 : rdata = 41'b00011111000000000110000000000000000000000;
			// PEs: 31, 31 -> 
			// srcs: (148, 3)(3) 1, (254) 0 --> (308) 0:NM0, ALU, *, 
			6'd3 : rdata = 41'b00011100000000000011111111100000000000000;
			// PEs: 31, 31 -> 31
			// srcs: (151, 4)(91) 3, (308) 0 --> (362) 3:NW0, ALU, -, NW0
			6'd4 : rdata = 41'b00010010000000000011111111100100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 32) begin
	always @(*) begin
		case(address)
			// PEs: 39 -> 40
			// srcs: (3, 0)(154) 6 --> (154) 6:PENB, pass, PUNB
			6'd0 : rdata = 41'b11000110111111100000000000000001000000000;
			// PEs: 38 -> 8
			// srcs: (9, 4)(202) 76 --> (202) 76:PEGB6, pass, PUGB1
			6'd1 : rdata = 41'b11000111000011000000000000000000000001001;
			// PEs: 48 -> 32
			// srcs: (12, 2)(126) 72 --> (126) 72:PUGB6, pass, NI0
			6'd2 : rdata = 41'b11000111000011010000000000010000000000000;
			// PEs: 8 -> 33
			// srcs: (14, 1)(176) 86 --> (176) 86:PUGB1, pass, PENB
			6'd3 : rdata = 41'b11000111000000110000000000000000100000000;
			// PEs: 35 -> 16
			// srcs: (15, 9)(201) 50 --> (201) 50:PEGB3, pass, PUGB2
			6'd4 : rdata = 41'b11000111000001100000000000000000000001010;
			// PEs: 32 -> 33
			// srcs: (21, 3)(126) 72 --> (126) 72:NI0, pass, PENB
			6'd5 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 33 -> 24
			// srcs: (28, 5)(177) 158 --> (177) 158:PEGB1, pass, PUGB3
			6'd6 : rdata = 41'b11000111000000100000000000000000000001011;
			// PEs: 16 -> 32
			// srcs: (34, 6)(182) 79 --> (182) 79:PUGB2, pass, NI0
			6'd7 : rdata = 41'b11000111000001010000000000010000000000000;
			// PEs: 48 -> 33
			// srcs: (35, 7)(184) 21 --> (184) 21:PUGB6, pass, PENB
			6'd8 : rdata = 41'b11000111000011010000000000000000100000000;
			// PEs: 32 -> 33
			// srcs: (41, 8)(182) 79 --> (182) 79:NI0, pass, PENB
			6'd9 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 33 -> 40
			// srcs: (48, 10)(185) 100 --> (185) 100:PEGB1, pass, PUNB
			6'd10 : rdata = 41'b11000111000000100000000000000001000000000;
			// PEs: 48 -> 32
			// srcs: (75, 11)(192) 697 --> (192) 697:PUGB6, pass, NI0
			6'd11 : rdata = 41'b11000111000011010000000000010000000000000;
			// PEs: 24 -> 33
			// srcs: (79, 12)(218) 480 --> (218) 480:PUNB, pass, PENB
			6'd12 : rdata = 41'b11000110111111110000000000000000100000000;
			// PEs: 32 -> 33
			// srcs: (89, 13)(192) 697 --> (192) 697:NI0, pass, PENB
			6'd13 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 34 -> 0
			// srcs: (100, 14)(221) -3 --> (221) -3:PEGB2, pass, PUGB0
			6'd14 : rdata = 41'b11000111000001000000000000000000000001000;
			// PEs: 34 -> 0
			// srcs: (104, 15)(221) -3 --> (221) -3:PEGB2, pass, PUGB0
			6'd15 : rdata = 41'b11000111000001000000000000000000000001000;
			// PEs: 34 -> 0
			// srcs: (105, 16)(221) -3 --> (221) -3:PEGB2, pass, PUGB0
			6'd16 : rdata = 41'b11000111000001000000000000000000000001000;
			// PEs: 34 -> 0
			// srcs: (106, 17)(221) -3 --> (221) -3:PEGB2, pass, PUGB0
			6'd17 : rdata = 41'b11000111000001000000000000000000000001000;
			// PEs: 34 -> 0
			// srcs: (107, 18)(221) -3 --> (221) -3:PEGB2, pass, PUGB0
			6'd18 : rdata = 41'b11000111000001000000000000000000000001000;
			// PEs: 34 -> 0
			// srcs: (108, 19)(221) -3 --> (221) -3:PEGB2, pass, PUGB0
			6'd19 : rdata = 41'b11000111000001000000000000000000000001000;
			// PEs: 34 -> 48
			// srcs: (109, 20)(221) -3 --> (221) -3:PEGB2, pass, PUGB6
			6'd20 : rdata = 41'b11000111000001000000000000000000000001110;
			// PEs: 34 -> 0
			// srcs: (110, 21)(221) -3 --> (221) -3:PEGB2, pass, PUGB0
			6'd21 : rdata = 41'b11000111000001000000000000000000000001000;
			// PEs: 34 -> 8
			// srcs: (111, 22)(221) -3 --> (221) -3:PEGB2, pass, PUGB1
			6'd22 : rdata = 41'b11000111000001000000000000000000000001001;
			// PEs: 34 -> 8
			// srcs: (112, 23)(221) -3 --> (221) -3:PEGB2, pass, PUGB1
			6'd23 : rdata = 41'b11000111000001000000000000000000000001001;
			// PEs: 34 -> 8
			// srcs: (113, 24)(221) -3 --> (221) -3:PEGB2, pass, PUGB1
			6'd24 : rdata = 41'b11000111000001000000000000000000000001001;
			// PEs: 34 -> 8
			// srcs: (114, 25)(221) -3 --> (221) -3:PEGB2, pass, PUGB1
			6'd25 : rdata = 41'b11000111000001000000000000000000000001001;
			// PEs: 34 -> 8
			// srcs: (115, 26)(221) -3 --> (221) -3:PEGB2, pass, PUGB1
			6'd26 : rdata = 41'b11000111000001000000000000000000000001001;
			// PEs: 34 -> 48
			// srcs: (116, 27)(221) -3 --> (221) -3:PEGB2, pass, PUGB6
			6'd27 : rdata = 41'b11000111000001000000000000000000000001110;
			// PEs: 34 -> 8
			// srcs: (117, 28)(221) -3 --> (221) -3:PEGB2, pass, PUGB1
			6'd28 : rdata = 41'b11000111000001000000000000000000000001001;
			// PEs: 34 -> 8
			// srcs: (118, 29)(221) -3 --> (221) -3:PEGB2, pass, PUGB1
			6'd29 : rdata = 41'b11000111000001000000000000000000000001001;
			// PEs: 34 -> 16
			// srcs: (119, 30)(221) -3 --> (221) -3:PEGB2, pass, PUGB2
			6'd30 : rdata = 41'b11000111000001000000000000000000000001010;
			// PEs: 34 -> 16
			// srcs: (120, 31)(221) -3 --> (221) -3:PEGB2, pass, PUGB2
			6'd31 : rdata = 41'b11000111000001000000000000000000000001010;
			// PEs: 34 -> 16
			// srcs: (121, 32)(221) -3 --> (221) -3:PEGB2, pass, PUGB2
			6'd32 : rdata = 41'b11000111000001000000000000000000000001010;
			// PEs: 34 -> 16
			// srcs: (122, 33)(221) -3 --> (221) -3:PEGB2, pass, PUGB2
			6'd33 : rdata = 41'b11000111000001000000000000000000000001010;
			// PEs: 34 -> 48
			// srcs: (123, 34)(221) -3 --> (221) -3:PEGB2, pass, PUGB6
			6'd34 : rdata = 41'b11000111000001000000000000000000000001110;
			// PEs: 34 -> 16
			// srcs: (124, 35)(221) -3 --> (221) -3:PEGB2, pass, PUGB2
			6'd35 : rdata = 41'b11000111000001000000000000000000000001010;
			// PEs: 34 -> 16
			// srcs: (125, 36)(221) -3 --> (221) -3:PEGB2, pass, PUGB2
			6'd36 : rdata = 41'b11000111000001000000000000000000000001010;
			// PEs: 34 -> 48
			// srcs: (126, 37)(221) -3 --> (221) -3:PEGB2, pass, PUGB6
			6'd37 : rdata = 41'b11000111000001000000000000000000000001110;
			// PEs: 34 -> 16
			// srcs: (127, 38)(221) -3 --> (221) -3:PEGB2, pass, PUGB2
			6'd38 : rdata = 41'b11000111000001000000000000000000000001010;
			// PEs: 34 -> 24
			// srcs: (128, 39)(221) -3 --> (221) -3:PEGB2, pass, PUGB3
			6'd39 : rdata = 41'b11000111000001000000000000000000000001011;
			// PEs: 34 -> 48
			// srcs: (129, 40)(221) -3 --> (221) -3:PEGB2, pass, PUGB6
			6'd40 : rdata = 41'b11000111000001000000000000000000000001110;
			// PEs: 34 -> 24
			// srcs: (130, 41)(221) -3 --> (221) -3:PEGB2, pass, PUGB3
			6'd41 : rdata = 41'b11000111000001000000000000000000000001011;
			// PEs: 34 -> 24
			// srcs: (131, 42)(221) -3 --> (221) -3:PEGB2, pass, PUGB3
			6'd42 : rdata = 41'b11000111000001000000000000000000000001011;
			// PEs: 34 -> 24
			// srcs: (132, 43)(221) -3 --> (221) -3:PEGB2, pass, PUGB3
			6'd43 : rdata = 41'b11000111000001000000000000000000000001011;
			// PEs: 34 -> 24
			// srcs: (133, 44)(221) -3 --> (221) -3:PEGB2, pass, PUGB3
			6'd44 : rdata = 41'b11000111000001000000000000000000000001011;
			// PEs: 34 -> 24
			// srcs: (134, 45)(221) -3 --> (221) -3:PEGB2, pass, PUGB3
			6'd45 : rdata = 41'b11000111000001000000000000000000000001011;
			// PEs: 34 -> 24
			// srcs: (135, 46)(221) -3 --> (221) -3:PEGB2, pass, PUGB3
			6'd46 : rdata = 41'b11000111000001000000000000000000000001011;
			// PEs: 34 -> 56
			// srcs: (136, 47)(221) -3 --> (221) -3:PEGB2, pass, PUGB7
			6'd47 : rdata = 41'b11000111000001000000000000000000000001111;
			// PEs: 34 -> 56
			// srcs: (142, 48)(221) -3 --> (221) -3:PEGB2, pass, PUGB7
			6'd48 : rdata = 41'b11000111000001000000000000000000000001111;
			// PEs: 34 -> 40
			// srcs: (144, 49)(221) -3 --> (221) -3:PEGB2, pass, PUNB
			6'd49 : rdata = 41'b11000111000001000000000000000001000000000;
			// PEs: 34 -> 40
			// srcs: (145, 50)(221) -3 --> (221) -3:PEGB2, pass, PUNB
			6'd50 : rdata = 41'b11000111000001000000000000000001000000000;
			// PEs: 34 -> 40
			// srcs: (146, 51)(221) -3 --> (221) -3:PEGB2, pass, PUNB
			6'd51 : rdata = 41'b11000111000001000000000000000001000000000;
			// PEs: 34 -> 40
			// srcs: (147, 52)(221) -3 --> (221) -3:PEGB2, pass, PUNB
			6'd52 : rdata = 41'b11000111000001000000000000000001000000000;
			// PEs: 34 -> 40
			// srcs: (148, 53)(221) -3 --> (221) -3:PEGB2, pass, PUNB
			6'd53 : rdata = 41'b11000111000001000000000000000001000000000;
			// PEs: 34 -> 56
			// srcs: (149, 54)(221) -3 --> (221) -3:PEGB2, pass, PUGB7
			6'd54 : rdata = 41'b11000111000001000000000000000000000001111;
			// PEs: 34 -> 40
			// srcs: (150, 55)(221) -3 --> (221) -3:PEGB2, pass, PUNB
			6'd55 : rdata = 41'b11000111000001000000000000000001000000000;
			// PEs: 34 -> 40
			// srcs: (151, 56)(221) -3 --> (221) -3:PEGB2, pass, PUNB
			6'd56 : rdata = 41'b11000111000001000000000000000001000000000;
			// PEs: 34 -> 56
			// srcs: (152, 57)(221) -3 --> (221) -3:PEGB2, pass, PUGB7
			6'd57 : rdata = 41'b11000111000001000000000000000000000001111;
			// PEs: 34 -> 48
			// srcs: (153, 58)(221) -3 --> (221) -3:PEGB2, pass, PUGB6
			6'd58 : rdata = 41'b11000111000001000000000000000000000001110;
			// PEs: 34 -> 48
			// srcs: (154, 59)(221) -3 --> (221) -3:PEGB2, pass, PUGB6
			6'd59 : rdata = 41'b11000111000001000000000000000000000001110;
			// PEs: 34 -> 56
			// srcs: (155, 60)(221) -3 --> (221) -3:PEGB2, pass, PUGB7
			6'd60 : rdata = 41'b11000111000001000000000000000000000001111;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 33) begin
	always @(*) begin
		case(address)
			// PEs: 33, 33 -> 34
			// srcs: (1, 0)(38) 1, (93) 3 --> (147) 3:ND0, NW0, *, PENB
			6'd0 : rdata = 41'b00011011000000000100000000000000100000000;
			// PEs: 32 -> 
			// srcs: (16, 1)(176) 86 --> (176) 86:PENB, pass, 
			6'd1 : rdata = 41'b11000110111111100000000000000000000000000;
			// PEs: 33, 32 -> 32
			// srcs: (23, 2)(176) 86, (126) 72 --> (177) 158:ALU, PENB, +, PEGB0
			6'd2 : rdata = 41'b00001001111111111101111111000000010000000;
			// PEs: 32 -> 
			// srcs: (37, 3)(184) 21 --> (184) 21:PENB, pass, 
			6'd3 : rdata = 41'b11000110111111100000000000000000000000000;
			// PEs: 32, 33 -> 32
			// srcs: (43, 4)(182) 79, (184) 21 --> (185) 100:PENB, ALU, +, PEGB0
			6'd4 : rdata = 41'b00001110111111100011111111100000010000000;
			// PEs: 32 -> 
			// srcs: (81, 5)(218) 480 --> (218) 480:PENB, pass, 
			6'd5 : rdata = 41'b11000110111111100000000000000000000000000;
			// PEs: 32, 33 -> 
			// srcs: (91, 6)(192) 697, (218) 480 --> (219) 1177:PENB, ALU, +, ALU
			6'd6 : rdata = 41'b00001110111111100011111111100000000000000;
			// PEs: 33 -> 34
			// srcs: (92, 7)(219) 1177 --> (220) 0:ALU, sigmoid, PENB
			6'd7 : rdata = 41'b10000001111111110000000000000000100000000;
			// PEs: 34, 33 -> 
			// srcs: (137, 8)(221) -3, (38) 1 --> (256) -3:PEGB2, ND0, *, 
			6'd8 : rdata = 41'b00011111000001000110000000000000000000000;
			// PEs: 33, 33 -> 
			// srcs: (140, 9)(3) 1, (256) -3 --> (310) -3:NM0, ALU, *, 
			6'd9 : rdata = 41'b00011100000000000011111111100000000000000;
			// PEs: 33, 33 -> 33
			// srcs: (143, 10)(93) 3, (310) -3 --> (364) 6:NW0, ALU, -, NW0
			6'd10 : rdata = 41'b00010010000000000011111111100100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 34) begin
	always @(*) begin
		case(address)
			// PEs: 34, 34 -> 
			// srcs: (1, 0)(39) 5, (94) 0 --> (148) 0:ND0, NW0, *, 
			6'd0 : rdata = 41'b00011011000000000100000000000000000000000;
			// PEs: 33, 34 -> 35
			// srcs: (4, 1)(147) 3, (148) 0 --> (199) 3:PENB, ALU, +, PENB
			6'd1 : rdata = 41'b00001110111111100011111111100000100000000;
			// PEs: 33, 34 -> 35, 32, 34
			// srcs: (95, 2)(220) 0, (58) 3 --> (221) -3:PENB, ND1, -, NI0, PENB, PEGB0
			6'd2 : rdata = 41'b00010110111111100110000000110000110000000;
			// PEs: 34 -> 32
			// srcs: (97, 3)(221) 0 --> (221) -3:ALU, pass, PEGB0
			6'd3 : rdata = 41'b11000001111111110000000000000000010000000;
			// PEs: 34 -> 32
			// srcs: (98, 4)(221) -3 --> (221) -3:NI0, pass, PEGB0
			6'd4 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 34 -> 32
			// srcs: (99, 5)(221) -3 --> (221) -3:NI0, pass, PEGB0
			6'd5 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 34 -> 32
			// srcs: (100, 6)(221) -3 --> (221) -3:NI0, pass, PEGB0
			6'd6 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 34 -> 32
			// srcs: (101, 7)(221) -3 --> (221) -3:NI0, pass, PEGB0
			6'd7 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 34 -> 32
			// srcs: (102, 8)(221) -3 --> (221) -3:NI0, pass, PEGB0
			6'd8 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 34 -> 32
			// srcs: (103, 9)(221) -3 --> (221) -3:NI0, pass, PEGB0
			6'd9 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 34 -> 32
			// srcs: (104, 10)(221) -3 --> (221) -3:NI0, pass, PEGB0
			6'd10 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 34 -> 32
			// srcs: (105, 11)(221) -3 --> (221) -3:NI0, pass, PEGB0
			6'd11 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 34 -> 32
			// srcs: (106, 12)(221) -3 --> (221) -3:NI0, pass, PEGB0
			6'd12 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 34 -> 32
			// srcs: (107, 13)(221) -3 --> (221) -3:NI0, pass, PEGB0
			6'd13 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 34 -> 32
			// srcs: (108, 14)(221) -3 --> (221) -3:NI0, pass, PEGB0
			6'd14 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 34 -> 32
			// srcs: (109, 15)(221) -3 --> (221) -3:NI0, pass, PEGB0
			6'd15 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 34 -> 32
			// srcs: (110, 16)(221) -3 --> (221) -3:NI0, pass, PEGB0
			6'd16 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 34 -> 32
			// srcs: (111, 17)(221) -3 --> (221) -3:NI0, pass, PEGB0
			6'd17 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 34 -> 32
			// srcs: (112, 18)(221) -3 --> (221) -3:NI0, pass, PEGB0
			6'd18 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 34 -> 32
			// srcs: (113, 19)(221) -3 --> (221) -3:NI0, pass, PEGB0
			6'd19 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 34 -> 32
			// srcs: (114, 20)(221) -3 --> (221) -3:NI0, pass, PEGB0
			6'd20 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 34 -> 32
			// srcs: (115, 21)(221) -3 --> (221) -3:NI0, pass, PEGB0
			6'd21 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 34 -> 32
			// srcs: (116, 22)(221) -3 --> (221) -3:NI0, pass, PEGB0
			6'd22 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 34 -> 32
			// srcs: (117, 23)(221) -3 --> (221) -3:NI0, pass, PEGB0
			6'd23 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 34 -> 32
			// srcs: (118, 24)(221) -3 --> (221) -3:NI0, pass, PEGB0
			6'd24 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 34 -> 32
			// srcs: (119, 25)(221) -3 --> (221) -3:NI0, pass, PEGB0
			6'd25 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 34 -> 32
			// srcs: (120, 26)(221) -3 --> (221) -3:NI0, pass, PEGB0
			6'd26 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 34 -> 32
			// srcs: (121, 27)(221) -3 --> (221) -3:NI0, pass, PEGB0
			6'd27 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 34 -> 32
			// srcs: (122, 28)(221) -3 --> (221) -3:NI0, pass, PEGB0
			6'd28 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 34 -> 32
			// srcs: (123, 29)(221) -3 --> (221) -3:NI0, pass, PEGB0
			6'd29 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 34 -> 32
			// srcs: (124, 30)(221) -3 --> (221) -3:NI0, pass, PEGB0
			6'd30 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 34 -> 32
			// srcs: (125, 31)(221) -3 --> (221) -3:NI0, pass, PEGB0
			6'd31 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 34 -> 32
			// srcs: (126, 32)(221) -3 --> (221) -3:NI0, pass, PEGB0
			6'd32 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 34 -> 32
			// srcs: (127, 33)(221) -3 --> (221) -3:NI0, pass, PEGB0
			6'd33 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 34 -> 32
			// srcs: (128, 34)(221) -3 --> (221) -3:NI0, pass, PEGB0
			6'd34 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 34 -> 32
			// srcs: (129, 35)(221) -3 --> (221) -3:NI0, pass, PEGB0
			6'd35 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 34 -> 33
			// srcs: (130, 36)(221) -3 --> (221) -3:NI0, pass, PEGB1
			6'd36 : rdata = 41'b11000101000000000000000000000000010010000;
			// PEs: 34, 34 -> 35
			// srcs: (131, 37)(221) -3, (39) 5 --> (257) -15:NI0, ND0, *, PENB
			6'd37 : rdata = 41'b00011101000000000110000000000000100000000;
			// PEs: 34 -> 36
			// srcs: (132, 38)(221) -3 --> (221) -3:NI0, pass, PEGB4
			6'd38 : rdata = 41'b11000101000000000000000000000000011000000;
			// PEs: 34 -> 37
			// srcs: (133, 39)(221) -3 --> (221) -3:NI0, pass, PEGB5
			6'd39 : rdata = 41'b11000101000000000000000000000000011010000;
			// PEs: 34 -> 38
			// srcs: (134, 40)(221) -3 --> (221) -3:NI0, pass, PEGB6
			6'd40 : rdata = 41'b11000101000000000000000000000000011100000;
			// PEs: 34 -> 32
			// srcs: (135, 41)(221) -3 --> (221) -3:NI0, pass, PEGB0
			6'd41 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 34 -> 39
			// srcs: (136, 42)(221) -3 --> (221) -3:NI0, pass, PEGB7
			6'd42 : rdata = 41'b11000101000000000000000000000000011110000;
			// PEs: 34 -> 32
			// srcs: (137, 43)(221) -3 --> (221) -3:NI0, pass, PEGB0
			6'd43 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 34 -> 32
			// srcs: (138, 44)(221) -3 --> (221) -3:NI0, pass, PEGB0
			6'd44 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 34 -> 32
			// srcs: (139, 45)(221) -3 --> (221) -3:NI0, pass, PEGB0
			6'd45 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 34 -> 32
			// srcs: (140, 46)(221) -3 --> (221) -3:NI0, pass, PEGB0
			6'd46 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 34 -> 32
			// srcs: (141, 47)(221) -3 --> (221) -3:NI0, pass, PEGB0
			6'd47 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 34 -> 32
			// srcs: (142, 48)(221) -3 --> (221) -3:NI0, pass, PEGB0
			6'd48 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 34 -> 32
			// srcs: (143, 49)(221) -3 --> (221) -3:NI0, pass, PEGB0
			6'd49 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 34 -> 32
			// srcs: (144, 50)(221) -3 --> (221) -3:NI0, pass, PEGB0
			6'd50 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 34 -> 32
			// srcs: (145, 51)(221) -3 --> (221) -3:NI0, pass, PEGB0
			6'd51 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 34 -> 32
			// srcs: (146, 52)(221) -3 --> (221) -3:NI0, pass, PEGB0
			6'd52 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 34 -> 32
			// srcs: (147, 53)(221) -3 --> (221) -3:NI0, pass, PEGB0
			6'd53 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 34 -> 32
			// srcs: (148, 54)(221) -3 --> (221) -3:NI0, pass, PEGB0
			6'd54 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 34, 35 -> 34
			// srcs: (149, 55)(94) 0, (311) -15 --> (365) 15:NW0, PEGB3, -, NW0
			6'd55 : rdata = 41'b00010010000000001110000011000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 35) begin
	always @(*) begin
		case(address)
			// PEs: 35, 35 -> 36
			// srcs: (1, 0)(40) 3, (95) 4 --> (149) 12:ND0, NW0, *, PENB
			6'd0 : rdata = 41'b00011011000000000100000000000000100000000;
			// PEs: 34, 36 -> 32
			// srcs: (10, 1)(199) 3, (200) 47 --> (201) 50:PENB, PEGB4, +, PEGB0
			6'd1 : rdata = 41'b00001110111111101110000100000000010000000;
			// PEs: 34, 35 -> 36
			// srcs: (98, 2)(221) -3, (40) 3 --> (258) -9:PENB, ND0, *, PENB
			6'd2 : rdata = 41'b00011110111111100110000000000000100000000;
			// PEs: 35, 36 -> 35
			// srcs: (107, 4)(95) 4, (312) -9 --> (366) 13:NW0, PEGB4, -, NW0
			6'd3 : rdata = 41'b00010010000000001110000100000100000000000;
			// PEs: 35, 34 -> 34
			// srcs: (134, 3)(3) 1, (257) -15 --> (311) -15:NM0, PENB, *, PEGB2
			6'd4 : rdata = 41'b00011100000000001101111111000000010100000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 36) begin
	always @(*) begin
		case(address)
			// PEs: 36, 36 -> 
			// srcs: (1, 0)(41) 5, (96) 7 --> (150) 35:ND0, NW0, *, 
			6'd0 : rdata = 41'b00011011000000000100000000000000000000000;
			// PEs: 35, 36 -> 35
			// srcs: (4, 1)(149) 12, (150) 35 --> (200) 47:PENB, ALU, +, PEGB3
			6'd1 : rdata = 41'b00001110111111100011111111100000010110000;
			// PEs: 36, 35 -> 35
			// srcs: (101, 3)(3) 1, (258) -9 --> (312) -9:NM0, PENB, *, PEGB3
			6'd2 : rdata = 41'b00011100000000001101111111000000010110000;
			// PEs: 34, 36 -> 37
			// srcs: (139, 2)(221) -3, (41) 5 --> (259) -15:PEGB2, ND0, *, PENB
			6'd3 : rdata = 41'b00011111000001000110000000000000100000000;
			// PEs: 36, 37 -> 36
			// srcs: (148, 4)(96) 7, (313) -15 --> (367) 22:NW0, PEGB5, -, NW0
			6'd4 : rdata = 41'b00010010000000001110000101000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 37) begin
	always @(*) begin
		case(address)
			// PEs: 37, 37 -> 38
			// srcs: (1, 0)(42) 3, (97) 4 --> (151) 12:ND0, NW0, *, PENB
			6'd0 : rdata = 41'b00011011000000000100000000000000100000000;
			// PEs: 34, 37 -> 37
			// srcs: (140, 1)(221) -3, (42) 3 --> (260) -9:PEGB2, ND0, *, NI0
			6'd1 : rdata = 41'b00011111000001000110000000010000000000000;
			// PEs: 37, 36 -> 36
			// srcs: (142, 2)(3) 1, (259) -15 --> (313) -15:NM0, PENB, *, PEGB4
			6'd2 : rdata = 41'b00011100000000001101111111000000011000000;
			// PEs: 37, 37 -> 
			// srcs: (143, 3)(3) 1, (260) -9 --> (314) -9:NM0, NI0, *, 
			6'd3 : rdata = 41'b00011100000000001010000000000000000000000;
			// PEs: 37, 37 -> 37
			// srcs: (146, 4)(97) 4, (314) -9 --> (368) 13:NW0, ALU, -, NW0
			6'd4 : rdata = 41'b00010010000000000011111111100100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 38) begin
	always @(*) begin
		case(address)
			// PEs: 38, 38 -> 
			// srcs: (1, 0)(43) 8, (98) 8 --> (152) 64:ND0, NW0, *, 
			6'd0 : rdata = 41'b00011011000000000100000000000000000000000;
			// PEs: 37, 38 -> 32
			// srcs: (4, 1)(151) 12, (152) 64 --> (202) 76:PENB, ALU, +, PEGB0
			6'd1 : rdata = 41'b00001110111111100011111111100000010000000;
			// PEs: 34, 38 -> 39
			// srcs: (141, 2)(221) -3, (43) 8 --> (261) -24:PEGB2, ND0, *, PENB
			6'd2 : rdata = 41'b00011111000001000110000000000000100000000;
			// PEs: 38, 39 -> 38
			// srcs: (150, 3)(98) 8, (315) -24 --> (369) 32:NW0, PEGB7, -, NW0
			6'd3 : rdata = 41'b00010010000000001110000111000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 39) begin
	always @(*) begin
		case(address)
			// PEs: 39, 39 -> 32
			// srcs: (1, 0)(45) 1, (100) 6 --> (154) 6:ND0, NW0, *, PENB
			6'd0 : rdata = 41'b00011011000000000100000000000000100000000;
			// PEs: 34, 39 -> 39
			// srcs: (143, 1)(221) -3, (45) 1 --> (263) -3:PEGB2, ND0, *, NI0
			6'd1 : rdata = 41'b00011111000001000110000000010000000000000;
			// PEs: 39, 38 -> 38
			// srcs: (144, 2)(3) 1, (261) -24 --> (315) -24:NM0, PENB, *, PEGB6
			6'd2 : rdata = 41'b00011100000000001101111111000000011100000;
			// PEs: 39, 39 -> 
			// srcs: (146, 3)(3) 1, (263) -3 --> (317) -3:NM0, NI0, *, 
			6'd3 : rdata = 41'b00011100000000001010000000000000000000000;
			// PEs: 39, 39 -> 39
			// srcs: (149, 4)(100) 6, (317) -3 --> (371) 9:NW0, ALU, -, NW0
			6'd4 : rdata = 41'b00010010000000000011111111100100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 40) begin
	always @(*) begin
		case(address)
			// PEs: 32 -> 41
			// srcs: (5, 0)(154) 6 --> (154) 6:PUNB, pass, PENB
			6'd0 : rdata = 41'b11000110111111110000000000000000100000000;
			// PEs: 47 -> 56
			// srcs: (6, 2)(212) 49 --> (212) 49:PENB, pass, PUGB7
			6'd1 : rdata = 41'b11000110111111100000000000000000000001111;
			// PEs: 56 -> 41
			// srcs: (13, 1)(160) 0 --> (160) 0:PUGB7, pass, PENB
			6'd2 : rdata = 41'b11000111000011110000000000000000100000000;
			// PEs: 42 -> 0
			// srcs: (25, 7)(211) 82 --> (211) 82:PEGB2, pass, PUGB0
			6'd3 : rdata = 41'b11000111000001000000000000000000000001000;
			// PEs: 56 -> 40
			// srcs: (33, 3)(187) 103 --> (187) 103:PUGB7, pass, NI0
			6'd4 : rdata = 41'b11000111000011110000000000010000000000000;
			// PEs: 24 -> 41
			// srcs: (34, 4)(189) 78 --> (189) 78:PUGB3, pass, PENB
			6'd5 : rdata = 41'b11000111000001110000000000000000100000000;
			// PEs: 40 -> 41
			// srcs: (40, 5)(187) 103 --> (187) 103:NI0, pass, PENB
			6'd6 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 32 -> 41
			// srcs: (50, 6)(185) 100 --> (185) 100:PUNB, pass, PENB
			6'd7 : rdata = 41'b11000110111111110000000000000000100000000;
			// PEs: 41 -> 48
			// srcs: (58, 8)(191) 281 --> (191) 281:PEGB1, pass, PUNB
			6'd8 : rdata = 41'b11000111000000100000000000000001000000000;
			// PEs: 32 -> 41
			// srcs: (146, 9)(221) -3 --> (221) -3:PUNB, pass, PENB
			6'd9 : rdata = 41'b11000110111111110000000000000000100000000;
			// PEs: 32 -> 42
			// srcs: (147, 10)(221) -3 --> (221) -3:PUNB, pass, PEGB2
			6'd10 : rdata = 41'b11000110111111110000000000000000010100000;
			// PEs: 32 -> 43
			// srcs: (148, 11)(221) -3 --> (221) -3:PUNB, pass, PEGB3
			6'd11 : rdata = 41'b11000110111111110000000000000000010110000;
			// PEs: 32 -> 44
			// srcs: (149, 12)(221) -3 --> (221) -3:PUNB, pass, PEGB4
			6'd12 : rdata = 41'b11000110111111110000000000000000011000000;
			// PEs: 32 -> 45
			// srcs: (150, 13)(221) -3 --> (221) -3:PUNB, pass, PEGB5
			6'd13 : rdata = 41'b11000110111111110000000000000000011010000;
			// PEs: 32 -> 46
			// srcs: (152, 14)(221) -3 --> (221) -3:PUNB, pass, PEGB6
			6'd14 : rdata = 41'b11000110111111110000000000000000011100000;
			// PEs: 32 -> 47
			// srcs: (153, 15)(221) -3 --> (221) -3:PUNB, pass, PEGB7
			6'd15 : rdata = 41'b11000110111111110000000000000000011110000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 41) begin
	always @(*) begin
		case(address)
			// PEs: 41, 41 -> 
			// srcs: (1, 0)(46) 5, (101) 9 --> (155) 45:ND0, NW0, *, 
			6'd0 : rdata = 41'b00011011000000000100000000000000000000000;
			// PEs: 40, 41 -> 42
			// srcs: (8, 1)(154) 6, (155) 45 --> (206) 51:PENB, ALU, +, PENB
			6'd1 : rdata = 41'b00001110111111100011111111100000100000000;
			// PEs: 45, 40 -> 42
			// srcs: (17, 2)(209) 31, (160) 0 --> (210) 31:PEGB5, PENB, +, PENB
			6'd2 : rdata = 41'b00001111000010101101111111000000100000000;
			// PEs: 40 -> 
			// srcs: (36, 3)(189) 78 --> (189) 78:PENB, pass, 
			6'd3 : rdata = 41'b11000110111111100000000000000000000000000;
			// PEs: 40, 41 -> 
			// srcs: (42, 4)(187) 103, (189) 78 --> (190) 181:PENB, ALU, +, 
			6'd4 : rdata = 41'b00001110111111100011111111100000000000000;
			// PEs: 40, 41 -> 40
			// srcs: (53, 5)(185) 100, (190) 181 --> (191) 281:PENB, ALU, +, PEGB0
			6'd5 : rdata = 41'b00001110111111100011111111100000010000000;
			// PEs: 40, 41 -> 42
			// srcs: (148, 6)(221) -3, (46) 5 --> (264) -15:PENB, ND0, *, PENB
			6'd6 : rdata = 41'b00011110111111100110000000000000100000000;
			// PEs: 41, 42 -> 41
			// srcs: (157, 7)(101) 9, (318) -15 --> (372) 24:NW0, PEGB2, -, NW0
			6'd7 : rdata = 41'b00010010000000001110000010000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 42) begin
	always @(*) begin
		case(address)
			// PEs: 42, 42 -> 43
			// srcs: (1, 0)(47) 0, (102) 2 --> (156) 0:ND0, NW0, *, PENB
			6'd0 : rdata = 41'b00011011000000000100000000000000100000000;
			// PEs: 41, 43 -> 
			// srcs: (14, 1)(206) 51, (207) 0 --> (208) 51:PENB, PEGB3, +, 
			6'd1 : rdata = 41'b00001110111111101110000011000000000000000;
			// PEs: 42, 41 -> 40
			// srcs: (20, 2)(208) 51, (210) 31 --> (211) 82:ALU, PENB, +, PEGB0
			6'd2 : rdata = 41'b00001001111111111101111111000000010000000;
			// PEs: 42, 41 -> 41
			// srcs: (151, 4)(3) 1, (264) -15 --> (318) -15:NM0, PENB, *, PEGB1
			6'd3 : rdata = 41'b00011100000000001101111111000000010010000;
			// PEs: 40, 42 -> 43
			// srcs: (152, 3)(221) -3, (47) 0 --> (265) 0:PEGB0, ND0, *, PENB
			6'd4 : rdata = 41'b00011111000000000110000000000000100000000;
			// PEs: 42, 43 -> 42
			// srcs: (161, 5)(102) 2, (319) 0 --> (373) 2:NW0, PEGB3, -, NW0
			6'd5 : rdata = 41'b00010010000000001110000011000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 43) begin
	always @(*) begin
		case(address)
			// PEs: 43, 43 -> 
			// srcs: (1, 0)(48) 0, (103) 6 --> (157) 0:ND0, NW0, *, 
			6'd0 : rdata = 41'b00011011000000000100000000000000000000000;
			// PEs: 42, 43 -> 42
			// srcs: (4, 1)(156) 0, (157) 0 --> (207) 0:PENB, ALU, +, PEGB2
			6'd1 : rdata = 41'b00001110111111100011111111100000010100000;
			// PEs: 40, 43 -> 44
			// srcs: (153, 2)(221) -3, (48) 0 --> (266) 0:PEGB0, ND0, *, PENB
			6'd2 : rdata = 41'b00011111000000000110000000000000100000000;
			// PEs: 43, 42 -> 42
			// srcs: (155, 3)(3) 1, (265) 0 --> (319) 0:NM0, PENB, *, PEGB2
			6'd3 : rdata = 41'b00011100000000001101111111000000010100000;
			// PEs: 43, 44 -> 43
			// srcs: (162, 4)(103) 6, (320) 0 --> (374) 6:NW0, PEGB4, -, NW0
			6'd4 : rdata = 41'b00010010000000001110000100000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 44) begin
	always @(*) begin
		case(address)
			// PEs: 44, 44 -> 45
			// srcs: (1, 0)(49) 4, (104) 7 --> (158) 28:ND0, NW0, *, PENB
			6'd0 : rdata = 41'b00011011000000000100000000000000100000000;
			// PEs: 40, 44 -> 44
			// srcs: (154, 1)(221) -3, (49) 4 --> (267) -12:PEGB0, ND0, *, NI0
			6'd1 : rdata = 41'b00011111000000000110000000010000000000000;
			// PEs: 44, 43 -> 43
			// srcs: (156, 2)(3) 1, (266) 0 --> (320) 0:NM0, PENB, *, PEGB3
			6'd2 : rdata = 41'b00011100000000001101111111000000010110000;
			// PEs: 44, 44 -> 
			// srcs: (157, 3)(3) 1, (267) -12 --> (321) -12:NM0, NI0, *, 
			6'd3 : rdata = 41'b00011100000000001010000000000000000000000;
			// PEs: 44, 44 -> 44
			// srcs: (160, 4)(104) 7, (321) -12 --> (375) 19:NW0, ALU, -, NW0
			6'd4 : rdata = 41'b00010010000000000011111111100100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 45) begin
	always @(*) begin
		case(address)
			// PEs: 45, 45 -> 
			// srcs: (1, 0)(50) 3, (105) 1 --> (159) 3:ND0, NW0, *, 
			6'd0 : rdata = 41'b00011011000000000100000000000000000000000;
			// PEs: 44, 45 -> 41
			// srcs: (4, 1)(158) 28, (159) 3 --> (209) 31:PENB, ALU, +, PEGB1
			6'd1 : rdata = 41'b00001110111111100011111111100000010010000;
			// PEs: 40, 45 -> 46
			// srcs: (155, 2)(221) -3, (50) 3 --> (268) -9:PEGB0, ND0, *, PENB
			6'd2 : rdata = 41'b00011111000000000110000000000000100000000;
			// PEs: 45, 46 -> 45
			// srcs: (164, 3)(105) 1, (322) -9 --> (376) 10:NW0, PEGB6, -, NW0
			6'd3 : rdata = 41'b00010010000000001110000110000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 46) begin
	always @(*) begin
		case(address)
			// PEs: 46, 46 -> 47
			// srcs: (1, 0)(52) 7, (107) 7 --> (161) 49:ND0, NW0, *, PENB
			6'd0 : rdata = 41'b00011011000000000100000000000000100000000;
			// PEs: 40, 46 -> 46
			// srcs: (157, 1)(221) -3, (52) 7 --> (270) -21:PEGB0, ND0, *, NI0
			6'd1 : rdata = 41'b00011111000000000110000000010000000000000;
			// PEs: 46, 45 -> 45
			// srcs: (158, 2)(3) 1, (268) -9 --> (322) -9:NM0, PENB, *, PEGB5
			6'd2 : rdata = 41'b00011100000000001101111111000000011010000;
			// PEs: 46, 46 -> 
			// srcs: (160, 3)(3) 1, (270) -21 --> (324) -21:NM0, NI0, *, 
			6'd3 : rdata = 41'b00011100000000001010000000000000000000000;
			// PEs: 46, 46 -> 46
			// srcs: (163, 4)(107) 7, (324) -21 --> (378) 28:NW0, ALU, -, NW0
			6'd4 : rdata = 41'b00010010000000000011111111100100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 47) begin
	always @(*) begin
		case(address)
			// PEs: 47, 47 -> 
			// srcs: (1, 0)(53) 0, (108) 8 --> (162) 0:ND0, NW0, *, 
			6'd0 : rdata = 41'b00011011000000000100000000000000000000000;
			// PEs: 46, 47 -> 40
			// srcs: (4, 1)(161) 49, (162) 0 --> (212) 49:PENB, ALU, +, PENB
			6'd1 : rdata = 41'b00001110111111100011111111100000100000000;
			// PEs: 40, 47 -> 
			// srcs: (158, 2)(221) -3, (53) 0 --> (271) 0:PEGB0, ND0, *, 
			6'd2 : rdata = 41'b00011111000000000110000000000000000000000;
			// PEs: 47, 47 -> 
			// srcs: (161, 3)(3) 1, (271) 0 --> (325) 0:NM0, ALU, *, 
			6'd3 : rdata = 41'b00011100000000000011111111100000000000000;
			// PEs: 47, 47 -> 47
			// srcs: (164, 4)(108) 8, (325) 0 --> (379) 8:NW0, ALU, -, NW0
			6'd4 : rdata = 41'b00010010000000000011111111100100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 48) begin
	always @(*) begin
		case(address)
			// PEs: 55 -> 24
			// srcs: (3, 4)(139) 49 --> (139) 49:PENB, pass, PUGB3
			6'd0 : rdata = 41'b11000110111111100000000000000000000001011;
			// PEs: 51 -> 16
			// srcs: (6, 0)(119) 18 --> (119) 18:PEGB3, pass, PUGB2
			6'd1 : rdata = 41'b11000111000001100000000000000000000001010;
			// PEs: 52 -> 32
			// srcs: (7, 1)(126) 72 --> (126) 72:PEGB4, pass, PUGB4
			6'd2 : rdata = 41'b11000111000010000000000000000000000001100;
			// PEs: 54 -> 56
			// srcs: (8, 3)(136) 16 --> (136) 16:PEGB6, pass, PUNB
			6'd3 : rdata = 41'b11000111000011000000000000000001000000000;
			// PEs: 50 -> 56
			// srcs: (9, 5)(214) 53 --> (214) 53:PEGB2, pass, PUNB
			6'd4 : rdata = 41'b11000111000001000000000000000001000000000;
			// PEs: 16 -> 49
			// srcs: (14, 2)(183) 3 --> (183) 3:PUGB2, pass, PENB
			6'd5 : rdata = 41'b11000111000001010000000000000000100000000;
			// PEs: 0 -> 48
			// srcs: (22, 6)(169) 74 --> (169) 74:PUGB0, pass, NI0
			6'd6 : rdata = 41'b11000111000000010000000000010000000000000;
			// PEs: 49 -> 32
			// srcs: (23, 9)(184) 21 --> (184) 21:PEGB1, pass, PUGB4
			6'd7 : rdata = 41'b11000111000000100000000000000000000001100;
			// PEs: 16 -> 49
			// srcs: (33, 7)(171) 37 --> (171) 37:PUGB2, pass, PENB
			6'd8 : rdata = 41'b11000111000001010000000000000000100000000;
			// PEs: 48 -> 49
			// srcs: (40, 8)(169) 74 --> (169) 74:NI0, pass, PENB
			6'd9 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 24 -> 49
			// srcs: (52, 10)(178) 305 --> (178) 305:PUGB3, pass, PENB
			6'd10 : rdata = 41'b11000111000001110000000000000000100000000;
			// PEs: 40 -> 49
			// srcs: (60, 11)(191) 281 --> (191) 281:PUNB, pass, PENB
			6'd11 : rdata = 41'b11000110111111110000000000000000100000000;
			// PEs: 49 -> 32
			// srcs: (70, 12)(192) 697 --> (192) 697:PEGB1, pass, PUGB4
			6'd12 : rdata = 41'b11000111000000100000000000000000000001100;
			// PEs: 32 -> 51
			// srcs: (114, 13)(221) -3 --> (221) -3:PUGB4, pass, PEGB3
			6'd13 : rdata = 41'b11000111000010010000000000000000010110000;
			// PEs: 32 -> 52
			// srcs: (121, 14)(221) -3 --> (221) -3:PUGB4, pass, PEGB4
			6'd14 : rdata = 41'b11000111000010010000000000000000011000000;
			// PEs: 32 -> 53
			// srcs: (128, 15)(221) -3 --> (221) -3:PUGB4, pass, PEGB5
			6'd15 : rdata = 41'b11000111000010010000000000000000011010000;
			// PEs: 32 -> 54
			// srcs: (131, 16)(221) -3 --> (221) -3:PUGB4, pass, PEGB6
			6'd16 : rdata = 41'b11000111000010010000000000000000011100000;
			// PEs: 32 -> 55
			// srcs: (134, 17)(221) -3 --> (221) -3:PUGB4, pass, PEGB7
			6'd17 : rdata = 41'b11000111000010010000000000000000011110000;
			// PEs: 32 -> 49
			// srcs: (158, 18)(221) -3 --> (221) -3:PUGB4, pass, PENB
			6'd18 : rdata = 41'b11000111000010010000000000000000100000000;
			// PEs: 32 -> 50
			// srcs: (159, 19)(221) -3 --> (221) -3:PUGB4, pass, PEGB2
			6'd19 : rdata = 41'b11000111000010010000000000000000010100000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 49) begin
	always @(*) begin
		case(address)
			// PEs: 49, 49 -> 50
			// srcs: (1, 0)(55) 5, (110) 7 --> (164) 35:ND0, NW0, *, PENB
			6'd0 : rdata = 41'b00011011000000000100000000000000100000000;
			// PEs: 48, 53 -> 48
			// srcs: (17, 1)(183) 3, (133) 18 --> (184) 21:PENB, PEGB5, +, PEGB0
			6'd1 : rdata = 41'b00001110111111101110000101000000010000000;
			// PEs: 48 -> 
			// srcs: (35, 2)(171) 37 --> (171) 37:PENB, pass, 
			6'd2 : rdata = 41'b11000110111111100000000000000000000000000;
			// PEs: 48, 49 -> 
			// srcs: (42, 3)(169) 74, (171) 37 --> (172) 111:PENB, ALU, +, 
			6'd3 : rdata = 41'b00001110111111100011111111100000000000000;
			// PEs: 49, 48 -> 
			// srcs: (55, 4)(172) 111, (178) 305 --> (179) 416:ALU, PENB, +, 
			6'd4 : rdata = 41'b00001001111111111101111111000000000000000;
			// PEs: 49, 48 -> 48
			// srcs: (65, 5)(179) 416, (191) 281 --> (192) 697:ALU, PENB, +, PEGB0
			6'd5 : rdata = 41'b00001001111111111101111111000000010000000;
			// PEs: 48, 49 -> 50
			// srcs: (160, 6)(221) -3, (55) 5 --> (273) -15:PENB, ND0, *, PENB
			6'd6 : rdata = 41'b00011110111111100110000000000000100000000;
			// PEs: 49, 50 -> 49
			// srcs: (169, 7)(110) 7, (327) -15 --> (381) 22:NW0, PEGB2, -, NW0
			6'd7 : rdata = 41'b00010010000000001110000010000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 50) begin
	always @(*) begin
		case(address)
			// PEs: 50, 50 -> 
			// srcs: (1, 0)(56) 2, (111) 9 --> (165) 18:ND0, NW0, *, 
			6'd0 : rdata = 41'b00011011000000000100000000000000000000000;
			// PEs: 49, 50 -> 48
			// srcs: (4, 1)(164) 35, (165) 18 --> (214) 53:PENB, ALU, +, PEGB0
			6'd1 : rdata = 41'b00001110111111100011111111100000010000000;
			// PEs: 50, 49 -> 49
			// srcs: (163, 3)(3) 1, (273) -15 --> (327) -15:NM0, PENB, *, PEGB1
			6'd2 : rdata = 41'b00011100000000001101111111000000010010000;
			// PEs: 48, 50 -> 51
			// srcs: (164, 2)(221) -3, (56) 2 --> (274) -6:PEGB0, ND0, *, PENB
			6'd3 : rdata = 41'b00011111000000000110000000000000100000000;
			// PEs: 50, 51 -> 50
			// srcs: (173, 4)(111) 9, (328) -6 --> (382) 15:NW0, PEGB3, -, NW0
			6'd4 : rdata = 41'b00010010000000001110000011000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 51) begin
	always @(*) begin
		case(address)
			// PEs: 51, 51 -> 48
			// srcs: (1, 0)(10) 6, (65) 3 --> (119) 18:ND0, NW0, *, PEGB0
			6'd0 : rdata = 41'b00011011000000000100000000000000010000000;
			// PEs: 48, 51 -> 
			// srcs: (119, 1)(221) -3, (10) 6 --> (228) -18:PEGB0, ND0, *, 
			6'd1 : rdata = 41'b00011111000000000110000000000000000000000;
			// PEs: 51, 51 -> 
			// srcs: (122, 2)(3) 1, (228) -18 --> (282) -18:NM0, ALU, *, 
			6'd2 : rdata = 41'b00011100000000000011111111100000000000000;
			// PEs: 51, 51 -> 51
			// srcs: (125, 4)(65) 3, (282) -18 --> (336) 21:NW0, ALU, -, NW0
			6'd3 : rdata = 41'b00010010000000000011111111100100000000000;
			// PEs: 51, 50 -> 50
			// srcs: (167, 3)(3) 1, (274) -6 --> (328) -6:NM0, PENB, *, PEGB2
			6'd4 : rdata = 41'b00011100000000001101111111000000010100000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 52) begin
	always @(*) begin
		case(address)
			// PEs: 52, 52 -> 48
			// srcs: (1, 0)(17) 9, (72) 8 --> (126) 72:ND0, NW0, *, PEGB0
			6'd0 : rdata = 41'b00011011000000000100000000000000010000000;
			// PEs: 48, 52 -> 
			// srcs: (126, 1)(221) -3, (17) 9 --> (235) -27:PEGB0, ND0, *, 
			6'd1 : rdata = 41'b00011111000000000110000000000000000000000;
			// PEs: 52, 52 -> 
			// srcs: (129, 2)(3) 1, (235) -27 --> (289) -27:NM0, ALU, *, 
			6'd2 : rdata = 41'b00011100000000000011111111100000000000000;
			// PEs: 52, 52 -> 52
			// srcs: (132, 3)(72) 8, (289) -27 --> (343) 35:NW0, ALU, -, NW0
			6'd3 : rdata = 41'b00010010000000000011111111100100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 53) begin
	always @(*) begin
		case(address)
			// PEs: 53, 53 -> 49
			// srcs: (1, 0)(24) 6, (79) 3 --> (133) 18:ND0, NW0, *, PEGB1
			6'd0 : rdata = 41'b00011011000000000100000000000000010010000;
			// PEs: 48, 53 -> 
			// srcs: (133, 1)(221) -3, (24) 6 --> (242) -18:PEGB0, ND0, *, 
			6'd1 : rdata = 41'b00011111000000000110000000000000000000000;
			// PEs: 53, 53 -> 
			// srcs: (136, 2)(3) 1, (242) -18 --> (296) -18:NM0, ALU, *, 
			6'd2 : rdata = 41'b00011100000000000011111111100000000000000;
			// PEs: 53, 53 -> 53
			// srcs: (139, 3)(79) 3, (296) -18 --> (350) 21:NW0, ALU, -, NW0
			6'd3 : rdata = 41'b00010010000000000011111111100100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 54) begin
	always @(*) begin
		case(address)
			// PEs: 54, 54 -> 48
			// srcs: (1, 0)(27) 2, (82) 8 --> (136) 16:ND0, NW0, *, PEGB0
			6'd0 : rdata = 41'b00011011000000000100000000000000010000000;
			// PEs: 48, 54 -> 
			// srcs: (136, 1)(221) -3, (27) 2 --> (245) -6:PEGB0, ND0, *, 
			6'd1 : rdata = 41'b00011111000000000110000000000000000000000;
			// PEs: 54, 54 -> 
			// srcs: (139, 2)(3) 1, (245) -6 --> (299) -6:NM0, ALU, *, 
			6'd2 : rdata = 41'b00011100000000000011111111100000000000000;
			// PEs: 54, 54 -> 54
			// srcs: (142, 3)(82) 8, (299) -6 --> (353) 14:NW0, ALU, -, NW0
			6'd3 : rdata = 41'b00010010000000000011111111100100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 55) begin
	always @(*) begin
		case(address)
			// PEs: 55, 55 -> 48
			// srcs: (1, 0)(30) 7, (85) 7 --> (139) 49:ND0, NW0, *, PENB
			6'd0 : rdata = 41'b00011011000000000100000000000000100000000;
			// PEs: 48, 55 -> 
			// srcs: (139, 1)(221) -3, (30) 7 --> (248) -21:PEGB0, ND0, *, 
			6'd1 : rdata = 41'b00011111000000000110000000000000000000000;
			// PEs: 55, 55 -> 
			// srcs: (142, 2)(3) 1, (248) -21 --> (302) -21:NM0, ALU, *, 
			6'd2 : rdata = 41'b00011100000000000011111111100000000000000;
			// PEs: 55, 55 -> 55
			// srcs: (145, 3)(85) 7, (302) -21 --> (356) 28:NW0, ALU, -, NW0
			6'd3 : rdata = 41'b00010010000000000011111111100100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 56) begin
	always @(*) begin
		case(address)
			// PEs: 57 -> 0
			// srcs: (6, 3)(146) 48 --> (146) 48:PEGB1, pass, PUNB
			6'd0 : rdata = 41'b11000111000000100000000000000001000000000;
			// PEs: 58 -> 8
			// srcs: (7, 4)(153) 0 --> (153) 0:PEGB2, pass, PUGB1
			6'd1 : rdata = 41'b11000111000001000000000000000000000001001;
			// PEs: 59 -> 40
			// srcs: (8, 5)(160) 0 --> (160) 0:PEGB3, pass, PUGB5
			6'd2 : rdata = 41'b11000111000001100000000000000000000001101;
			// PEs: 48 -> 56
			// srcs: (10, 1)(136) 16 --> (136) 16:PUNB, pass, NI0
			6'd3 : rdata = 41'b11000110111111110000000000010000000000000;
			// PEs: 16 -> 57
			// srcs: (15, 0)(186) 87 --> (186) 87:PUGB2, pass, PENB
			6'd4 : rdata = 41'b11000111000001010000000000000000100000000;
			// PEs: 56 -> 57
			// srcs: (21, 2)(136) 16 --> (136) 16:NI0, pass, PENB
			6'd5 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 40 -> 57
			// srcs: (22, 6)(212) 49 --> (212) 49:PUGB5, pass, PENB
			6'd6 : rdata = 41'b11000111000010110000000000000000100000000;
			// PEs: 48 -> 57
			// srcs: (23, 7)(214) 53 --> (214) 53:PUNB, pass, PENB
			6'd7 : rdata = 41'b11000110111111110000000000000000100000000;
			// PEs: 57 -> 40
			// srcs: (28, 8)(187) 103 --> (187) 103:PEGB1, pass, PUGB5
			6'd8 : rdata = 41'b11000111000000100000000000000000000001101;
			// PEs: 58 -> 0
			// srcs: (39, 9)(216) 112 --> (216) 112:PEGB2, pass, PUNB
			6'd9 : rdata = 41'b11000111000001000000000000000001000000000;
			// PEs: 32 -> 57
			// srcs: (141, 10)(221) -3 --> (221) -3:PUGB4, pass, PENB
			6'd10 : rdata = 41'b11000111000010010000000000000000100000000;
			// PEs: 32 -> 58
			// srcs: (147, 11)(221) -3 --> (221) -3:PUGB4, pass, PEGB2
			6'd11 : rdata = 41'b11000111000010010000000000000000010100000;
			// PEs: 32 -> 59
			// srcs: (154, 12)(221) -3 --> (221) -3:PUGB4, pass, PEGB3
			6'd12 : rdata = 41'b11000111000010010000000000000000010110000;
			// PEs: 32 -> 60
			// srcs: (157, 13)(221) -3 --> (221) -3:PUGB4, pass, PEGB4
			6'd13 : rdata = 41'b11000111000010010000000000000000011000000;
			// PEs: 32 -> 61
			// srcs: (160, 14)(221) -3 --> (221) -3:PUGB4, pass, PEGB5
			6'd14 : rdata = 41'b11000111000010010000000000000000011010000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 57) begin
	always @(*) begin
		case(address)
			// PEs: 57, 57 -> 56
			// srcs: (1, 0)(37) 8, (92) 6 --> (146) 48:ND0, NW0, *, PEGB0
			6'd0 : rdata = 41'b00011011000000000100000000000000010000000;
			// PEs: 56 -> 
			// srcs: (17, 1)(186) 87 --> (186) 87:PENB, pass, 
			6'd1 : rdata = 41'b11000110111111100000000000000000000000000;
			// PEs: 57, 56 -> 56
			// srcs: (23, 2)(186) 87, (136) 16 --> (187) 103:ALU, PENB, +, PEGB0
			6'd2 : rdata = 41'b00001001111111111101111111000000010000000;
			// PEs: 56, 60 -> 57
			// srcs: (24, 3)(212) 49, (163) 6 --> (213) 55:PENB, PEGB4, +, NI0
			6'd3 : rdata = 41'b00001110111111101110000100010000000000000;
			// PEs: 56, 61 -> 58
			// srcs: (25, 4)(214) 53, (166) 4 --> (215) 57:PENB, PEGB5, +, PENB
			6'd4 : rdata = 41'b00001110111111101110000101000000100000000;
			// PEs: 57 -> 58
			// srcs: (32, 5)(213) 55 --> (213) 55:NI0, pass, PENB
			6'd5 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 56, 57 -> 58
			// srcs: (143, 6)(221) -3, (37) 8 --> (255) -24:PENB, ND0, *, PENB
			6'd6 : rdata = 41'b00011110111111100110000000000000100000000;
			// PEs: 57, 58 -> 57
			// srcs: (152, 7)(92) 6, (309) -24 --> (363) 30:NW0, PEGB2, -, NW0
			6'd7 : rdata = 41'b00010010000000001110000010000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 58) begin
	always @(*) begin
		case(address)
			// PEs: 58, 58 -> 56
			// srcs: (1, 0)(44) 8, (99) 0 --> (153) 0:ND0, NW0, *, PEGB0
			6'd0 : rdata = 41'b00011011000000000100000000000000010000000;
			// PEs: 57 -> 
			// srcs: (27, 1)(215) 57 --> (215) 57:PENB, pass, 
			6'd1 : rdata = 41'b11000110111111100000000000000000000000000;
			// PEs: 57, 58 -> 56
			// srcs: (34, 2)(213) 55, (215) 57 --> (216) 112:PENB, ALU, +, PEGB0
			6'd2 : rdata = 41'b00001110111111100011111111100000010000000;
			// PEs: 58, 57 -> 57
			// srcs: (146, 4)(3) 1, (255) -24 --> (309) -24:NM0, PENB, *, PEGB1
			6'd3 : rdata = 41'b00011100000000001101111111000000010010000;
			// PEs: 56, 58 -> 59
			// srcs: (152, 3)(221) -3, (44) 8 --> (262) -24:PEGB0, ND0, *, PENB
			6'd4 : rdata = 41'b00011111000000000110000000000000100000000;
			// PEs: 58, 59 -> 58
			// srcs: (161, 5)(99) 0, (316) -24 --> (370) 24:NW0, PEGB3, -, NW0
			6'd5 : rdata = 41'b00010010000000001110000011000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 59) begin
	always @(*) begin
		case(address)
			// PEs: 59, 59 -> 56
			// srcs: (1, 0)(51) 0, (106) 5 --> (160) 0:ND0, NW0, *, PEGB0
			6'd0 : rdata = 41'b00011011000000000100000000000000010000000;
			// PEs: 59, 58 -> 58
			// srcs: (155, 2)(3) 1, (262) -24 --> (316) -24:NM0, PENB, *, PEGB2
			6'd1 : rdata = 41'b00011100000000001101111111000000010100000;
			// PEs: 56, 59 -> 
			// srcs: (159, 1)(221) -3, (51) 0 --> (269) 0:PEGB0, ND0, *, 
			6'd2 : rdata = 41'b00011111000000000110000000000000000000000;
			// PEs: 59, 59 -> 
			// srcs: (162, 3)(3) 1, (269) 0 --> (323) 0:NM0, ALU, *, 
			6'd3 : rdata = 41'b00011100000000000011111111100000000000000;
			// PEs: 59, 59 -> 59
			// srcs: (165, 4)(106) 5, (323) 0 --> (377) 5:NW0, ALU, -, NW0
			6'd4 : rdata = 41'b00010010000000000011111111100100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 60) begin
	always @(*) begin
		case(address)
			// PEs: 60, 60 -> 57
			// srcs: (1, 0)(54) 6, (109) 1 --> (163) 6:ND0, NW0, *, PEGB1
			6'd0 : rdata = 41'b00011011000000000100000000000000010010000;
			// PEs: 56, 60 -> 
			// srcs: (162, 1)(221) -3, (54) 6 --> (272) -18:PEGB0, ND0, *, 
			6'd1 : rdata = 41'b00011111000000000110000000000000000000000;
			// PEs: 60, 60 -> 
			// srcs: (165, 2)(3) 1, (272) -18 --> (326) -18:NM0, ALU, *, 
			6'd2 : rdata = 41'b00011100000000000011111111100000000000000;
			// PEs: 60, 60 -> 60
			// srcs: (168, 3)(109) 1, (326) -18 --> (380) 19:NW0, ALU, -, NW0
			6'd3 : rdata = 41'b00010010000000000011111111100100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 61) begin
	always @(*) begin
		case(address)
			// PEs: 61, 61 -> 57
			// srcs: (1, 0)(57) 4, (112) 1 --> (166) 4:ND0, NW0, *, PEGB1
			6'd0 : rdata = 41'b00011011000000000100000000000000010010000;
			// PEs: 56, 61 -> 62
			// srcs: (165, 1)(221) -3, (57) 4 --> (275) -12:PEGB0, ND0, *, PENB
			6'd1 : rdata = 41'b00011111000000000110000000000000100000000;
			// PEs: 61, 62 -> 61
			// srcs: (174, 2)(112) 1, (329) -12 --> (383) 13:NW0, PEGB6, -, NW0
			6'd2 : rdata = 41'b00010010000000001110000110000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 62) begin
	always @(*) begin
		case(address)
			// PEs: 62, 61 -> 61
			// srcs: (168, 0)(3) 1, (275) -12 --> (329) -12:NM0, PENB, *, PEGB5
			6'd0 : rdata = 41'b00011100000000001101111111000000011010000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 63) begin
	always @(*) begin
		case(address)
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

endgenerate
/*****************************************************************************/
endmodule
