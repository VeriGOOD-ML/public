`timescale 1ns/1ps

module ROM_ASIC #(
// Parameters
    parameter   DATA_WIDTH          = 16,
    parameter   ADDR_WIDTH          = 7,
    parameter   INIT                = "weight.txt",
    parameter   TYPE                = "block",
    parameter   ROM_DEPTH           = 1<<ADDR_WIDTH
) (
// Port Declarations
    input  wire                         CLK,
    input  wire                         RESET,
    input  wire  [ADDR_WIDTH-1:0]       ADDRESS,
    input  wire                         ENABLE,
    output reg   [DATA_WIDTH-1:0]       DATA_OUT,
    output reg                          DATA_OUT_VALID
);

// ******************************************************************
// Internal variables
// ******************************************************************

  localparam DEPTH = ROM_DEPTH;

  reg     [DATA_WIDTH-1:0]        rdata;
  wire     [ADDR_WIDTH-1:0]        address;

  assign address = ADDRESS;


  // `include "instructions.v"   // TODO
  always @(*) begin
	case(address)
/*****************************************************************************************/
//
// read [True, False, False, False]
// ['x(0,)', 'x(1,)', 'x(2,)', 'x(3,)', 'x(88,)', 'x(89,)', 'x(91,)', 'x(92,)', 'x(177,)', 'x(178,)', 'x(179,)', 'x(180,)', 'x(174,)', 'x(181,)', 'x(184,)', 'x(187,)']
// Data values: [0, -3, -1, -3, 1, -3, -2, -1, 1, 0, 1, 1, 0, 1, 0, 2]
// Dest PEs: [1, 2, 3, 4, 10, 11, 12, 13, 19, 20, 21, 22, 28, 29, 30, 31]
7'd0: rdata =    56'b00000000000000000000000000000000000000000000000000000001;
//
// shift amount: 15, Lanes IDs: [1, 2, 3, 4]
7'd1: rdata =    56'b00000000000000000000000000000000000100100100100001011111;
//
// read [True, False, False, False]
// ['x(4,)', 'x(5,)', 'x(7,)', 'x(8,)', 'x(88,)', 'x(89,)', 'x(91,)', 'x(92,)', 'x(177,)', 'x(178,)', 'x(179,)', 'x(180,)', 'x(174,)', 'x(181,)', 'x(184,)', 'x(187,)']
// Data values: [-2, 2, -1, 2, 1, -3, -2, -1, 1, 0, 1, 1, 0, 1, 0, 2]
// Dest PEs: [5, 6, 7, 9, 10, 11, 12, 13, 19, 20, 21, 22, 28, 29, 30, 31]
7'd2: rdata =    56'b00000000000000000000000000000000000000000000000000000001;
//
// shift amount: 10, Lanes IDs: [9]
7'd3: rdata =    56'b00000000000000000000100000000000000000000000000001011010;
//
// shift amount: 11, Lanes IDs: [5, 6, 7]
7'd4: rdata =    56'b00000000000000000000000000100100100000000000000001011011;
//
// read [True, True, False, False]
// ['x(10,)', 'x(11,)', 'x(13,)', 'x(14,)', 'x(88,)', 'x(89,)', 'x(91,)', 'x(92,)', 'x(177,)', 'x(178,)', 'x(179,)', 'x(180,)', 'x(174,)', 'x(181,)', 'x(184,)', 'x(187,)']
// Data values: [-3, 1, -1, 0, 1, -3, -2, -1, 1, 0, 1, 1, 0, 1, 0, 2]
// Dest PEs: [10, 11, 12, 13, 10, 11, 12, 13, 19, 20, 21, 22, 28, 29, 30, 31]
7'd5: rdata =    56'b00000000000000000000000000000000000000000000000000000011;
//
// shift amount: 6, Lanes IDs: [10, 11, 12, 13]
7'd6: rdata =    56'b00000000100100100100000000000000000000000000000001010110;
//
// shift amount: 10, Lanes IDs: [10, 11, 12, 13]
7'd7: rdata =    56'b00000000100100100100000000000000000000000000000001011010;
//
// read [True, True, False, False]
// ['x(16,)', 'x(17,)', 'x(19,)', 'x(20,)', 'x(94,)', 'x(95,)', 'x(97,)', 'x(98,)', 'x(177,)', 'x(178,)', 'x(179,)', 'x(180,)', 'x(174,)', 'x(181,)', 'x(184,)', 'x(187,)']
// Data values: [-1, 0, 1, -2, 0, 1, 0, 1, 1, 0, 1, 1, 0, 1, 0, 2]
// Dest PEs: [14, 15, 17, 18, 14, 15, 17, 18, 19, 20, 21, 22, 28, 29, 30, 31]
7'd8: rdata =    56'b00000000000000000000000000000000000000000000000000000011;
//
// shift amount: 1, Lanes IDs: [1, 2]
7'd9: rdata =    56'b00000000000000000000000000000000000000001101100001010001;
//
// shift amount: 2, Lanes IDs: [14, 15]
7'd10: rdata =   56'b00100100000000000000000000000000000000000000000001010010;
//
// shift amount: 5, Lanes IDs: [1, 2]
7'd11: rdata =   56'b00000000000000000000000000000000000000001101100001010101;
//
// shift amount: 6, Lanes IDs: [14, 15]
7'd12: rdata =   56'b00100100000000000000000000000000000000000000000001010110;
//
// read [True, True, True, False]
// ['x(22,)', 'x(23,)', 'x(25,)', 'x(26,)', 'x(100,)', 'x(101,)', 'x(102,)', 'x(103,)', 'x(177,)', 'x(178,)', 'x(179,)', 'x(180,)', 'x(174,)', 'x(181,)', 'x(184,)', 'x(187,)']
// Data values: [-2, 0, -3, 2, 1, 1, -2, 2, 1, 0, 1, 1, 0, 1, 0, 2]
// Dest PEs: [19, 20, 21, 22, 19, 20, 21, 22, 19, 20, 21, 22, 28, 29, 30, 31]
7'd13: rdata =   56'b00000000000000000000000000000000000000000000000000000111;
//
// shift amount: 13, Lanes IDs: [3, 4, 5, 6]
7'd14: rdata =   56'b00000000000000000000000000001101101101100000000001011101;
//
// shift amount: 1, Lanes IDs: [3, 4, 5, 6]
7'd15: rdata =   56'b00000000000000000000000000001101101101100000000001010001;
//
// shift amount: 5, Lanes IDs: [3, 4, 5, 6]
7'd16: rdata =   56'b00000000000000000000000000001101101101100000000001010101;
//
// read [True, True, True, False]
// ['x(27,)', 'x(28,)', 'x(29,)', 'x(30,)', 'x(104,)', 'x(105,)', 'x(107,)', 'x(108,)', 'x(182,)', 'x(183,)', 'x(185,)', 'x(186,)', 'x(174,)', 'x(181,)', 'x(184,)', 'x(187,)']
// Data values: [0, -1, 0, 2, 1, 2, 1, 2, 0, 2, -1, -3, 0, 1, 0, 2]
// Dest PEs: [23, 25, 26, 27, 23, 25, 26, 27, 23, 25, 26, 27, 28, 29, 30, 31]
7'd17: rdata =   56'b00000000000000000000000000000000000000000000000000000111;
//
// shift amount: 8, Lanes IDs: [9, 10, 11]
7'd18: rdata =   56'b00000000000001101101100000000000000000000000000001011000;
//
// shift amount: 9, Lanes IDs: [7]
7'd19: rdata =   56'b00000000000000000000000001100000000000000000000001011001;
//
// shift amount: 12, Lanes IDs: [9, 10, 11]
7'd20: rdata =   56'b00000000000001101101100000000000000000000000000001011100;
//
// shift amount: 0, Lanes IDs: [9, 10, 11]
7'd21: rdata =   56'b00000000000001101101100000000000000000000000000001010000;
//
// shift amount: 13, Lanes IDs: [7]
7'd22: rdata =   56'b00000000000000000000000001100000000000000000000001011101;
//
// shift amount: 1, Lanes IDs: [7]
7'd23: rdata =   56'b00000000000000000000000001100000000000000000000001010001;
//
// read [True, True, True, True]
// ['x(32,)', 'x(33,)', 'x(35,)', 'x(36,)', 'x(110,)', 'x(111,)', 'x(113,)', 'x(114,)', 'x(188,)', 'x(189,)', 'x(191,)', 'x(192,)', 'x(174,)', 'x(181,)', 'x(184,)', 'x(187,)']
// Data values: [-2, 0, -3, 2, -3, -1, -2, -1, 1, 2, -3, 1, 0, 1, 0, 2]
// Dest PEs: [28, 29, 30, 31, 28, 29, 30, 31, 28, 29, 30, 31, 28, 29, 30, 31]
7'd24: rdata =   56'b00000000000000000000000000000000000000000000000000001111;
//
// shift amount: 4, Lanes IDs: [12, 13, 14, 15]
7'd25: rdata =   56'b01101101101100000000000000000000000000000000000001010100;
//
// shift amount: 8, Lanes IDs: [12, 13, 14, 15]
7'd26: rdata =   56'b01101101101100000000000000000000000000000000000001011000;
//
// shift amount: 12, Lanes IDs: [12, 13, 14, 15]
7'd27: rdata =   56'b01101101101100000000000000000000000000000000000001011100;
//
// shift amount: 0, Lanes IDs: [12, 13, 14, 15]
7'd28: rdata =   56'b01101101101100000000000000000000000000000000000001010000;
//
// read [True, True, True, True]
// ['x(38,)', 'x(39,)', 'x(41,)', 'x(42,)', 'x(116,)', 'x(117,)', 'x(119,)', 'x(120,)', 'x(194,)', 'x(195,)', 'x(197,)', 'x(198,)', 'x(190,)', 'x(193,)', 'x(196,)', 'x(199,)']
// Data values: [-2, 1, 0, 2, 1, 0, 2, -3, 1, 0, 2, 0, 0, -3, 0, 2]
// Dest PEs: [33, 34, 35, 36, 33, 34, 35, 36, 33, 34, 35, 36, 33, 34, 35, 36]
7'd29: rdata =   56'b00000000000000000000000000000000000000000000000000001111;
//
// shift amount: 15, Lanes IDs: [1, 2, 3, 4]
7'd30: rdata =   56'b00000000000000000000000000000000010110110110100001011111;
//
// shift amount: 3, Lanes IDs: [1, 2, 3, 4]
7'd31: rdata =   56'b00000000000000000000000000000000010110110110100001010011;
//
// shift amount: 7, Lanes IDs: [1, 2, 3, 4]
7'd32: rdata =   56'b00000000000000000000000000000000010110110110100001010111;
//
// shift amount: 11, Lanes IDs: [1, 2, 3, 4]
7'd33: rdata =   56'b00000000000000000000000000000000010110110110100001011011;
//
// read [True, True, True, True]
// ['x(44,)', 'x(45,)', 'x(47,)', 'x(48,)', 'x(122,)', 'x(123,)', 'x(125,)', 'x(126,)', 'x(6,)', 'x(9,)', 'x(12,)', 'x(15,)', 'y', None, None, None]
// Data values: [-3, 1, 2, 1, -3, -3, 1, 2, -3, 2, -3, -3, -1, None, None, None]
// Dest PEs: [37, 38, 39, 41, 37, 38, 39, 41, 37, 38, 39, 41, 37, None, None, None]
7'd34: rdata =   56'b00000000000000000000000000000000000000000000000000001111;
//
// shift amount: 10, Lanes IDs: [9]
7'd35: rdata =   56'b00000000000000000010100000000000000000000000000001011010;
//
// shift amount: 11, Lanes IDs: [5, 6, 7]
7'd36: rdata =   56'b00000000000000000000000010110110100000000000000001011011;
//
// shift amount: 14, Lanes IDs: [9]
7'd37: rdata =   56'b00000000000000000010100000000000000000000000000001011110;
//
// shift amount: 2, Lanes IDs: [9]
7'd38: rdata =   56'b00000000000000000010100000000000000000000000000001010010;
//
// shift amount: 15, Lanes IDs: [5, 6, 7]
7'd39: rdata =   56'b00000000000000000000000010110110100000000000000001011111;
//
// shift amount: 3, Lanes IDs: [5, 6, 7]
7'd40: rdata =   56'b00000000000000000000000010110110100000000000000001010011;
//
// shift amount: 7, Lanes IDs: [5]
7'd41: rdata =   56'b00000000000000000000000000000010100000000000000001010111;
//
// read [True, True, True, False]
// ['x(50,)', 'x(51,)', 'x(52,)', 'x(53,)', 'x(127,)', 'x(128,)', 'x(129,)', 'x(130,)', 'x(18,)', 'x(21,)', 'x(24,)', 'x(31,)', None, None, None, None]
// Data values: [2, 0, -3, -1, 1, -1, -3, -3, 2, 1, 1, 1, None, None, None, None]
// Dest PEs: [42, 43, 44, 45, 42, 43, 44, 45, 42, 43, 44, 45, None, None, None, None]
7'd42: rdata =   56'b00000000000000000000000000000000000000000000000000000111;
//
// shift amount: 6, Lanes IDs: [10, 11, 12, 13]
7'd43: rdata =   56'b00000010110110110100000000000000000000000000000001010110;
//
// shift amount: 10, Lanes IDs: [10, 11, 12, 13]
7'd44: rdata =   56'b00000010110110110100000000000000000000000000000001011010;
//
// shift amount: 14, Lanes IDs: [10, 11, 12, 13]
7'd45: rdata =   56'b00000010110110110100000000000000000000000000000001011110;
//
// read [True, True, True, False]
// ['x(54,)', 'x(55,)', 'x(57,)', 'x(58,)', 'x(132,)', 'x(133,)', 'x(135,)', 'x(136,)', 'x(34,)', 'x(37,)', 'x(40,)', 'x(43,)', None, None, None, None]
// Data values: [1, -3, 1, -3, 0, -1, 0, 1, 0, -2, -2, -2, None, None, None, None]
// Dest PEs: [46, 47, 49, 50, 46, 47, 49, 50, 46, 47, 49, 50, None, None, None, None]
7'd46: rdata =   56'b00000000000000000000000000000000000000000000000000000111;
//
// shift amount: 1, Lanes IDs: [1, 2]
7'd47: rdata =   56'b00000000000000000000000000000000000000011111100001010001;
//
// shift amount: 2, Lanes IDs: [14, 15]
7'd48: rdata =   56'b10110100000000000000000000000000000000000000000001010010;
//
// shift amount: 5, Lanes IDs: [1, 2]
7'd49: rdata =   56'b00000000000000000000000000000000000000011111100001010101;
//
// shift amount: 6, Lanes IDs: [14, 15]
7'd50: rdata =   56'b10110100000000000000000000000000000000000000000001010110;
//
// shift amount: 9, Lanes IDs: [1, 2]
7'd51: rdata =   56'b00000000000000000000000000000000000000011111100001011001;
//
// shift amount: 10, Lanes IDs: [14, 15]
7'd52: rdata =   56'b10110100000000000000000000000000000000000000000001011010;
//
// read [True, True, True, False]
// ['x(60,)', 'x(61,)', 'x(63,)', 'x(64,)', 'x(138,)', 'x(139,)', 'x(141,)', 'x(142,)', 'x(46,)', 'x(49,)', 'x(56,)', 'x(59,)', None, None, None, None]
// Data values: [-1, 2, -3, 0, -1, 0, -3, 0, -2, -2, 0, -2, None, None, None, None]
// Dest PEs: [51, 52, 53, 54, 51, 52, 53, 54, 51, 52, 53, 54, None, None, None, None]
7'd53: rdata =   56'b00000000000000000000000000000000000000000000000000000111;
//
// shift amount: 13, Lanes IDs: [3, 4, 5, 6]
7'd54: rdata =   56'b00000000000000000000000000011111111111100000000001011101;
//
// shift amount: 1, Lanes IDs: [3, 4, 5, 6]
7'd55: rdata =   56'b00000000000000000000000000011111111111100000000001010001;
//
// shift amount: 5, Lanes IDs: [3, 4, 5, 6]
7'd56: rdata =   56'b00000000000000000000000000011111111111100000000001010101;
//
// read [True, True, True, False]
// ['x(66,)', 'x(67,)', 'x(69,)', 'x(70,)', 'x(144,)', 'x(145,)', 'x(147,)', 'x(148,)', 'x(62,)', 'x(65,)', 'x(68,)', 'x(71,)', None, None, None, None]
// Data values: [-1, 0, -3, -1, -3, -2, 2, -3, -1, -1, 1, 2, None, None, None, None]
// Dest PEs: [55, 57, 58, 59, 55, 57, 58, 59, 55, 57, 58, 59, None, None, None, None]
7'd57: rdata =   56'b00000000000000000000000000000000000000000000000000000111;
//
// shift amount: 8, Lanes IDs: [9, 10, 11]
7'd58: rdata =   56'b00000000000011111111100000000000000000000000000001011000;
//
// shift amount: 9, Lanes IDs: [7]
7'd59: rdata =   56'b00000000000000000000000011100000000000000000000001011001;
//
// shift amount: 12, Lanes IDs: [9, 10, 11]
7'd60: rdata =   56'b00000000000011111111100000000000000000000000000001011100;
//
// shift amount: 0, Lanes IDs: [9, 10, 11]
7'd61: rdata =   56'b00000000000011111111100000000000000000000000000001010000;
//
// shift amount: 13, Lanes IDs: [7]
7'd62: rdata =   56'b00000000000000000000000011100000000000000000000001011101;
//
// shift amount: 1, Lanes IDs: [7]
7'd63: rdata =   56'b00000000000000000000000011100000000000000000000001010001;
//
// read [True, True, True, False]
// ['x(72,)', 'x(73,)', 'x(75,)', 'x(76,)', 'x(150,)', 'x(151,)', 'x(152,)', 'x(153,)', 'x(74,)', 'x(81,)', 'x(84,)', 'x(87,)', None, None, None, None]
// Data values: [0, -3, -2, -1, 2, -3, -2, 0, -2, -2, 2, -2, None, None, None, None]
// Dest PEs: [60, 61, 62, 63, 60, 61, 62, 63, 60, 61, 62, 63, None, None, None, None]
7'd64: rdata =   56'b00000000000000000000000000000000000000000000000000000111;
//
// shift amount: 4, Lanes IDs: [12, 13, 14, 15]
7'd65: rdata =   56'b11111111111100000000000000000000000000000000000001010100;
//
// shift amount: 8, Lanes IDs: [12, 13, 14, 15]
7'd66: rdata =   56'b11111111111100000000000000000000000000000000000001011000;
//
// shift amount: 12, Lanes IDs: [12, 13, 14, 15]
7'd67: rdata =   56'b11111111111100000000000000000000000000000000000001011100;
//
// read [True, True, True, False]
// ['x(77,)', 'x(78,)', 'x(79,)', 'x(80,)', 'x(154,)', 'x(155,)', 'x(157,)', 'x(158,)', 'x(90,)', 'x(93,)', 'x(96,)', 'x(99,)', None, None, None, None]
// Data values: [0, -2, -2, 2, -1, -2, 2, -1, -1, -2, -3, -2, None, None, None, None]
// Dest PEs: [1, 2, 3, 4, 1, 2, 3, 4, 1, 2, 3, 4, None, None, None, None]
7'd68: rdata =   56'b00000000000000000000000000000000000000000000000000000111;
//
// shift amount: 15, Lanes IDs: [1, 2, 3, 4]
7'd69: rdata =   56'b00000000000000000000000000000000000100100100100001011111;
//
// shift amount: 3, Lanes IDs: [1, 2, 3, 4]
7'd70: rdata =   56'b00000000000000000000000000000000000100100100100001010011;
//
// shift amount: 7, Lanes IDs: [1, 2, 3, 4]
7'd71: rdata =   56'b00000000000000000000000000000000000100100100100001010111;
//
// read [True, True, True, False]
// ['x(82,)', 'x(83,)', 'x(85,)', 'x(86,)', 'x(160,)', 'x(161,)', 'x(163,)', 'x(164,)', 'x(106,)', 'x(109,)', 'x(112,)', 'x(115,)', None, None, None, None]
// Data values: [2, 0, 2, -3, -2, -3, -1, -1, 2, -2, -2, -1, None, None, None, None]
// Dest PEs: [5, 6, 7, 9, 5, 6, 7, 9, 5, 6, 7, 9, None, None, None, None]
7'd72: rdata =   56'b00000000000000000000000000000000000000000000000000000111;
//
// shift amount: 10, Lanes IDs: [9]
7'd73: rdata =   56'b00000000000000000000100000000000000000000000000001011010;
//
// shift amount: 11, Lanes IDs: [5, 6, 7]
7'd74: rdata =   56'b00000000000000000000000000100100100000000000000001011011;
//
// shift amount: 14, Lanes IDs: [9]
7'd75: rdata =   56'b00000000000000000000100000000000000000000000000001011110;
//
// shift amount: 2, Lanes IDs: [9]
7'd76: rdata =   56'b00000000000000000000100000000000000000000000000001010010;
//
// shift amount: 15, Lanes IDs: [5, 6, 7]
7'd77: rdata =   56'b00000000000000000000000000100100100000000000000001011111;
//
// shift amount: 3, Lanes IDs: [5, 6, 7]
7'd78: rdata =   56'b00000000000000000000000000100100100000000000000001010011;
//
// read [False, True, True, False]
// [None, None, None, None, 'x(166,)', 'x(167,)', 'x(169,)', 'x(170,)', 'x(118,)', 'x(121,)', 'x(124,)', 'x(131,)', None, None, None, None]
// Data values: [None, None, None, None, -2, 1, -3, 0, -3, -1, -3, 2, None, None, None, None]
// Dest PEs: [None, None, None, None, 10, 11, 12, 13, 10, 11, 12, 13, None, None, None, None]
7'd79: rdata =   56'b00000000000000000000000000000000000000000000000000000110;
//
// shift amount: 10, Lanes IDs: [10, 11, 12, 13]
7'd80: rdata =   56'b00000000100100100100000000000000000000000000000001011010;
//
// shift amount: 14, Lanes IDs: [10, 11, 12, 13]
7'd81: rdata =   56'b00000000100100100100000000000000000000000000000001011110;
//
// read [False, True, True, False]
// [None, None, None, None, 'x(172,)', 'x(173,)', 'x(175,)', 'x(176,)', 'x(134,)', 'x(137,)', 'x(140,)', 'x(143,)', None, None, None, None]
// Data values: [None, None, None, None, -2, -2, 2, -1, -2, -3, 1, 0, None, None, None, None]
// Dest PEs: [None, None, None, None, 14, 15, 17, 18, 14, 15, 17, 18, None, None, None, None]
7'd82: rdata =   56'b00000000000000000000000000000000000000000000000000000110;
//
// shift amount: 5, Lanes IDs: [1, 2]
7'd83: rdata =   56'b00000000000000000000000000000000000000001101100001010101;
//
// shift amount: 9, Lanes IDs: [1, 2]
7'd84: rdata =   56'b00000000000000000000000000000000000000001101100001011001;
//
// shift amount: 6, Lanes IDs: [14, 15]
7'd85: rdata =   56'b00100100000000000000000000000000000000000000000001010110;
//
// shift amount: 10, Lanes IDs: [14, 15]
7'd86: rdata =   56'b00100100000000000000000000000000000000000000000001011010;
//
// read [False, False, True, False]
// [None, None, None, None, None, None, None, None, 'x(146,)', 'x(149,)', 'x(156,)', 'x(159,)', None, None, None, None]
// Data values: [None, None, None, None, None, None, None, None, -3, 0, 2, 2, None, None, None, None]
// Dest PEs: [None, None, None, None, None, None, None, None, 19, 20, 21, 22, None, None, None, None]
7'd87: rdata =   56'b00000000000000000000000000000000000000000000000000000100;
//
// shift amount: 5, Lanes IDs: [3, 4, 5, 6]
7'd88: rdata =   56'b00000000000000000000000000001101101101100000000001010101;
//
// read [False, False, True, False]
// [None, None, None, None, None, None, None, None, 'x(162,)', 'x(165,)', 'x(168,)', 'x(171,)', None, None, None, None]
// Data values: [None, None, None, None, None, None, None, None, 1, -1, 1, -1, None, None, None, None]
// Dest PEs: [None, None, None, None, None, None, None, None, 23, 25, 26, 27, None, None, None, None]
7'd89: rdata =   56'b00000000000000000000000000000000000000000000000000000100;
//
// shift amount: 0, Lanes IDs: [9, 10, 11]
7'd90: rdata =   56'b00000000000001101101100000000000000000000000000001010000;
//
// shift amount: 1, Lanes IDs: [7]
7'd91: rdata =   56'b00000000000000000000000001100000000000000000000001010001;
//
// wfi
7'd92: rdata =   56'b00000000000000000000000000000000000000000000000001100000;
//
// loop
7'd93: rdata =   56'b00000000000000000000000000000000000000000000000001110000;/****************************************************************************************/
default: rdata = 56'b00000000000000000000000000000000000000000000000001110000;

	endcase
	end

    //reg     [ADDR_WIDTH-1:0]        address;

// ******************************************************************
// Read Logic
// ******************************************************************

    always @ (posedge CLK)
    begin : READ_VALID
        if (RESET) begin
            DATA_OUT_VALID <= 1'b0;
        end else if (ENABLE) begin
            DATA_OUT_VALID <= 1'b1;
        end
    end



 always @(posedge CLK) begin
    if (ENABLE)
        DATA_OUT <= rdata;
end

endmodule
