`timescale 1ns/1ps

module ROM_ASIC #(
// Parameters
    parameter   DATA_WIDTH          = 16,
    parameter   ADDR_WIDTH          = 9,
    parameter   INIT                = "weight.txt",
    parameter   TYPE                = "block",
    parameter   ROM_DEPTH           = 1<<ADDR_WIDTH
) (
// Port Declarations
    input  wire                         CLK,
    input  wire                         RESET,
    input  wire  [ADDR_WIDTH-1:0]       ADDRESS,
    input  wire                         ENABLE,
    output reg   [DATA_WIDTH-1:0]       DATA_OUT,
    output reg                          DATA_OUT_VALID
);

// ******************************************************************
// Internal variables
// ******************************************************************

  localparam DEPTH = ROM_DEPTH;

  reg     [DATA_WIDTH-1:0]        rdata;
  wire     [ADDR_WIDTH-1:0]        address;

  assign address = ADDRESS;


  // `include "instructions.v"   // TODO
  always @(*) begin
	case(address)
/*****************************************************************************************/
//
// read [True, False, False, False]
// ['x(0,)', 'x(1,)', 'x(2,)', 'x(3,)', 'x(92,)', 'x(93,)', 'x(95,)', 'x(96,)', 'x(184,)', 'x(185,)', 'x(187,)', 'x(188,)', 'x(276,)', 'x(277,)', 'x(279,)', 'x(280,)']
// Data values: [-3, -1, 0, 0, -1, 2, -3, 0, 2, 0, -2, 1, 0, -3, 1, -2]
// Dest PEs: [1, 2, 3, 4, 10, 11, 12, 13, 19, 20, 21, 22, 28, 29, 30, 31]
9'd0: rdata =    56'b00000000000000000000000000000000000000000000000000000001;
//
// shift amount: 15, Lanes IDs: [1, 2, 3, 4]
9'd1: rdata =    56'b00000000000000000000000000000000000100100100100001011111;
//
// read [True, False, False, False]
// ['x(4,)', 'x(5,)', 'x(7,)', 'x(8,)', 'x(92,)', 'x(93,)', 'x(95,)', 'x(96,)', 'x(184,)', 'x(185,)', 'x(187,)', 'x(188,)', 'x(276,)', 'x(277,)', 'x(279,)', 'x(280,)']
// Data values: [2, 2, 2, -1, -1, 2, -3, 0, 2, 0, -2, 1, 0, -3, 1, -2]
// Dest PEs: [5, 6, 7, 9, 10, 11, 12, 13, 19, 20, 21, 22, 28, 29, 30, 31]
9'd2: rdata =    56'b00000000000000000000000000000000000000000000000000000001;
//
// shift amount: 10, Lanes IDs: [9]
9'd3: rdata =    56'b00000000000000000000100000000000000000000000000001011010;
//
// shift amount: 11, Lanes IDs: [5, 6, 7]
9'd4: rdata =    56'b00000000000000000000000000100100100000000000000001011011;
//
// read [True, True, False, False]
// ['x(10,)', 'x(11,)', 'x(13,)', 'x(14,)', 'x(92,)', 'x(93,)', 'x(95,)', 'x(96,)', 'x(184,)', 'x(185,)', 'x(187,)', 'x(188,)', 'x(276,)', 'x(277,)', 'x(279,)', 'x(280,)']
// Data values: [2, 2, -2, -3, -1, 2, -3, 0, 2, 0, -2, 1, 0, -3, 1, -2]
// Dest PEs: [10, 11, 12, 13, 10, 11, 12, 13, 19, 20, 21, 22, 28, 29, 30, 31]
9'd5: rdata =    56'b00000000000000000000000000000000000000000000000000000011;
//
// shift amount: 6, Lanes IDs: [10, 11, 12, 13]
9'd6: rdata =    56'b00000000100100100100000000000000000000000000000001010110;
//
// shift amount: 10, Lanes IDs: [10, 11, 12, 13]
9'd7: rdata =    56'b00000000100100100100000000000000000000000000000001011010;
//
// read [True, True, False, False]
// ['x(16,)', 'x(17,)', 'x(19,)', 'x(20,)', 'x(98,)', 'x(99,)', 'x(100,)', 'x(101,)', 'x(184,)', 'x(185,)', 'x(187,)', 'x(188,)', 'x(276,)', 'x(277,)', 'x(279,)', 'x(280,)']
// Data values: [-2, -1, -3, -3, 2, -1, 0, 0, 2, 0, -2, 1, 0, -3, 1, -2]
// Dest PEs: [14, 15, 17, 18, 14, 15, 17, 18, 19, 20, 21, 22, 28, 29, 30, 31]
9'd8: rdata =    56'b00000000000000000000000000000000000000000000000000000011;
//
// shift amount: 1, Lanes IDs: [1, 2]
9'd9: rdata =    56'b00000000000000000000000000000000000000001101100001010001;
//
// shift amount: 2, Lanes IDs: [14, 15]
9'd10: rdata =   56'b00100100000000000000000000000000000000000000000001010010;
//
// shift amount: 5, Lanes IDs: [1, 2]
9'd11: rdata =   56'b00000000000000000000000000000000000000001101100001010101;
//
// shift amount: 6, Lanes IDs: [14, 15]
9'd12: rdata =   56'b00100100000000000000000000000000000000000000000001010110;
//
// read [True, True, True, False]
// ['x(22,)', 'x(23,)', 'x(25,)', 'x(26,)', 'x(102,)', 'x(103,)', 'x(105,)', 'x(106,)', 'x(184,)', 'x(185,)', 'x(187,)', 'x(188,)', 'x(276,)', 'x(277,)', 'x(279,)', 'x(280,)']
// Data values: [0, -3, 2, 1, -2, 2, -1, 2, 2, 0, -2, 1, 0, -3, 1, -2]
// Dest PEs: [19, 20, 21, 22, 19, 20, 21, 22, 19, 20, 21, 22, 28, 29, 30, 31]
9'd13: rdata =   56'b00000000000000000000000000000000000000000000000000000111;
//
// shift amount: 13, Lanes IDs: [3, 4, 5, 6]
9'd14: rdata =   56'b00000000000000000000000000001101101101100000000001011101;
//
// shift amount: 1, Lanes IDs: [3, 4, 5, 6]
9'd15: rdata =   56'b00000000000000000000000000001101101101100000000001010001;
//
// shift amount: 5, Lanes IDs: [3, 4, 5, 6]
9'd16: rdata =   56'b00000000000000000000000000001101101101100000000001010101;
//
// read [True, True, True, False]
// ['x(28,)', 'x(29,)', 'x(31,)', 'x(32,)', 'x(108,)', 'x(109,)', 'x(111,)', 'x(112,)', 'x(190,)', 'x(191,)', 'x(193,)', 'x(194,)', 'x(276,)', 'x(277,)', 'x(279,)', 'x(280,)']
// Data values: [-2, 2, 1, 2, -1, -2, 1, 2, 0, 2, -3, 0, 0, -3, 1, -2]
// Dest PEs: [23, 25, 26, 27, 23, 25, 26, 27, 23, 25, 26, 27, 28, 29, 30, 31]
9'd17: rdata =   56'b00000000000000000000000000000000000000000000000000000111;
//
// shift amount: 8, Lanes IDs: [9, 10, 11]
9'd18: rdata =   56'b00000000000001101101100000000000000000000000000001011000;
//
// shift amount: 9, Lanes IDs: [7]
9'd19: rdata =   56'b00000000000000000000000001100000000000000000000001011001;
//
// shift amount: 12, Lanes IDs: [9, 10, 11]
9'd20: rdata =   56'b00000000000001101101100000000000000000000000000001011100;
//
// shift amount: 0, Lanes IDs: [9, 10, 11]
9'd21: rdata =   56'b00000000000001101101100000000000000000000000000001010000;
//
// shift amount: 13, Lanes IDs: [7]
9'd22: rdata =   56'b00000000000000000000000001100000000000000000000001011101;
//
// shift amount: 1, Lanes IDs: [7]
9'd23: rdata =   56'b00000000000000000000000001100000000000000000000001010001;
//
// read [True, True, True, True]
// ['x(34,)', 'x(35,)', 'x(37,)', 'x(38,)', 'x(114,)', 'x(115,)', 'x(117,)', 'x(118,)', 'x(196,)', 'x(197,)', 'x(198,)', 'x(199,)', 'x(276,)', 'x(277,)', 'x(279,)', 'x(280,)']
// Data values: [2, -3, -3, 2, -2, -3, -3, -3, 2, 0, 1, 0, 0, -3, 1, -2]
// Dest PEs: [28, 29, 30, 31, 28, 29, 30, 31, 28, 29, 30, 31, 28, 29, 30, 31]
9'd24: rdata =   56'b00000000000000000000000000000000000000000000000000001111;
//
// shift amount: 4, Lanes IDs: [12, 13, 14, 15]
9'd25: rdata =   56'b01101101101100000000000000000000000000000000000001010100;
//
// shift amount: 8, Lanes IDs: [12, 13, 14, 15]
9'd26: rdata =   56'b01101101101100000000000000000000000000000000000001011000;
//
// shift amount: 12, Lanes IDs: [12, 13, 14, 15]
9'd27: rdata =   56'b01101101101100000000000000000000000000000000000001011100;
//
// shift amount: 0, Lanes IDs: [12, 13, 14, 15]
9'd28: rdata =   56'b01101101101100000000000000000000000000000000000001010000;
//
// read [True, True, True, True]
// ['x(40,)', 'x(41,)', 'x(43,)', 'x(44,)', 'x(120,)', 'x(121,)', 'x(123,)', 'x(124,)', 'x(200,)', 'x(201,)', 'x(203,)', 'x(204,)', 'x(282,)', 'x(283,)', 'x(285,)', 'x(286,)']
// Data values: [-1, -2, 2, -2, -1, -3, -1, -2, 0, -1, -3, -2, 2, 0, -2, 2]
// Dest PEs: [33, 34, 35, 36, 33, 34, 35, 36, 33, 34, 35, 36, 33, 34, 35, 36]
9'd29: rdata =   56'b00000000000000000000000000000000000000000000000000001111;
//
// shift amount: 15, Lanes IDs: [1, 2, 3, 4]
9'd30: rdata =   56'b00000000000000000000000000000000010110110110100001011111;
//
// shift amount: 3, Lanes IDs: [1, 2, 3, 4]
9'd31: rdata =   56'b00000000000000000000000000000000010110110110100001010011;
//
// shift amount: 7, Lanes IDs: [1, 2, 3, 4]
9'd32: rdata =   56'b00000000000000000000000000000000010110110110100001010111;
//
// shift amount: 11, Lanes IDs: [1, 2, 3, 4]
9'd33: rdata =   56'b00000000000000000000000000000000010110110110100001011011;
//
// read [True, True, True, True]
// ['x(46,)', 'x(47,)', 'x(49,)', 'x(50,)', 'x(126,)', 'x(127,)', 'x(129,)', 'x(130,)', 'x(206,)', 'x(207,)', 'x(209,)', 'x(210,)', 'x(288,)', 'x(289,)', 'x(291,)', 'x(292,)']
// Data values: [-2, 0, -3, 0, 1, -2, -2, -3, 1, -3, -1, 1, -1, 1, 1, 1]
// Dest PEs: [37, 38, 39, 41, 37, 38, 39, 41, 37, 38, 39, 41, 37, 38, 39, 41]
9'd34: rdata =   56'b00000000000000000000000000000000000000000000000000001111;
//
// shift amount: 10, Lanes IDs: [9]
9'd35: rdata =   56'b00000000000000000010100000000000000000000000000001011010;
//
// shift amount: 11, Lanes IDs: [5, 6, 7]
9'd36: rdata =   56'b00000000000000000000000010110110100000000000000001011011;
//
// shift amount: 14, Lanes IDs: [9]
9'd37: rdata =   56'b00000000000000000010100000000000000000000000000001011110;
//
// shift amount: 2, Lanes IDs: [9]
9'd38: rdata =   56'b00000000000000000010100000000000000000000000000001010010;
//
// shift amount: 6, Lanes IDs: [9]
9'd39: rdata =   56'b00000000000000000010100000000000000000000000000001010110;
//
// shift amount: 15, Lanes IDs: [5, 6, 7]
9'd40: rdata =   56'b00000000000000000000000010110110100000000000000001011111;
//
// shift amount: 3, Lanes IDs: [5, 6, 7]
9'd41: rdata =   56'b00000000000000000000000010110110100000000000000001010011;
//
// shift amount: 7, Lanes IDs: [5, 6, 7]
9'd42: rdata =   56'b00000000000000000000000010110110100000000000000001010111;
//
// read [True, True, True, True]
// ['x(51,)', 'x(52,)', 'x(53,)', 'x(54,)', 'x(132,)', 'x(133,)', 'x(135,)', 'x(136,)', 'x(212,)', 'x(213,)', 'x(215,)', 'x(216,)', 'x(294,)', 'x(295,)', 'x(296,)', 'x(297,)']
// Data values: [2, -2, 0, -3, -3, 2, 0, 0, 1, 1, -1, 2, -3, 1, 0, 0]
// Dest PEs: [42, 43, 44, 45, 42, 43, 44, 45, 42, 43, 44, 45, 42, 43, 44, 45]
9'd43: rdata =   56'b00000000000000000000000000000000000000000000000000001111;
//
// shift amount: 6, Lanes IDs: [10, 11, 12, 13]
9'd44: rdata =   56'b00000010110110110100000000000000000000000000000001010110;
//
// shift amount: 10, Lanes IDs: [10, 11, 12, 13]
9'd45: rdata =   56'b00000010110110110100000000000000000000000000000001011010;
//
// shift amount: 14, Lanes IDs: [10, 11, 12, 13]
9'd46: rdata =   56'b00000010110110110100000000000000000000000000000001011110;
//
// shift amount: 2, Lanes IDs: [10, 11, 12, 13]
9'd47: rdata =   56'b00000010110110110100000000000000000000000000000001010010;
//
// read [True, True, True, True]
// ['x(56,)', 'x(57,)', 'x(59,)', 'x(60,)', 'x(138,)', 'x(139,)', 'x(141,)', 'x(142,)', 'x(218,)', 'x(219,)', 'x(221,)', 'x(222,)', 'x(298,)', 'x(299,)', 'x(301,)', 'x(302,)']
// Data values: [-2, -2, 0, 2, 1, -3, -3, -2, -1, 0, -2, -2, -1, -1, 1, 0]
// Dest PEs: [46, 47, 49, 50, 46, 47, 49, 50, 46, 47, 49, 50, 46, 47, 49, 50]
9'd48: rdata =   56'b00000000000000000000000000000000000000000000000000001111;
//
// shift amount: 1, Lanes IDs: [1, 2]
9'd49: rdata =   56'b00000000000000000000000000000000000000011111100001010001;
//
// shift amount: 2, Lanes IDs: [14, 15]
9'd50: rdata =   56'b10110100000000000000000000000000000000000000000001010010;
//
// shift amount: 5, Lanes IDs: [1, 2]
9'd51: rdata =   56'b00000000000000000000000000000000000000011111100001010101;
//
// shift amount: 6, Lanes IDs: [14, 15]
9'd52: rdata =   56'b10110100000000000000000000000000000000000000000001010110;
//
// shift amount: 9, Lanes IDs: [1, 2]
9'd53: rdata =   56'b00000000000000000000000000000000000000011111100001011001;
//
// shift amount: 10, Lanes IDs: [14, 15]
9'd54: rdata =   56'b10110100000000000000000000000000000000000000000001011010;
//
// shift amount: 13, Lanes IDs: [1, 2]
9'd55: rdata =   56'b00000000000000000000000000000000000000011111100001011101;
//
// shift amount: 14, Lanes IDs: [14, 15]
9'd56: rdata =   56'b10110100000000000000000000000000000000000000000001011110;
//
// read [True, True, True, True]
// ['x(62,)', 'x(63,)', 'x(65,)', 'x(66,)', 'x(144,)', 'x(145,)', 'x(147,)', 'x(148,)', 'x(224,)', 'x(225,)', 'x(227,)', 'x(228,)', 'x(304,)', 'x(305,)', 'x(307,)', 'x(308,)']
// Data values: [1, 1, 1, -1, -3, 2, -2, -1, 2, 1, 2, 0, 0, 1, 1, -1]
// Dest PEs: [51, 52, 53, 54, 51, 52, 53, 54, 51, 52, 53, 54, 51, 52, 53, 54]
9'd57: rdata =   56'b00000000000000000000000000000000000000000000000000001111;
//
// shift amount: 13, Lanes IDs: [3, 4, 5, 6]
9'd58: rdata =   56'b00000000000000000000000000011111111111100000000001011101;
//
// shift amount: 1, Lanes IDs: [3, 4, 5, 6]
9'd59: rdata =   56'b00000000000000000000000000011111111111100000000001010001;
//
// shift amount: 5, Lanes IDs: [3, 4, 5, 6]
9'd60: rdata =   56'b00000000000000000000000000011111111111100000000001010101;
//
// shift amount: 9, Lanes IDs: [3, 4, 5, 6]
9'd61: rdata =   56'b00000000000000000000000000011111111111100000000001011001;
//
// read [True, True, True, True]
// ['x(68,)', 'x(69,)', 'x(71,)', 'x(72,)', 'x(149,)', 'x(150,)', 'x(151,)', 'x(152,)', 'x(230,)', 'x(231,)', 'x(233,)', 'x(234,)', 'x(310,)', 'x(311,)', 'x(313,)', 'x(314,)']
// Data values: [2, 1, -1, 2, 2, 0, -2, -2, -2, -2, 2, 2, 1, 1, -3, -2]
// Dest PEs: [55, 57, 58, 59, 55, 57, 58, 59, 55, 57, 58, 59, 55, 57, 58, 59]
9'd62: rdata =   56'b00000000000000000000000000000000000000000000000000001111;
//
// shift amount: 8, Lanes IDs: [9, 10, 11]
9'd63: rdata =   56'b00000000000011111111100000000000000000000000000001011000;
//
// shift amount: 9, Lanes IDs: [7]
9'd64: rdata =   56'b00000000000000000000000011100000000000000000000001011001;
//
// shift amount: 12, Lanes IDs: [9, 10, 11]
9'd65: rdata =   56'b00000000000011111111100000000000000000000000000001011100;
//
// shift amount: 0, Lanes IDs: [9, 10, 11]
9'd66: rdata =   56'b00000000000011111111100000000000000000000000000001010000;
//
// shift amount: 4, Lanes IDs: [9, 10, 11]
9'd67: rdata =   56'b00000000000011111111100000000000000000000000000001010100;
//
// shift amount: 13, Lanes IDs: [7]
9'd68: rdata =   56'b00000000000000000000000011100000000000000000000001011101;
//
// shift amount: 1, Lanes IDs: [7]
9'd69: rdata =   56'b00000000000000000000000011100000000000000000000001010001;
//
// shift amount: 5, Lanes IDs: [7]
9'd70: rdata =   56'b00000000000000000000000011100000000000000000000001010101;
//
// read [True, True, True, True]
// ['x(74,)', 'x(75,)', 'x(77,)', 'x(78,)', 'x(154,)', 'x(155,)', 'x(157,)', 'x(158,)', 'x(236,)', 'x(237,)', 'x(239,)', 'x(240,)', 'x(316,)', 'x(317,)', 'x(319,)', 'x(320,)']
// Data values: [-2, -3, -3, -1, 2, -2, -1, -2, -3, -3, -3, 1, -3, 2, 2, -3]
// Dest PEs: [60, 61, 62, 63, 60, 61, 62, 63, 60, 61, 62, 63, 60, 61, 62, 63]
9'd71: rdata =   56'b00000000000000000000000000000000000000000000000000001111;
//
// shift amount: 4, Lanes IDs: [12, 13, 14, 15]
9'd72: rdata =   56'b11111111111100000000000000000000000000000000000001010100;
//
// shift amount: 8, Lanes IDs: [12, 13, 14, 15]
9'd73: rdata =   56'b11111111111100000000000000000000000000000000000001011000;
//
// shift amount: 12, Lanes IDs: [12, 13, 14, 15]
9'd74: rdata =   56'b11111111111100000000000000000000000000000000000001011100;
//
// shift amount: 0, Lanes IDs: [12, 13, 14, 15]
9'd75: rdata =   56'b11111111111100000000000000000000000000000000000001010000;
//
// read [True, True, True, True]
// ['x(80,)', 'x(81,)', 'x(83,)', 'x(84,)', 'x(160,)', 'x(161,)', 'x(163,)', 'x(164,)', 'x(242,)', 'x(243,)', 'x(245,)', 'x(246,)', 'x(322,)', 'x(323,)', 'x(325,)', 'x(326,)']
// Data values: [-3, 2, 1, -1, -2, -1, 1, 0, -3, 0, 1, -3, -2, 1, 2, 1]
// Dest PEs: [1, 2, 3, 4, 1, 2, 3, 4, 1, 2, 3, 4, 1, 2, 3, 4]
9'd76: rdata =   56'b00000000000000000000000000000000000000000000000000001111;
//
// shift amount: 15, Lanes IDs: [1, 2, 3, 4]
9'd77: rdata =   56'b00000000000000000000000000000000000100100100100001011111;
//
// shift amount: 3, Lanes IDs: [1, 2, 3, 4]
9'd78: rdata =   56'b00000000000000000000000000000000000100100100100001010011;
//
// shift amount: 7, Lanes IDs: [1, 2, 3, 4]
9'd79: rdata =   56'b00000000000000000000000000000000000100100100100001010111;
//
// shift amount: 11, Lanes IDs: [1, 2, 3, 4]
9'd80: rdata =   56'b00000000000000000000000000000000000100100100100001011011;
//
// read [True, True, True, True]
// ['x(86,)', 'x(87,)', 'x(89,)', 'x(90,)', 'x(166,)', 'x(167,)', 'x(169,)', 'x(170,)', 'x(247,)', 'x(248,)', 'x(249,)', 'x(250,)', 'x(328,)', 'x(329,)', 'x(331,)', 'x(332,)']
// Data values: [-2, 0, 1, -3, -1, 0, -3, -1, 1, 0, 0, -1, 2, 2, 2, 1]
// Dest PEs: [5, 6, 7, 9, 5, 6, 7, 9, 5, 6, 7, 9, 5, 6, 7, 9]
9'd81: rdata =   56'b00000000000000000000000000000000000000000000000000001111;
//
// shift amount: 10, Lanes IDs: [9]
9'd82: rdata =   56'b00000000000000000000100000000000000000000000000001011010;
//
// shift amount: 11, Lanes IDs: [5, 6, 7]
9'd83: rdata =   56'b00000000000000000000000000100100100000000000000001011011;
//
// shift amount: 14, Lanes IDs: [9]
9'd84: rdata =   56'b00000000000000000000100000000000000000000000000001011110;
//
// shift amount: 2, Lanes IDs: [9]
9'd85: rdata =   56'b00000000000000000000100000000000000000000000000001010010;
//
// shift amount: 6, Lanes IDs: [9]
9'd86: rdata =   56'b00000000000000000000100000000000000000000000000001010110;
//
// shift amount: 15, Lanes IDs: [5, 6, 7]
9'd87: rdata =   56'b00000000000000000000000000100100100000000000000001011111;
//
// shift amount: 3, Lanes IDs: [5, 6, 7]
9'd88: rdata =   56'b00000000000000000000000000100100100000000000000001010011;
//
// shift amount: 7, Lanes IDs: [5, 6, 7]
9'd89: rdata =   56'b00000000000000000000000000100100100000000000000001010111;
//
// read [True, True, True, True]
// ['x(368,)', 'x(369,)', 'x(371,)', 'x(372,)', 'x(172,)', 'x(173,)', 'x(175,)', 'x(176,)', 'x(252,)', 'x(253,)', 'x(255,)', 'x(256,)', 'x(334,)', 'x(335,)', 'x(337,)', 'x(338,)']
// Data values: [0, -1, -2, -2, -1, 1, 1, 1, -1, -1, 0, -3, -2, -3, -2, -3]
// Dest PEs: [37, 38, 39, 41, 10, 11, 12, 13, 10, 11, 12, 13, 10, 11, 12, 13]
9'd90: rdata =   56'b00000000000000000000000000000000000000000000000000001111;
//
// shift amount: 10, Lanes IDs: [9, 10, 11, 12, 13]
9'd91: rdata =   56'b00000000100100100110100000000000000000000000000001011010;
//
// shift amount: 11, Lanes IDs: [5, 6, 7]
9'd92: rdata =   56'b00000000000000000000000010110110100000000000000001011011;
//
// shift amount: 14, Lanes IDs: [10, 11, 12, 13]
9'd93: rdata =   56'b00000000100100100100000000000000000000000000000001011110;
//
// shift amount: 2, Lanes IDs: [10, 11, 12, 13]
9'd94: rdata =   56'b00000000100100100100000000000000000000000000000001010010;
//
// read [True, True, True, True]
// ['x(374,)', 'x(375,)', 'x(377,)', 'x(378,)', 'x(178,)', 'x(179,)', 'x(181,)', 'x(182,)', 'x(258,)', 'x(259,)', 'x(261,)', 'x(262,)', 'x(340,)', 'x(341,)', 'x(343,)', 'x(344,)']
// Data values: [1, 2, -3, -2, -3, 1, 0, -2, 1, -3, 0, 1, -2, 2, 1, 0]
// Dest PEs: [42, 43, 44, 45, 14, 15, 17, 18, 14, 15, 17, 18, 14, 15, 17, 18]
9'd95: rdata =   56'b00000000000000000000000000000000000000000000000000001111;
//
// shift amount: 5, Lanes IDs: [1, 2]
9'd96: rdata =   56'b00000000000000000000000000000000000000001101100001010101;
//
// shift amount: 6, Lanes IDs: [10, 11, 12, 13, 14, 15]
9'd97: rdata =   56'b00100110110110110100000000000000000000000000000001010110;
//
// shift amount: 9, Lanes IDs: [1, 2]
9'd98: rdata =   56'b00000000000000000000000000000000000000001101100001011001;
//
// shift amount: 10, Lanes IDs: [14, 15]
9'd99: rdata =   56'b00100100000000000000000000000000000000000000000001011010;
//
// shift amount: 13, Lanes IDs: [1, 2]
9'd100: rdata =  56'b00000000000000000000000000000000000000001101100001011101;
//
// shift amount: 14, Lanes IDs: [14, 15]
9'd101: rdata =  56'b00100100000000000000000000000000000000000000000001011110;
//
// read [True, True, True, True]
// ['x(380,)', 'x(381,)', 'x(383,)', 'x(384,)', 'x(460,)', 'x(461,)', 'x(463,)', 'x(464,)', 'x(264,)', 'x(265,)', 'x(267,)', 'x(268,)', 'x(345,)', 'x(346,)', 'x(347,)', 'x(348,)']
// Data values: [-3, -3, 2, -2, -3, 1, 0, 1, -1, -1, -1, 1, -1, 2, -3, -3]
// Dest PEs: [46, 47, 49, 50, 46, 47, 49, 50, 19, 20, 21, 22, 19, 20, 21, 22]
9'd102: rdata =  56'b00000000000000000000000000000000000000000000000000001111;
//
// shift amount: 1, Lanes IDs: [1, 2]
9'd103: rdata =  56'b00000000000000000000000000000000000000011111100001010001;
//
// shift amount: 2, Lanes IDs: [14, 15]
9'd104: rdata =  56'b10110100000000000000000000000000000000000000000001010010;
//
// shift amount: 5, Lanes IDs: [1, 2, 3, 4, 5, 6]
9'd105: rdata =  56'b00000000000000000000000000001101101101111111100001010101;
//
// shift amount: 6, Lanes IDs: [14, 15]
9'd106: rdata =  56'b10110100000000000000000000000000000000000000000001010110;
//
// shift amount: 9, Lanes IDs: [3, 4, 5, 6]
9'd107: rdata =  56'b00000000000000000000000000001101101101100000000001011001;
//
// read [True, True, True, True]
// ['x(386,)', 'x(387,)', 'x(389,)', 'x(390,)', 'x(466,)', 'x(467,)', 'x(469,)', 'x(470,)', 'x(270,)', 'x(271,)', 'x(273,)', 'x(274,)', 'x(350,)', 'x(351,)', 'x(353,)', 'x(354,)']
// Data values: [0, -3, -3, 0, -3, -2, -2, -3, 1, -3, 0, -1, -3, -2, -1, 2]
// Dest PEs: [51, 52, 53, 54, 51, 52, 53, 54, 23, 25, 26, 27, 23, 25, 26, 27]
9'd108: rdata =  56'b00000000000000000000000000000000000000000000000000001111;
//
// shift amount: 0, Lanes IDs: [9, 10, 11]
9'd109: rdata =  56'b00000000000001101101100000000000000000000000000001010000;
//
// shift amount: 4, Lanes IDs: [9, 10, 11]
9'd110: rdata =  56'b00000000000001101101100000000000000000000000000001010100;
//
// shift amount: 13, Lanes IDs: [3, 4, 5, 6]
9'd111: rdata =  56'b00000000000000000000000000011111111111100000000001011101;
//
// shift amount: 1, Lanes IDs: [3, 4, 5, 6, 7]
9'd112: rdata =  56'b00000000000000000000000001111111111111100000000001010001;
//
// shift amount: 5, Lanes IDs: [7]
9'd113: rdata =  56'b00000000000000000000000001100000000000000000000001010101;
//
// read [True, True, True, True]
// ['x(392,)', 'x(393,)', 'x(394,)', 'x(395,)', 'x(472,)', 'x(473,)', 'x(475,)', 'x(476,)', 'x(552,)', 'x(553,)', 'x(555,)', 'x(556,)', 'x(356,)', 'x(357,)', 'x(359,)', 'x(360,)']
// Data values: [-3, -2, 0, 0, -1, -2, 1, 0, 2, -2, -2, -3, -1, -3, 2, 2]
// Dest PEs: [55, 57, 58, 59, 55, 57, 58, 59, 55, 57, 58, 59, 28, 29, 30, 31]
9'd114: rdata =  56'b00000000000000000000000000000000000000000000000000001111;
//
// shift amount: 8, Lanes IDs: [9, 10, 11]
9'd115: rdata =  56'b00000000000011111111100000000000000000000000000001011000;
//
// shift amount: 9, Lanes IDs: [7]
9'd116: rdata =  56'b00000000000000000000000011100000000000000000000001011001;
//
// shift amount: 12, Lanes IDs: [9, 10, 11]
9'd117: rdata =  56'b00000000000011111111100000000000000000000000000001011100;
//
// shift amount: 0, Lanes IDs: [9, 10, 11, 12, 13, 14, 15]
9'd118: rdata =  56'b01101101101111111111100000000000000000000000000001010000;
//
// shift amount: 13, Lanes IDs: [7]
9'd119: rdata =  56'b00000000000000000000000011100000000000000000000001011101;
//
// shift amount: 1, Lanes IDs: [7]
9'd120: rdata =  56'b00000000000000000000000011100000000000000000000001010001;
//
// read [True, True, True, True]
// ['x(396,)', 'x(397,)', 'x(399,)', 'x(400,)', 'x(478,)', 'x(479,)', 'x(481,)', 'x(482,)', 'x(558,)', 'x(559,)', 'x(561,)', 'x(562,)', 'x(362,)', 'x(363,)', 'x(365,)', 'x(366,)']
// Data values: [2, 1, 2, -3, 2, 0, -3, 0, 1, 1, -2, 1, -2, 1, -1, 1]
// Dest PEs: [60, 61, 62, 63, 60, 61, 62, 63, 60, 61, 62, 63, 33, 34, 35, 36]
9'd121: rdata =  56'b00000000000000000000000000000000000000000000000000001111;
//
// shift amount: 11, Lanes IDs: [1, 2, 3, 4]
9'd122: rdata =  56'b00000000000000000000000000000000010110110110100001011011;
//
// shift amount: 4, Lanes IDs: [12, 13, 14, 15]
9'd123: rdata =  56'b11111111111100000000000000000000000000000000000001010100;
//
// shift amount: 8, Lanes IDs: [12, 13, 14, 15]
9'd124: rdata =  56'b11111111111100000000000000000000000000000000000001011000;
//
// shift amount: 12, Lanes IDs: [12, 13, 14, 15]
9'd125: rdata =  56'b11111111111100000000000000000000000000000000000001011100;
//
// read [True, True, True, True]
// ['x(402,)', 'x(403,)', 'x(405,)', 'x(406,)', 'x(484,)', 'x(485,)', 'x(487,)', 'x(488,)', 'x(564,)', 'x(565,)', 'x(567,)', 'x(568,)', 'x(644,)', 'x(645,)', 'x(647,)', 'x(648,)']
// Data values: [-2, 1, 0, 1, -1, 1, -3, -1, 1, 0, -2, 2, 2, -1, 1, -3]
// Dest PEs: [1, 2, 3, 4, 1, 2, 3, 4, 1, 2, 3, 4, 1, 2, 3, 4]
9'd126: rdata =  56'b00000000000000000000000000000000000000000000000000001111;
//
// shift amount: 15, Lanes IDs: [1, 2, 3, 4]
9'd127: rdata =  56'b00000000000000000000000000000000000100100100100001011111;
//
// shift amount: 3, Lanes IDs: [1, 2, 3, 4]
9'd128: rdata =  56'b00000000000000000000000000000000000100100100100001010011;
//
// shift amount: 7, Lanes IDs: [1, 2, 3, 4]
9'd129: rdata =  56'b00000000000000000000000000000000000100100100100001010111;
//
// shift amount: 11, Lanes IDs: [1, 2, 3, 4]
9'd130: rdata =  56'b00000000000000000000000000000000000100100100100001011011;
//
// read [True, True, True, True]
// ['x(408,)', 'x(409,)', 'x(411,)', 'x(412,)', 'x(490,)', 'x(491,)', 'x(492,)', 'x(493,)', 'x(570,)', 'x(571,)', 'x(573,)', 'x(574,)', 'x(650,)', 'x(651,)', 'x(653,)', 'x(654,)']
// Data values: [-3, -1, 1, -1, 0, -3, -1, 0, -2, 2, -2, 1, 1, 1, 0, 1]
// Dest PEs: [5, 6, 7, 9, 5, 6, 7, 9, 5, 6, 7, 9, 5, 6, 7, 9]
9'd131: rdata =  56'b00000000000000000000000000000000000000000000000000001111;
//
// shift amount: 10, Lanes IDs: [9]
9'd132: rdata =  56'b00000000000000000000100000000000000000000000000001011010;
//
// shift amount: 11, Lanes IDs: [5, 6, 7]
9'd133: rdata =  56'b00000000000000000000000000100100100000000000000001011011;
//
// shift amount: 14, Lanes IDs: [9]
9'd134: rdata =  56'b00000000000000000000100000000000000000000000000001011110;
//
// shift amount: 2, Lanes IDs: [9]
9'd135: rdata =  56'b00000000000000000000100000000000000000000000000001010010;
//
// shift amount: 6, Lanes IDs: [9]
9'd136: rdata =  56'b00000000000000000000100000000000000000000000000001010110;
//
// shift amount: 15, Lanes IDs: [5, 6, 7]
9'd137: rdata =  56'b00000000000000000000000000100100100000000000000001011111;
//
// shift amount: 3, Lanes IDs: [5, 6, 7]
9'd138: rdata =  56'b00000000000000000000000000100100100000000000000001010011;
//
// shift amount: 7, Lanes IDs: [5, 6, 7]
9'd139: rdata =  56'b00000000000000000000000000100100100000000000000001010111;
//
// read [True, True, True, True]
// ['x(414,)', 'x(415,)', 'x(417,)', 'x(418,)', 'x(494,)', 'x(495,)', 'x(497,)', 'x(498,)', 'x(576,)', 'x(577,)', 'x(579,)', 'x(580,)', 'x(656,)', 'x(657,)', 'x(659,)', 'x(660,)']
// Data values: [-2, -2, -1, 1, 1, 0, 2, -1, -2, 1, 0, 2, -3, -3, 2, 1]
// Dest PEs: [10, 11, 12, 13, 10, 11, 12, 13, 10, 11, 12, 13, 10, 11, 12, 13]
9'd140: rdata =  56'b00000000000000000000000000000000000000000000000000001111;
//
// shift amount: 6, Lanes IDs: [10, 11, 12, 13]
9'd141: rdata =  56'b00000000100100100100000000000000000000000000000001010110;
//
// shift amount: 10, Lanes IDs: [10, 11, 12, 13]
9'd142: rdata =  56'b00000000100100100100000000000000000000000000000001011010;
//
// shift amount: 14, Lanes IDs: [10, 11, 12, 13]
9'd143: rdata =  56'b00000000100100100100000000000000000000000000000001011110;
//
// shift amount: 2, Lanes IDs: [10, 11, 12, 13]
9'd144: rdata =  56'b00000000100100100100000000000000000000000000000001010010;
//
// read [True, True, True, True]
// ['x(420,)', 'x(421,)', 'x(423,)', 'x(424,)', 'x(500,)', 'x(501,)', 'x(503,)', 'x(504,)', 'x(582,)', 'x(583,)', 'x(585,)', 'x(586,)', 'x(662,)', 'x(663,)', 'x(665,)', 'x(666,)']
// Data values: [0, -3, -3, -3, 1, -2, -3, -1, 1, -2, 1, 1, -1, -2, 1, 2]
// Dest PEs: [14, 15, 17, 18, 14, 15, 17, 18, 14, 15, 17, 18, 14, 15, 17, 18]
9'd145: rdata =  56'b00000000000000000000000000000000000000000000000000001111;
//
// shift amount: 1, Lanes IDs: [1, 2]
9'd146: rdata =  56'b00000000000000000000000000000000000000001101100001010001;
//
// shift amount: 2, Lanes IDs: [14, 15]
9'd147: rdata =  56'b00100100000000000000000000000000000000000000000001010010;
//
// shift amount: 5, Lanes IDs: [1, 2]
9'd148: rdata =  56'b00000000000000000000000000000000000000001101100001010101;
//
// shift amount: 6, Lanes IDs: [14, 15]
9'd149: rdata =  56'b00100100000000000000000000000000000000000000000001010110;
//
// shift amount: 9, Lanes IDs: [1, 2]
9'd150: rdata =  56'b00000000000000000000000000000000000000001101100001011001;
//
// shift amount: 10, Lanes IDs: [14, 15]
9'd151: rdata =  56'b00100100000000000000000000000000000000000000000001011010;
//
// shift amount: 13, Lanes IDs: [1, 2]
9'd152: rdata =  56'b00000000000000000000000000000000000000001101100001011101;
//
// shift amount: 14, Lanes IDs: [14, 15]
9'd153: rdata =  56'b00100100000000000000000000000000000000000000000001011110;
//
// read [True, True, True, True]
// ['x(426,)', 'x(427,)', 'x(429,)', 'x(430,)', 'x(506,)', 'x(507,)', 'x(509,)', 'x(510,)', 'x(588,)', 'x(589,)', 'x(590,)', 'x(591,)', 'x(668,)', 'x(669,)', 'x(671,)', 'x(672,)']
// Data values: [-2, -3, -2, 2, 1, 0, 2, 2, 0, 2, -3, 2, 2, 1, 2, -3]
// Dest PEs: [19, 20, 21, 22, 19, 20, 21, 22, 19, 20, 21, 22, 19, 20, 21, 22]
9'd154: rdata =  56'b00000000000000000000000000000000000000000000000000001111;
//
// shift amount: 13, Lanes IDs: [3, 4, 5, 6]
9'd155: rdata =  56'b00000000000000000000000000001101101101100000000001011101;
//
// shift amount: 1, Lanes IDs: [3, 4, 5, 6]
9'd156: rdata =  56'b00000000000000000000000000001101101101100000000001010001;
//
// shift amount: 5, Lanes IDs: [3, 4, 5, 6]
9'd157: rdata =  56'b00000000000000000000000000001101101101100000000001010101;
//
// shift amount: 9, Lanes IDs: [3, 4, 5, 6]
9'd158: rdata =  56'b00000000000000000000000000001101101101100000000001011001;
//
// read [True, True, True, True]
// ['x(432,)', 'x(433,)', 'x(435,)', 'x(436,)', 'x(512,)', 'x(513,)', 'x(515,)', 'x(516,)', 'x(592,)', 'x(593,)', 'x(595,)', 'x(596,)', 'x(674,)', 'x(675,)', 'x(677,)', 'x(678,)']
// Data values: [-1, -3, 2, -3, 0, -1, 2, -1, -1, 0, 0, 2, 1, 1, 2, 0]
// Dest PEs: [23, 25, 26, 27, 23, 25, 26, 27, 23, 25, 26, 27, 23, 25, 26, 27]
9'd159: rdata =  56'b00000000000000000000000000000000000000000000000000001111;
//
// shift amount: 8, Lanes IDs: [9, 10, 11]
9'd160: rdata =  56'b00000000000001101101100000000000000000000000000001011000;
//
// shift amount: 9, Lanes IDs: [7]
9'd161: rdata =  56'b00000000000000000000000001100000000000000000000001011001;
//
// shift amount: 12, Lanes IDs: [9, 10, 11]
9'd162: rdata =  56'b00000000000001101101100000000000000000000000000001011100;
//
// shift amount: 0, Lanes IDs: [9, 10, 11]
9'd163: rdata =  56'b00000000000001101101100000000000000000000000000001010000;
//
// shift amount: 4, Lanes IDs: [9, 10, 11]
9'd164: rdata =  56'b00000000000001101101100000000000000000000000000001010100;
//
// shift amount: 13, Lanes IDs: [7]
9'd165: rdata =  56'b00000000000000000000000001100000000000000000000001011101;
//
// shift amount: 1, Lanes IDs: [7]
9'd166: rdata =  56'b00000000000000000000000001100000000000000000000001010001;
//
// shift amount: 5, Lanes IDs: [7]
9'd167: rdata =  56'b00000000000000000000000001100000000000000000000001010101;
//
// read [True, True, True, True]
// ['x(438,)', 'x(439,)', 'x(441,)', 'x(442,)', 'x(518,)', 'x(519,)', 'x(521,)', 'x(522,)', 'x(598,)', 'x(599,)', 'x(601,)', 'x(602,)', 'x(680,)', 'x(681,)', 'x(683,)', 'x(684,)']
// Data values: [2, 2, 0, 2, 0, -1, 2, -1, 2, 0, -3, -3, -1, 2, 1, -1]
// Dest PEs: [28, 29, 30, 31, 28, 29, 30, 31, 28, 29, 30, 31, 28, 29, 30, 31]
9'd168: rdata =  56'b00000000000000000000000000000000000000000000000000001111;
//
// shift amount: 4, Lanes IDs: [12, 13, 14, 15]
9'd169: rdata =  56'b01101101101100000000000000000000000000000000000001010100;
//
// shift amount: 8, Lanes IDs: [12, 13, 14, 15]
9'd170: rdata =  56'b01101101101100000000000000000000000000000000000001011000;
//
// shift amount: 12, Lanes IDs: [12, 13, 14, 15]
9'd171: rdata =  56'b01101101101100000000000000000000000000000000000001011100;
//
// shift amount: 0, Lanes IDs: [12, 13, 14, 15]
9'd172: rdata =  56'b01101101101100000000000000000000000000000000000001010000;
//
// read [True, True, True, True]
// ['x(443,)', 'x(444,)', 'x(445,)', 'x(446,)', 'x(524,)', 'x(525,)', 'x(527,)', 'x(528,)', 'x(604,)', 'x(605,)', 'x(607,)', 'x(608,)', 'x(686,)', 'x(687,)', 'x(688,)', 'x(689,)']
// Data values: [1, 0, -1, 0, -2, 0, -3, -3, 0, -1, 1, -2, 0, 1, 2, 1]
// Dest PEs: [33, 34, 35, 36, 33, 34, 35, 36, 33, 34, 35, 36, 33, 34, 35, 36]
9'd173: rdata =  56'b00000000000000000000000000000000000000000000000000001111;
//
// shift amount: 15, Lanes IDs: [1, 2, 3, 4]
9'd174: rdata =  56'b00000000000000000000000000000000010110110110100001011111;
//
// shift amount: 3, Lanes IDs: [1, 2, 3, 4]
9'd175: rdata =  56'b00000000000000000000000000000000010110110110100001010011;
//
// shift amount: 7, Lanes IDs: [1, 2, 3, 4]
9'd176: rdata =  56'b00000000000000000000000000000000010110110110100001010111;
//
// shift amount: 11, Lanes IDs: [1, 2, 3, 4]
9'd177: rdata =  56'b00000000000000000000000000000000010110110110100001011011;
//
// read [True, True, True, True]
// ['x(448,)', 'x(449,)', 'x(451,)', 'x(452,)', 'x(530,)', 'x(531,)', 'x(533,)', 'x(534,)', 'x(610,)', 'x(611,)', 'x(613,)', 'x(614,)', 'x(690,)', 'x(691,)', 'x(693,)', 'x(694,)']
// Data values: [-2, 0, 2, 0, 1, 2, -3, -3, -1, 1, -1, 1, 2, 1, -3, 2]
// Dest PEs: [37, 38, 39, 41, 37, 38, 39, 41, 37, 38, 39, 41, 37, 38, 39, 41]
9'd178: rdata =  56'b00000000000000000000000000000000000000000000000000001111;
//
// shift amount: 10, Lanes IDs: [9]
9'd179: rdata =  56'b00000000000000000010100000000000000000000000000001011010;
//
// shift amount: 11, Lanes IDs: [5, 6, 7]
9'd180: rdata =  56'b00000000000000000000000010110110100000000000000001011011;
//
// shift amount: 14, Lanes IDs: [9]
9'd181: rdata =  56'b00000000000000000010100000000000000000000000000001011110;
//
// shift amount: 2, Lanes IDs: [9]
9'd182: rdata =  56'b00000000000000000010100000000000000000000000000001010010;
//
// shift amount: 6, Lanes IDs: [9]
9'd183: rdata =  56'b00000000000000000010100000000000000000000000000001010110;
//
// shift amount: 15, Lanes IDs: [5, 6, 7]
9'd184: rdata =  56'b00000000000000000000000010110110100000000000000001011111;
//
// shift amount: 3, Lanes IDs: [5, 6, 7]
9'd185: rdata =  56'b00000000000000000000000010110110100000000000000001010011;
//
// shift amount: 7, Lanes IDs: [5, 6, 7]
9'd186: rdata =  56'b00000000000000000000000010110110100000000000000001010111;
//
// read [True, True, True, True]
// ['x(454,)', 'x(455,)', 'x(457,)', 'x(458,)', 'x(536,)', 'x(537,)', 'x(539,)', 'x(540,)', 'x(616,)', 'x(617,)', 'x(619,)', 'x(620,)', 'x(696,)', 'x(697,)', 'x(699,)', 'x(700,)']
// Data values: [-3, 2, 1, -1, -2, -2, -3, 1, -1, -1, 1, 2, -3, -3, -2, -1]
// Dest PEs: [42, 43, 44, 45, 42, 43, 44, 45, 42, 43, 44, 45, 42, 43, 44, 45]
9'd187: rdata =  56'b00000000000000000000000000000000000000000000000000001111;
//
// shift amount: 6, Lanes IDs: [10, 11, 12, 13]
9'd188: rdata =  56'b00000010110110110100000000000000000000000000000001010110;
//
// shift amount: 10, Lanes IDs: [10, 11, 12, 13]
9'd189: rdata =  56'b00000010110110110100000000000000000000000000000001011010;
//
// shift amount: 14, Lanes IDs: [10, 11, 12, 13]
9'd190: rdata =  56'b00000010110110110100000000000000000000000000000001011110;
//
// shift amount: 2, Lanes IDs: [10, 11, 12, 13]
9'd191: rdata =  56'b00000010110110110100000000000000000000000000000001010010;
//
// read [True, True, True, True]
// ['x(737,)', 'x(738,)', 'x(739,)', 'x(740,)', 'x(541,)', 'x(542,)', 'x(543,)', 'x(544,)', 'x(622,)', 'x(623,)', 'x(625,)', 'x(626,)', 'x(702,)', 'x(703,)', 'x(705,)', 'x(706,)']
// Data values: [-3, 0, -3, 0, -2, -1, -1, 1, 1, 2, 2, -2, 1, 1, 1, -2]
// Dest PEs: [10, 11, 12, 13, 46, 47, 49, 50, 46, 47, 49, 50, 46, 47, 49, 50]
9'd192: rdata =  56'b00000000000000000000000000000000000000000000000000001111;
//
// shift amount: 5, Lanes IDs: [1, 2]
9'd193: rdata =  56'b00000000000000000000000000000000000000011111100001010101;
//
// shift amount: 6, Lanes IDs: [10, 11, 12, 13, 14, 15]
9'd194: rdata =  56'b10110100100100100100000000000000000000000000000001010110;
//
// shift amount: 9, Lanes IDs: [1, 2]
9'd195: rdata =  56'b00000000000000000000000000000000000000011111100001011001;
//
// shift amount: 10, Lanes IDs: [14, 15]
9'd196: rdata =  56'b10110100000000000000000000000000000000000000000001011010;
//
// shift amount: 13, Lanes IDs: [1, 2]
9'd197: rdata =  56'b00000000000000000000000000000000000000011111100001011101;
//
// shift amount: 14, Lanes IDs: [14, 15]
9'd198: rdata =  56'b10110100000000000000000000000000000000000000000001011110;
//
// read [True, True, True, True]
// ['x(742,)', 'x(743,)', 'x(745,)', 'x(746,)', 'x(546,)', 'x(547,)', 'x(549,)', 'x(550,)', 'x(628,)', 'x(629,)', 'x(631,)', 'x(632,)', 'x(708,)', 'x(709,)', 'x(711,)', 'x(712,)']
// Data values: [1, 2, 1, 0, -2, -3, -1, -2, -1, -2, 1, -1, 2, -2, 2, -2]
// Dest PEs: [14, 15, 17, 18, 51, 52, 53, 54, 51, 52, 53, 54, 51, 52, 53, 54]
9'd199: rdata =  56'b00000000000000000000000000000000000000000000000000001111;
//
// shift amount: 1, Lanes IDs: [1, 2, 3, 4, 5, 6]
9'd200: rdata =  56'b00000000000000000000000000011111111111101101100001010001;
//
// shift amount: 2, Lanes IDs: [14, 15]
9'd201: rdata =  56'b00100100000000000000000000000000000000000000000001010010;
//
// shift amount: 5, Lanes IDs: [3, 4, 5, 6]
9'd202: rdata =  56'b00000000000000000000000000011111111111100000000001010101;
//
// shift amount: 9, Lanes IDs: [3, 4, 5, 6]
9'd203: rdata =  56'b00000000000000000000000000011111111111100000000001011001;
//
// read [True, True, True, True]
// ['x(748,)', 'x(749,)', 'x(751,)', 'x(752,)', 'x(110,)', 'x(113,)', 'x(116,)', 'x(119,)', 'x(634,)', 'x(635,)', 'x(637,)', 'x(638,)', 'x(714,)', 'x(715,)', 'x(717,)', 'x(718,)']
// Data values: [2, -2, 2, 2, 1, 1, -2, 0, 2, -1, 1, -1, 0, -1, 1, -2]
// Dest PEs: [19, 20, 21, 22, 19, 20, 21, 22, 55, 57, 58, 59, 55, 57, 58, 59]
9'd204: rdata =  56'b00000000000000000000000000000000000000000000000000001111;
//
// shift amount: 0, Lanes IDs: [9, 10, 11]
9'd205: rdata =  56'b00000000000011111111100000000000000000000000000001010000;
//
// shift amount: 4, Lanes IDs: [9, 10, 11]
9'd206: rdata =  56'b00000000000011111111100000000000000000000000000001010100;
//
// shift amount: 13, Lanes IDs: [3, 4, 5, 6]
9'd207: rdata =  56'b00000000000000000000000000001101101101100000000001011101;
//
// shift amount: 1, Lanes IDs: [3, 4, 5, 6, 7]
9'd208: rdata =  56'b00000000000000000000000011101101101101100000000001010001;
//
// shift amount: 5, Lanes IDs: [7]
9'd209: rdata =  56'b00000000000000000000000011100000000000000000000001010101;
//
// read [True, True, True, True]
// ['x(754,)', 'x(755,)', 'x(757,)', 'x(758,)', 'x(122,)', 'x(125,)', 'x(128,)', 'x(131,)', 'x(639,)', 'x(640,)', 'x(641,)', 'x(642,)', 'x(720,)', 'x(721,)', 'x(723,)', 'x(724,)']
// Data values: [-3, -1, 2, 0, -1, 2, -1, 2, -3, 1, 1, -2, -3, -1, 2, 0]
// Dest PEs: [23, 25, 26, 27, 23, 25, 26, 27, 60, 61, 62, 63, 60, 61, 62, 63]
9'd210: rdata =  56'b00000000000000000000000000000000000000000000000000001111;
//
// shift amount: 8, Lanes IDs: [9, 10, 11]
9'd211: rdata =  56'b00000000000001101101100000000000000000000000000001011000;
//
// shift amount: 9, Lanes IDs: [7]
9'd212: rdata =  56'b00000000000000000000000001100000000000000000000001011001;
//
// shift amount: 12, Lanes IDs: [9, 10, 11, 12, 13, 14, 15]
9'd213: rdata =  56'b11111111111101101101100000000000000000000000000001011100;
//
// shift amount: 0, Lanes IDs: [12, 13, 14, 15]
9'd214: rdata =  56'b11111111111100000000000000000000000000000000000001010000;
//
// shift amount: 13, Lanes IDs: [7]
9'd215: rdata =  56'b00000000000000000000000001100000000000000000000001011101;
//
// read [True, True, True, True]
// ['x(760,)', 'x(761,)', 'x(763,)', 'x(764,)', 'x(134,)', 'x(137,)', 'x(140,)', 'x(143,)', 'x(318,)', 'x(321,)', 'x(324,)', 'x(327,)', 'x(726,)', 'x(727,)', 'x(729,)', 'x(730,)']
// Data values: [-2, 0, -2, 0, -3, -2, -2, 2, 1, -2, -2, 0, 1, 1, 0, 0]
// Dest PEs: [28, 29, 30, 31, 28, 29, 30, 31, 28, 29, 30, 31, 1, 2, 3, 4]
9'd216: rdata =  56'b00000000000000000000000000000000000000000000000000001111;
//
// shift amount: 11, Lanes IDs: [1, 2, 3, 4]
9'd217: rdata =  56'b00000000000000000000000000000000000100100100100001011011;
//
// shift amount: 4, Lanes IDs: [12, 13, 14, 15]
9'd218: rdata =  56'b01101101101100000000000000000000000000000000000001010100;
//
// shift amount: 8, Lanes IDs: [12, 13, 14, 15]
9'd219: rdata =  56'b01101101101100000000000000000000000000000000000001011000;
//
// shift amount: 12, Lanes IDs: [12, 13, 14, 15]
9'd220: rdata =  56'b01101101101100000000000000000000000000000000000001011100;
//
// read [True, True, True, True]
// ['x(766,)', 'x(767,)', 'x(769,)', 'x(770,)', 'x(146,)', 'x(153,)', 'x(156,)', 'x(159,)', 'x(330,)', 'x(333,)', 'x(336,)', 'x(339,)', 'x(732,)', 'x(733,)', 'x(735,)', 'x(736,)']
// Data values: [-1, 1, -2, -2, -2, -3, 1, -3, -3, -3, -2, -3, 2, -2, -2, -3]
// Dest PEs: [33, 34, 35, 36, 33, 34, 35, 36, 33, 34, 35, 36, 5, 6, 7, 9]
9'd221: rdata =  56'b00000000000000000000000000000000000000000000000000001111;
//
// shift amount: 6, Lanes IDs: [9]
9'd222: rdata =  56'b00000000000000000000100000000000000000000000000001010110;
//
// shift amount: 15, Lanes IDs: [1, 2, 3, 4]
9'd223: rdata =  56'b00000000000000000000000000000000010110110110100001011111;
//
// shift amount: 3, Lanes IDs: [1, 2, 3, 4]
9'd224: rdata =  56'b00000000000000000000000000000000010110110110100001010011;
//
// shift amount: 7, Lanes IDs: [1, 2, 3, 4, 5, 6, 7]
9'd225: rdata =  56'b00000000000000000000000000100100110110110110100001010111;
//
// read [True, True, True, True]
// ['x(772,)', 'x(773,)', 'x(775,)', 'x(776,)', 'x(162,)', 'x(165,)', 'x(168,)', 'x(171,)', 'x(342,)', 'x(349,)', 'x(352,)', 'x(355,)', 'x(526,)', 'x(529,)', 'x(532,)', 'x(535,)']
// Data values: [-3, 1, 1, 0, 2, -2, 1, 1, -2, -2, -1, 1, 1, 0, 1, -3]
// Dest PEs: [37, 38, 39, 41, 37, 38, 39, 41, 37, 38, 39, 41, 37, 38, 39, 41]
9'd226: rdata =  56'b00000000000000000000000000000000000000000000000000001111;
//
// shift amount: 10, Lanes IDs: [9]
9'd227: rdata =  56'b00000000000000000010100000000000000000000000000001011010;
//
// shift amount: 11, Lanes IDs: [5, 6, 7]
9'd228: rdata =  56'b00000000000000000000000010110110100000000000000001011011;
//
// shift amount: 14, Lanes IDs: [9]
9'd229: rdata =  56'b00000000000000000010100000000000000000000000000001011110;
//
// shift amount: 2, Lanes IDs: [9]
9'd230: rdata =  56'b00000000000000000010100000000000000000000000000001010010;
//
// shift amount: 6, Lanes IDs: [9]
9'd231: rdata =  56'b00000000000000000010100000000000000000000000000001010110;
//
// shift amount: 15, Lanes IDs: [5, 6, 7]
9'd232: rdata =  56'b00000000000000000000000010110110100000000000000001011111;
//
// shift amount: 3, Lanes IDs: [5, 6, 7]
9'd233: rdata =  56'b00000000000000000000000010110110100000000000000001010011;
//
// shift amount: 7, Lanes IDs: [5, 6, 7]
9'd234: rdata =  56'b00000000000000000000000010110110100000000000000001010111;
//
// read [True, True, True, True]
// ['x(778,)', 'x(779,)', 'x(781,)', 'x(782,)', 'x(174,)', 'x(177,)', 'x(180,)', 'x(183,)', 'x(358,)', 'x(361,)', 'x(364,)', 'x(367,)', 'x(538,)', 'x(545,)', 'x(548,)', 'x(551,)']
// Data values: [1, -3, -2, 0, 1, 0, -2, 2, -1, 1, -3, 1, 0, 2, -1, -3]
// Dest PEs: [42, 43, 44, 45, 42, 43, 44, 45, 42, 43, 44, 45, 42, 43, 44, 45]
9'd235: rdata =  56'b00000000000000000000000000000000000000000000000000001111;
//
// shift amount: 6, Lanes IDs: [10, 11, 12, 13]
9'd236: rdata =  56'b00000010110110110100000000000000000000000000000001010110;
//
// shift amount: 10, Lanes IDs: [10, 11, 12, 13]
9'd237: rdata =  56'b00000010110110110100000000000000000000000000000001011010;
//
// shift amount: 14, Lanes IDs: [10, 11, 12, 13]
9'd238: rdata =  56'b00000010110110110100000000000000000000000000000001011110;
//
// shift amount: 2, Lanes IDs: [10, 11, 12, 13]
9'd239: rdata =  56'b00000010110110110100000000000000000000000000000001010010;
//
// read [True, True, True, True]
// ['x(6,)', 'x(9,)', 'x(12,)', 'x(15,)', 'x(186,)', 'x(189,)', 'x(192,)', 'x(195,)', 'x(370,)', 'x(373,)', 'x(376,)', 'x(379,)', 'x(554,)', 'x(557,)', 'x(560,)', 'x(563,)']
// Data values: [-3, -3, -3, -1, -2, 0, 0, 1, 2, -2, -2, -3, 2, 2, 2, -3]
// Dest PEs: [46, 47, 49, 50, 46, 47, 49, 50, 46, 47, 49, 50, 46, 47, 49, 50]
9'd240: rdata =  56'b00000000000000000000000000000000000000000000000000001111;
//
// shift amount: 1, Lanes IDs: [1, 2]
9'd241: rdata =  56'b00000000000000000000000000000000000000011111100001010001;
//
// shift amount: 2, Lanes IDs: [14, 15]
9'd242: rdata =  56'b10110100000000000000000000000000000000000000000001010010;
//
// shift amount: 5, Lanes IDs: [1, 2]
9'd243: rdata =  56'b00000000000000000000000000000000000000011111100001010101;
//
// shift amount: 6, Lanes IDs: [14, 15]
9'd244: rdata =  56'b10110100000000000000000000000000000000000000000001010110;
//
// shift amount: 9, Lanes IDs: [1, 2]
9'd245: rdata =  56'b00000000000000000000000000000000000000011111100001011001;
//
// shift amount: 10, Lanes IDs: [14, 15]
9'd246: rdata =  56'b10110100000000000000000000000000000000000000000001011010;
//
// shift amount: 13, Lanes IDs: [1, 2]
9'd247: rdata =  56'b00000000000000000000000000000000000000011111100001011101;
//
// shift amount: 14, Lanes IDs: [14, 15]
9'd248: rdata =  56'b10110100000000000000000000000000000000000000000001011110;
//
// read [True, True, True, True]
// ['x(18,)', 'x(21,)', 'x(24,)', 'x(27,)', 'x(202,)', 'x(205,)', 'x(208,)', 'x(211,)', 'x(382,)', 'x(385,)', 'x(388,)', 'x(391,)', 'x(566,)', 'x(569,)', 'x(572,)', 'x(575,)']
// Data values: [-2, 1, 0, 2, -3, -3, 2, -2, 0, -2, -1, -3, -1, 1, -1, 1]
// Dest PEs: [51, 52, 53, 54, 51, 52, 53, 54, 51, 52, 53, 54, 51, 52, 53, 54]
9'd249: rdata =  56'b00000000000000000000000000000000000000000000000000001111;
//
// shift amount: 13, Lanes IDs: [3, 4, 5, 6]
9'd250: rdata =  56'b00000000000000000000000000011111111111100000000001011101;
//
// shift amount: 1, Lanes IDs: [3, 4, 5, 6]
9'd251: rdata =  56'b00000000000000000000000000011111111111100000000001010001;
//
// shift amount: 5, Lanes IDs: [3, 4, 5, 6]
9'd252: rdata =  56'b00000000000000000000000000011111111111100000000001010101;
//
// shift amount: 9, Lanes IDs: [3, 4, 5, 6]
9'd253: rdata =  56'b00000000000000000000000000011111111111100000000001011001;
//
// read [True, True, True, True]
// ['x(30,)', 'x(33,)', 'x(36,)', 'x(39,)', 'x(214,)', 'x(217,)', 'x(220,)', 'x(223,)', 'x(398,)', 'x(401,)', 'x(404,)', 'x(407,)', 'x(578,)', 'x(581,)', 'x(584,)', 'x(587,)']
// Data values: [-3, -2, -2, 0, 1, 1, 1, 2, 2, -3, 0, 2, 0, -2, -2, 2]
// Dest PEs: [55, 57, 58, 59, 55, 57, 58, 59, 55, 57, 58, 59, 55, 57, 58, 59]
9'd254: rdata =  56'b00000000000000000000000000000000000000000000000000001111;
//
// shift amount: 8, Lanes IDs: [9, 10, 11]
9'd255: rdata =  56'b00000000000011111111100000000000000000000000000001011000;
//
// shift amount: 9, Lanes IDs: [7]
9'd256: rdata =  56'b00000000000000000000000011100000000000000000000001011001;
//
// shift amount: 12, Lanes IDs: [9, 10, 11]
9'd257: rdata =  56'b00000000000011111111100000000000000000000000000001011100;
//
// shift amount: 0, Lanes IDs: [9, 10, 11]
9'd258: rdata =  56'b00000000000011111111100000000000000000000000000001010000;
//
// shift amount: 4, Lanes IDs: [9, 10, 11]
9'd259: rdata =  56'b00000000000011111111100000000000000000000000000001010100;
//
// shift amount: 13, Lanes IDs: [7]
9'd260: rdata =  56'b00000000000000000000000011100000000000000000000001011101;
//
// shift amount: 1, Lanes IDs: [7]
9'd261: rdata =  56'b00000000000000000000000011100000000000000000000001010001;
//
// shift amount: 5, Lanes IDs: [7]
9'd262: rdata =  56'b00000000000000000000000011100000000000000000000001010101;
//
// read [True, True, True, True]
// ['x(42,)', 'x(45,)', 'x(48,)', 'x(55,)', 'x(226,)', 'x(229,)', 'x(232,)', 'x(235,)', 'x(410,)', 'x(413,)', 'x(416,)', 'x(419,)', 'x(594,)', 'x(597,)', 'x(600,)', 'x(603,)']
// Data values: [-1, -3, 2, -2, 2, -1, 0, 0, 1, 0, -2, -2, -1, 2, 0, -1]
// Dest PEs: [60, 61, 62, 63, 60, 61, 62, 63, 60, 61, 62, 63, 60, 61, 62, 63]
9'd263: rdata =  56'b00000000000000000000000000000000000000000000000000001111;
//
// shift amount: 4, Lanes IDs: [12, 13, 14, 15]
9'd264: rdata =  56'b11111111111100000000000000000000000000000000000001010100;
//
// shift amount: 8, Lanes IDs: [12, 13, 14, 15]
9'd265: rdata =  56'b11111111111100000000000000000000000000000000000001011000;
//
// shift amount: 12, Lanes IDs: [12, 13, 14, 15]
9'd266: rdata =  56'b11111111111100000000000000000000000000000000000001011100;
//
// shift amount: 0, Lanes IDs: [12, 13, 14, 15]
9'd267: rdata =  56'b11111111111100000000000000000000000000000000000001010000;
//
// read [True, True, True, True]
// ['x(58,)', 'x(61,)', 'x(64,)', 'x(67,)', 'x(238,)', 'x(241,)', 'x(244,)', 'x(251,)', 'x(422,)', 'x(425,)', 'x(428,)', 'x(431,)', 'x(606,)', 'x(609,)', 'x(612,)', 'x(615,)']
// Data values: [0, -3, 0, -1, -2, 2, 1, -3, 2, 0, -2, -2, -3, -3, -2, 2]
// Dest PEs: [1, 2, 3, 4, 1, 2, 3, 4, 1, 2, 3, 4, 1, 2, 3, 4]
9'd268: rdata =  56'b00000000000000000000000000000000000000000000000000001111;
//
// shift amount: 15, Lanes IDs: [1, 2, 3, 4]
9'd269: rdata =  56'b00000000000000000000000000000000000100100100100001011111;
//
// shift amount: 3, Lanes IDs: [1, 2, 3, 4]
9'd270: rdata =  56'b00000000000000000000000000000000000100100100100001010011;
//
// shift amount: 7, Lanes IDs: [1, 2, 3, 4]
9'd271: rdata =  56'b00000000000000000000000000000000000100100100100001010111;
//
// shift amount: 11, Lanes IDs: [1, 2, 3, 4]
9'd272: rdata =  56'b00000000000000000000000000000000000100100100100001011011;
//
// read [True, True, True, True]
// ['x(70,)', 'x(73,)', 'x(76,)', 'x(79,)', 'x(254,)', 'x(257,)', 'x(260,)', 'x(263,)', 'x(434,)', 'x(437,)', 'x(440,)', 'x(447,)', 'x(618,)', 'x(621,)', 'x(624,)', 'x(627,)']
// Data values: [-2, 0, 2, -3, -3, -1, 1, -2, 0, 2, -2, 1, -2, -1, 1, -3]
// Dest PEs: [5, 6, 7, 9, 5, 6, 7, 9, 5, 6, 7, 9, 5, 6, 7, 9]
9'd273: rdata =  56'b00000000000000000000000000000000000000000000000000001111;
//
// shift amount: 10, Lanes IDs: [9]
9'd274: rdata =  56'b00000000000000000000100000000000000000000000000001011010;
//
// shift amount: 11, Lanes IDs: [5, 6, 7]
9'd275: rdata =  56'b00000000000000000000000000100100100000000000000001011011;
//
// shift amount: 14, Lanes IDs: [9]
9'd276: rdata =  56'b00000000000000000000100000000000000000000000000001011110;
//
// shift amount: 2, Lanes IDs: [9]
9'd277: rdata =  56'b00000000000000000000100000000000000000000000000001010010;
//
// shift amount: 6, Lanes IDs: [9]
9'd278: rdata =  56'b00000000000000000000100000000000000000000000000001010110;
//
// shift amount: 15, Lanes IDs: [5, 6, 7]
9'd279: rdata =  56'b00000000000000000000000000100100100000000000000001011111;
//
// shift amount: 3, Lanes IDs: [5, 6, 7]
9'd280: rdata =  56'b00000000000000000000000000100100100000000000000001010011;
//
// shift amount: 7, Lanes IDs: [5, 6, 7]
9'd281: rdata =  56'b00000000000000000000000000100100100000000000000001010111;
//
// read [True, True, True, True]
// ['x(82,)', 'x(85,)', 'x(88,)', 'x(91,)', 'x(266,)', 'x(269,)', 'x(272,)', 'x(275,)', 'x(450,)', 'x(453,)', 'x(456,)', 'x(459,)', 'x(630,)', 'x(633,)', 'x(636,)', 'x(643,)']
// Data values: [-3, 2, 1, -3, 2, -3, 0, -2, 1, 1, 2, 1, 1, -1, 1, 1]
// Dest PEs: [10, 11, 12, 13, 10, 11, 12, 13, 10, 11, 12, 13, 10, 11, 12, 13]
9'd282: rdata =  56'b00000000000000000000000000000000000000000000000000001111;
//
// shift amount: 6, Lanes IDs: [10, 11, 12, 13]
9'd283: rdata =  56'b00000000100100100100000000000000000000000000000001010110;
//
// shift amount: 10, Lanes IDs: [10, 11, 12, 13]
9'd284: rdata =  56'b00000000100100100100000000000000000000000000000001011010;
//
// shift amount: 14, Lanes IDs: [10, 11, 12, 13]
9'd285: rdata =  56'b00000000100100100100000000000000000000000000000001011110;
//
// shift amount: 2, Lanes IDs: [10, 11, 12, 13]
9'd286: rdata =  56'b00000000100100100100000000000000000000000000000001010010;
//
// read [True, True, True, True]
// ['x(94,)', 'x(97,)', 'x(104,)', 'x(107,)', 'x(278,)', 'x(281,)', 'x(284,)', 'x(287,)', 'x(462,)', 'x(465,)', 'x(468,)', 'x(471,)', 'x(646,)', 'x(649,)', 'x(652,)', 'x(655,)']
// Data values: [2, -3, 2, -1, 2, 0, 1, -1, -1, -2, -1, 0, 0, 2, -1, 0]
// Dest PEs: [14, 15, 17, 18, 14, 15, 17, 18, 14, 15, 17, 18, 14, 15, 17, 18]
9'd287: rdata =  56'b00000000000000000000000000000000000000000000000000001111;
//
// shift amount: 1, Lanes IDs: [1, 2]
9'd288: rdata =  56'b00000000000000000000000000000000000000001101100001010001;
//
// shift amount: 2, Lanes IDs: [14, 15]
9'd289: rdata =  56'b00100100000000000000000000000000000000000000000001010010;
//
// shift amount: 5, Lanes IDs: [1, 2]
9'd290: rdata =  56'b00000000000000000000000000000000000000001101100001010101;
//
// shift amount: 6, Lanes IDs: [14, 15]
9'd291: rdata =  56'b00100100000000000000000000000000000000000000000001010110;
//
// shift amount: 9, Lanes IDs: [1, 2]
9'd292: rdata =  56'b00000000000000000000000000000000000000001101100001011001;
//
// shift amount: 10, Lanes IDs: [14, 15]
9'd293: rdata =  56'b00100100000000000000000000000000000000000000000001011010;
//
// shift amount: 13, Lanes IDs: [1, 2]
9'd294: rdata =  56'b00000000000000000000000000000000000000001101100001011101;
//
// shift amount: 14, Lanes IDs: [14, 15]
9'd295: rdata =  56'b00100100000000000000000000000000000000000000000001011110;
//
// read [True, True, True, True]
// ['x(734,)', 'x(741,)', 'x(744,)', 'x(747,)', 'x(290,)', 'x(293,)', 'x(300,)', 'x(303,)', 'x(474,)', 'x(477,)', 'x(480,)', 'x(483,)', 'x(658,)', 'x(661,)', 'x(664,)', 'x(667,)']
// Data values: [2, -2, 2, 2, -2, 1, 1, 2, 2, -1, -2, 0, 1, 0, 1, 0]
// Dest PEs: [46, 47, 49, 50, 19, 20, 21, 22, 19, 20, 21, 22, 19, 20, 21, 22]
9'd296: rdata =  56'b00000000000000000000000000000000000000000000000000001111;
//
// shift amount: 1, Lanes IDs: [1, 2, 3, 4, 5, 6]
9'd297: rdata =  56'b00000000000000000000000000001101101101111111100001010001;
//
// shift amount: 2, Lanes IDs: [14, 15]
9'd298: rdata =  56'b10110100000000000000000000000000000000000000000001010010;
//
// shift amount: 5, Lanes IDs: [3, 4, 5, 6]
9'd299: rdata =  56'b00000000000000000000000000001101101101100000000001010101;
//
// shift amount: 9, Lanes IDs: [3, 4, 5, 6]
9'd300: rdata =  56'b00000000000000000000000000001101101101100000000001011001;
//
// read [True, True, True, True]
// ['x(750,)', 'x(753,)', 'x(756,)', 'x(759,)', 'x(306,)', 'x(309,)', 'x(312,)', 'x(315,)', 'x(486,)', 'x(489,)', 'x(496,)', 'x(499,)', 'x(670,)', 'x(673,)', 'x(676,)', 'x(679,)']
// Data values: [-2, -2, 2, 1, 2, -3, -1, 2, 0, 0, 0, -1, -1, -1, 2, -1]
// Dest PEs: [51, 52, 53, 54, 23, 25, 26, 27, 23, 25, 26, 27, 23, 25, 26, 27]
9'd301: rdata =  56'b00000000000000000000000000000000000000000000000000001111;
//
// shift amount: 12, Lanes IDs: [9, 10, 11]
9'd302: rdata =  56'b00000000000001101101100000000000000000000000000001011100;
//
// shift amount: 0, Lanes IDs: [9, 10, 11]
9'd303: rdata =  56'b00000000000001101101100000000000000000000000000001010000;
//
// shift amount: 4, Lanes IDs: [9, 10, 11]
9'd304: rdata =  56'b00000000000001101101100000000000000000000000000001010100;
//
// shift amount: 13, Lanes IDs: [3, 4, 5, 6, 7]
9'd305: rdata =  56'b00000000000000000000000001111111111111100000000001011101;
//
// shift amount: 1, Lanes IDs: [7]
9'd306: rdata =  56'b00000000000000000000000001100000000000000000000001010001;
//
// shift amount: 5, Lanes IDs: [7]
9'd307: rdata =  56'b00000000000000000000000001100000000000000000000001010101;
//
// read [True, False, True, True]
// ['x(762,)', 'x(765,)', 'x(768,)', 'x(771,)', None, None, None, None, 'x(502,)', 'x(505,)', 'x(508,)', 'x(511,)', 'x(682,)', 'x(685,)', 'x(692,)', 'x(695,)']
// Data values: [1, 0, 2, 0, None, None, None, None, -1, 2, -2, 1, 0, 2, 2, 1]
// Dest PEs: [55, 57, 58, 59, None, None, None, None, 28, 29, 30, 31, 28, 29, 30, 31]
9'd308: rdata =  56'b00000000000000000000000000000000000000000000000000001101;
//
// shift amount: 8, Lanes IDs: [9, 10, 11]
9'd309: rdata =  56'b00000000000011111111100000000000000000000000000001011000;
//
// shift amount: 9, Lanes IDs: [7]
9'd310: rdata =  56'b00000000000000000000000011100000000000000000000001011001;
//
// shift amount: 12, Lanes IDs: [12, 13, 14, 15]
9'd311: rdata =  56'b01101101101100000000000000000000000000000000000001011100;
//
// shift amount: 0, Lanes IDs: [12, 13, 14, 15]
9'd312: rdata =  56'b01101101101100000000000000000000000000000000000001010000;
//
// read [True, False, True, True]
// ['x(774,)', 'x(777,)', 'x(780,)', 'x(783,)', None, None, None, None, 'x(514,)', 'x(517,)', 'x(520,)', 'x(523,)', 'x(698,)', 'x(701,)', 'x(704,)', 'x(707,)']
// Data values: [1, 1, -1, 0, None, None, None, None, 2, 1, 2, 2, 2, -2, 0, 0]
// Dest PEs: [60, 61, 62, 63, None, None, None, None, 33, 34, 35, 36, 33, 34, 35, 36]
9'd313: rdata =  56'b00000000000000000000000000000000000000000000000000001101;
//
// shift amount: 4, Lanes IDs: [12, 13, 14, 15]
9'd314: rdata =  56'b11111111111100000000000000000000000000000000000001010100;
//
// shift amount: 7, Lanes IDs: [1, 2, 3, 4]
9'd315: rdata =  56'b00000000000000000000000000000000010110110110100001010111;
//
// shift amount: 11, Lanes IDs: [1, 2, 3, 4]
9'd316: rdata =  56'b00000000000000000000000000000000010110110110100001011011;
//
// read [True, False, False, True]
// ['y', None, None, None, None, None, None, None, None, None, None, None, 'x(710,)', 'x(713,)', 'x(716,)', 'x(719,)']
// Data values: [2, None, None, None, None, None, None, None, None, None, None, None, -3, 1, 0, -2]
// Dest PEs: [10, None, None, None, None, None, None, None, None, None, None, None, 37, 38, 39, 41]
9'd317: rdata =  56'b00000000000000000000000000000000000000000000000000001001;
//
// shift amount: 6, Lanes IDs: [9, 10]
9'd318: rdata =  56'b00000000000000000110100000000000000000000000000001010110;
//
// shift amount: 7, Lanes IDs: [5, 6, 7]
9'd319: rdata =  56'b00000000000000000000000010110110100000000000000001010111;
//
// read [False, False, False, True]
// [None, None, None, None, None, None, None, None, None, None, None, None, 'x(722,)', 'x(725,)', 'x(728,)', 'x(731,)']
// Data values: [None, None, None, None, None, None, None, None, None, None, None, None, 1, 0, -1, -1]
// Dest PEs: [None, None, None, None, None, None, None, None, None, None, None, None, 42, 43, 44, 45]
9'd320: rdata =  56'b00000000000000000000000000000000000000000000000000001000;
//
// shift amount: 2, Lanes IDs: [10, 11, 12, 13]
9'd321: rdata =  56'b00000010110110110100000000000000000000000000000001010010;
//
// wfi
9'd322: rdata =  56'b00000000000000000000000000000000000000000000000001100000;
//
// loop
9'd323: rdata =  56'b00000000000000000000000000000000000000000000000001110000;/****************************************************************************************/
default: rdata = 56'b00000000000000000000000000000000000000000000000001110000;

	endcase
	end

    //reg     [ADDR_WIDTH-1:0]        address;

// ******************************************************************
// Read Logic
// ******************************************************************

    always @ (posedge CLK)
    begin : READ_VALID
        if (RESET) begin
            DATA_OUT_VALID <= 1'b0;
        end else if (ENABLE) begin
            DATA_OUT_VALID <= 1'b1;
        end
    end



 always @(posedge CLK) begin
    if (ENABLE)
        DATA_OUT <= rdata;
end

endmodule
