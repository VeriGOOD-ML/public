`define INPUT_BITWIDTH 8
`define BITWIDTH 16
`define NUM_CYCLE 4
`define LOG_NUM_CYCLE 2
`define SIZE 35
`define NUMBER_UNIT 10
`define INST_BITWIDTH 3

//`define SVM 1
//`define LINEAR 1
//`define LOGISTIC 1
`define RECO 1
