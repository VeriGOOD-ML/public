`define WEIGHT_COUNT_MACRO(lanes,pe) (\
(lanes == 0 && pe == 0) ? 16'd0 : \
(lanes == 0 && pe == 1) ? 16'd0 : \
(lanes == 0 && pe == 2) ? 16'd0 : \
(lanes == 0 && pe == 3) ? 16'd0 : \
(lanes == 0 && pe == 4) ? 16'd0 : \
(lanes == 1 && pe == 0) ? 16'd269 : \
(lanes == 1 && pe == 1) ? 16'd140 : \
(lanes == 1 && pe == 2) ? 16'd141 : \
(lanes == 1 && pe == 3) ? 16'd141 : \
(lanes == 1 && pe == 4) ? 16'd691 : \
(lanes == 2 && pe == 0) ? 16'd328 : \
(lanes == 2 && pe == 1) ? 16'd216 : \
(lanes == 2 && pe == 2) ? 16'd156 : \
(lanes == 2 && pe == 3) ? 16'd193 : \
(lanes == 2 && pe == 4) ? 16'd893 : \
(lanes == 3 && pe == 0) ? 16'd293 : \
(lanes == 3 && pe == 1) ? 16'd146 : \
(lanes == 3 && pe == 2) ? 16'd187 : \
(lanes == 3 && pe == 3) ? 16'd165 : \
(lanes == 3 && pe == 4) ? 16'd791 : \
(lanes == 4 && pe == 0) ? 16'd266 : \
(lanes == 4 && pe == 1) ? 16'd135 : \
(lanes == 4 && pe == 2) ? 16'd152 : \
(lanes == 4 && pe == 3) ? 16'd140 : \
(lanes == 4 && pe == 4) ? 16'd693 : \
(lanes == 5 && pe == 0) ? 16'd265 : \
(lanes == 5 && pe == 1) ? 16'd129 : \
(lanes == 5 && pe == 2) ? 16'd143 : \
(lanes == 5 && pe == 3) ? 16'd140 : \
(lanes == 5 && pe == 4) ? 16'd677 : \
(lanes == 6 && pe == 0) ? 16'd266 : \
(lanes == 6 && pe == 1) ? 16'd137 : \
(lanes == 6 && pe == 2) ? 16'd152 : \
(lanes == 6 && pe == 3) ? 16'd138 : \
(lanes == 6 && pe == 4) ? 16'd693 : \
(lanes == 7 && pe == 0) ? 16'd265 : \
(lanes == 7 && pe == 1) ? 16'd133 : \
(lanes == 7 && pe == 2) ? 16'd143 : \
(lanes == 7 && pe == 3) ? 16'd139 : \
(lanes == 7 && pe == 4) ? 16'd680 : \
(lanes == 8 && pe == 0) ? 16'd0 : \
(lanes == 8 && pe == 1) ? 16'd0 : \
(lanes == 8 && pe == 2) ? 16'd0 : \
(lanes == 8 && pe == 3) ? 16'd0 : \
(lanes == 8 && pe == 4) ? 16'd0 : \
(lanes == 9 && pe == 0) ? 16'd268 : \
(lanes == 9 && pe == 1) ? 16'd143 : \
(lanes == 9 && pe == 2) ? 16'd143 : \
(lanes == 9 && pe == 3) ? 16'd139 : \
(lanes == 9 && pe == 4) ? 16'd693 : \
(lanes == 10 && pe == 0) ? 16'd186 : \
(lanes == 10 && pe == 1) ? 16'd173 : \
(lanes == 10 && pe == 2) ? 16'd234 : \
(lanes == 10 && pe == 3) ? 16'd229 : \
(lanes == 10 && pe == 4) ? 16'd822 : \
(lanes == 11 && pe == 0) ? 16'd165 : \
(lanes == 11 && pe == 1) ? 16'd182 : \
(lanes == 11 && pe == 2) ? 16'd146 : \
(lanes == 11 && pe == 3) ? 16'd147 : \
(lanes == 11 && pe == 4) ? 16'd640 : \
(lanes == 12 && pe == 0) ? 16'd147 : \
(lanes == 12 && pe == 1) ? 16'd139 : \
(lanes == 12 && pe == 2) ? 16'd135 : \
(lanes == 12 && pe == 3) ? 16'd137 : \
(lanes == 12 && pe == 4) ? 16'd558 : \
(lanes == 13 && pe == 0) ? 16'd141 : \
(lanes == 13 && pe == 1) ? 16'd139 : \
(lanes == 13 && pe == 2) ? 16'd141 : \
(lanes == 13 && pe == 3) ? 16'd136 : \
(lanes == 13 && pe == 4) ? 16'd557 : \
(lanes == 14 && pe == 0) ? 16'd130 : \
(lanes == 14 && pe == 1) ? 16'd139 : \
(lanes == 14 && pe == 2) ? 16'd128 : \
(lanes == 14 && pe == 3) ? 16'd130 : \
(lanes == 14 && pe == 4) ? 16'd527 : \
(lanes == 15 && pe == 0) ? 16'd147 : \
(lanes == 15 && pe == 1) ? 16'd141 : \
(lanes == 15 && pe == 2) ? 16'd131 : \
(lanes == 15 && pe == 3) ? 16'd138 : \
16'd557)