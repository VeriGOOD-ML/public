`define INPUT_BITWIDTH 16
`define BITWIDTH 32
`define NUM_CYCLE 4
`define LOG_NUM_CYCLE 2
`define SIZE 14
`define NUM_UNIT 1

`define SVM 1