`timescale 1ns/1ps
module decoder #( parameter inputLen = 3,
	parameter outputLen = 1 << inputLen 
	)(
	in , 
 	decoder_out 
);

	//--------------------------------------------------------------------------------------
	
	//--------------------------------------------------------------------------------------
	
	//--------------------------------------------------------------------------------------
	input [inputLen - 1 : 0] in;
	output [outputLen - 1 : 0] decoder_out ; 
    //--------------------------------------------------------------------------------------
    
    //-------------------------------------------------------------------------------------- 	
	assign decoder_out = (1 << in) ;
	//--------------------------------------------------------------------------------------
	
endmodule
