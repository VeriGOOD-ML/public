`define INPUT_BITWIDTH 16
`define BITWIDTH 32
`define NUM_CYCLE 25
`define LOG_NUM_CYCLE 5
`define SIZE 10
`define NUMBER_UNIT 10
`define INST_BITWIDTH 3
`define IP_NUM_STAGE 0
`define SGD_NUM_STAGE 0

//`define SVM 1
//`define LINEAR 1
//`define LOGISTIC 1
`define RECO 1
