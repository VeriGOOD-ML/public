`define INPUT_BITWIDTH
`define BITWIDTH
`define NUM_CYCLE
`define LOG_NUM_CYCLE
`define SIZE

//`define SVM 1
//`define LINEAR 1
//`define LOGISTIC 1
//`define RECO 1