`timescale 1ns/1ps

module iBuffer_ASIC #(
    parameter integer addrLen = 5,
	parameter integer dataLen = 32,
	parameter integer peId	= 1
)(
	clk,
	rdAddr,
	noStall,
	dataOut
);

	input clk;
	input noStall;
	input[addrLen - 1: 0] rdAddr;
	output reg[dataLen - 1: 0] dataOut;

	//--------------------------------------------------------------------------------------
	reg[dataLen - 1: 0] mem	[0: (1 << addrLen) - 1];
	
	// ******************************************************************
	// Initialization
	// ******************************************************************

    localparam DATA_WIDTH = dataLen;
    localparam DEPTH = (1<<addrLen);
    wire     [addrLen-1:0]        address;
    reg     [DATA_WIDTH-1:0]        rdata;

    assign address = rdAddr;
	
	always @(posedge clk) begin
 		if(noStall) dataOut <= rdata;
	end
	
    // `include "instructions.v" // TODO

	//-------------------------------------------------------------------------------------
 	
generate
if(peId == 0) begin
	always @(*) begin
		case(address)
			4'd0 : rdata = 55'b0001101000000000011000000001000000000000000000000000000;
			4'd1 : rdata = 55'b1100011011111110000000000000000000000000000001000000000;
			4'd2 : rdata = 55'b1100011100001100000000000000000000000000000001000000000;
			4'd3 : rdata = 55'b0000111100000110101000000001000000010000000000000000000;
			4'd4 : rdata = 55'b0001110100000001011000000011000000100000000000000000000;
			4'd5 : rdata = 55'b0001010100000010011000000101000000110000000000100000000;
			4'd6 : rdata = 55'b0001110100000011011000000001000001000000000000000000000;
			4'd7 : rdata = 55'b0001110000000000101000001001000001010000000000000000000;
			4'd8 : rdata = 55'b0001001000000000101000001010000000001000000000000000000;
			4'd9 : rdata = 55'b1100011100000011000000000000000000000000000000011111111;
			4'd10 : rdata = 55'b1100011100000011000000000000000000000000000000011101110;
			default : rdata = 55'b0000000000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 1) begin
	always @(*) begin
		case(address)
			4'd0 : rdata = 55'b0001101000000000011000000001000000000000000000000000000;
			4'd1 : rdata = 55'b0000111100001000101000000001000000010000000000000000000;
			4'd2 : rdata = 55'b0001110100000001011000000101000000100000000000000000000;
			4'd3 : rdata = 55'b0001010100000010011000000111000010010000000000100000000;
			4'd4 : rdata = 55'b1100010100000011000000000000000000000000000000100000000;
			4'd5 : rdata = 55'b0001111011111110011000000011000001000000000000000000000;
			4'd6 : rdata = 55'b0001110000000000101000001001000001010000000000000000000;
			4'd7 : rdata = 55'b0001001000000001101000001010000000001000000010010111011;
			4'd8 : rdata = 55'b1100011100000100000000000000000000001000000000000000000;
			default : rdata = 55'b0000000000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 2) begin
	always @(*) begin
		case(address)
			4'd0 : rdata = 55'b0001101000000000011000000001000000000000000000000000000;
			4'd1 : rdata = 55'b0000111100001010101000000001000000010000000000000000000;
			4'd2 : rdata = 55'b0001110100000001011000000101000000100000000000000000000;
			4'd3 : rdata = 55'b0001010100000010011000000111000011110000000000100000000;
			4'd4 : rdata = 55'b1100010100000011000000000000000000000000000000100000000;
			4'd5 : rdata = 55'b0001111011111110011000000001000001000000000000000000000;
			4'd6 : rdata = 55'b0001111011111110011000000011000001100000000000000000000;
			4'd7 : rdata = 55'b0001110000000000101000001001000001010000000000000000000;
			4'd8 : rdata = 55'b0001110000000000101000001101000001110000000000000000000;
			4'd9 : rdata = 55'b0001001000000001101000001010000000001000000010010011001;
			4'd10 : rdata = 55'b0001001000000010101000001110000000001000000100011001100;
			4'd11 : rdata = 55'b1100011100000110000000000000000000001000000000000000000;
			default : rdata = 55'b0000000000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 3) begin
	always @(*) begin
		case(address)
			4'd0 : rdata = 55'b0001101000000000011000000000000000000000000000010001000;
			4'd1 : rdata = 55'b0001111011111110011000000011000000000000000000000000000;
			4'd2 : rdata = 55'b0001111011111110011000000001000000100000000000000000000;
			4'd3 : rdata = 55'b0001110000000000101000000001000000010000000000000000000;
			4'd4 : rdata = 55'b0001110000000000101000000101000000110000000000000000000;
			4'd5 : rdata = 55'b0001001000000001101000000010000000001000000010010101010;
			4'd6 : rdata = 55'b0001001000000010101000000110000000001000000100011011101;
			4'd7 : rdata = 55'b1100011100000010000000000000000000001000000000000000000;
			default : rdata = 55'b0000000000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 4) begin
	always @(*) begin
		case(address)
			4'd0 : rdata = 55'b0001101000000000011000000000000000000000000000010011001;
			4'd1 : rdata = 55'b1100011100000100000000000000000000001000000000000000000;
			default : rdata = 55'b0000000000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 5) begin
	always @(*) begin
		case(address)
			4'd0 : rdata = 55'b0001101000000000011000000000000000000000000000010101010;
			4'd1 : rdata = 55'b1100011100000110000000000000000000001000000000000000000;
			default : rdata = 55'b0000000000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 6) begin
	always @(*) begin
		case(address)
			4'd0 : rdata = 55'b0001101100000000010000000000000000000000000000010001000;
			4'd1 : rdata = 55'b1100011100000000000000000000000000001000000000000000000;
			default : rdata = 55'b0000000000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 7) begin
	always @(*) begin
		case(address)
			4'd0 : rdata = 55'b0001101100000000010000000000000000000000000000100000000;
			4'd1 : rdata = 55'b1100011100000000000000000000000000001000000000000000000;
			default : rdata = 55'b0000000000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 8) begin
	always @(*) begin
		case(address)
			4'd0 : rdata = 55'b0001101100000000010000000000000000000000000000100000000;
			4'd1 : rdata = 55'b0000111100000100110111111111000000110000000000000000000;
			4'd2 : rdata = 55'b0000111100000010110111111111000000000000000000000000000;
			4'd3 : rdata = 55'b0001110100000011011000000111000001000000000000000000000;
			4'd4 : rdata = 55'b0001110100000000011000000011000000010000000000000000000;
			4'd5 : rdata = 55'b0001010100000100011000001001000001010000000000100000000;
			4'd6 : rdata = 55'b0001010100000001011000000101000000100000000000100000000;
			4'd7 : rdata = 55'b0001110100000101011000000001000010000000000000000000000;
			4'd8 : rdata = 55'b0001110100000010011000000001000001100000000000000000000;
			4'd9 : rdata = 55'b0001110000000000101000010001000010010000000000000000000;
			4'd10 : rdata = 55'b0001110000000000101000001101000001110000000000000000000;
			4'd11 : rdata = 55'b0001001000000010101000010010000000001000000100000000000;
			4'd12 : rdata = 55'b0001001000000001101000001110000000001000000010000000000;
			4'd13 : rdata = 55'b1100011100000100000000000000000000001000000000000000000;
			default : rdata = 55'b0000000000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 9) begin
	always @(*) begin
		case(address)
			4'd0 : rdata = 55'b0001101100000000010000000000000000000000000000010001000;
			4'd1 : rdata = 55'b0000111100000110110111111101000000000000000000000000000;
			4'd2 : rdata = 55'b0001110100000000011000000011000000010000000000000000000;
			4'd3 : rdata = 55'b0001010100000001011000000101010000110000000000100000000;
			4'd4 : rdata = 55'b1100010100000010000000000000000000000000000000100000000;
			4'd5 : rdata = 55'b0001111011111110011000000001000001010000000000000000000;
			4'd6 : rdata = 55'b0001111011111110011000000001000000110000000000000000000;
			4'd7 : rdata = 55'b0001110000000000101000001011000001100000000000000000000;
			4'd8 : rdata = 55'b0001110000000000101000000111000001000000000000000000000;
			4'd9 : rdata = 55'b0001001000000001101000001100000000001000000010100000000;
			4'd10 : rdata = 55'b0001001000000000101000001000000000001000000000000000000;
			default : rdata = 55'b0000000000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 10) begin
	always @(*) begin
		case(address)
			4'd0 : rdata = 55'b0001101100000000010000000000000000000000000000010001000;
			4'd1 : rdata = 55'b0001111011111110011000000011000000000000000000000000000;
			4'd2 : rdata = 55'b0001111011111110011000000001000000100000000000000000000;
			4'd3 : rdata = 55'b0001110000000000101000000001000000010000000000000000000;
			4'd4 : rdata = 55'b0001110000000000101000000101000000110000000000000000000;
			4'd5 : rdata = 55'b0001001000000001101000000010000000001000000010010001000;
			4'd6 : rdata = 55'b0001001000000010101000000110000000001000000100100000000;
			4'd7 : rdata = 55'b1100011011111110000000000000000000001000000000000000000;
			default : rdata = 55'b0000000000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 11) begin
	always @(*) begin
		case(address)
			4'd0 : rdata = 55'b0001101100000000010000000000000000000000000000010011001;
			4'd1 : rdata = 55'b1100011011111110000000000000000000001000000000000000000;
			default : rdata = 55'b0000000000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 12) begin
	always @(*) begin
		case(address)
			default : rdata = 55'b0000000000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 13) begin
	always @(*) begin
		case(address)
			default : rdata = 55'b0000000000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 14) begin
	always @(*) begin
		case(address)
			default : rdata = 55'b0000000000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 15) begin
	always @(*) begin
		case(address)
			default : rdata = 55'b0000000000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 16) begin
	always @(*) begin
		case(address)
			default : rdata = 55'b0000000000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 17) begin
	always @(*) begin
		case(address)
			default : rdata = 55'b0000000000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 18) begin
	always @(*) begin
		case(address)
			default : rdata = 55'b0000000000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 19) begin
	always @(*) begin
		case(address)
			default : rdata = 55'b0000000000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 20) begin
	always @(*) begin
		case(address)
			default : rdata = 55'b0000000000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 21) begin
	always @(*) begin
		case(address)
			default : rdata = 55'b0000000000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 22) begin
	always @(*) begin
		case(address)
			default : rdata = 55'b0000000000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 23) begin
	always @(*) begin
		case(address)
			default : rdata = 55'b0000000000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 24) begin
	always @(*) begin
		case(address)
			default : rdata = 55'b0000000000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 25) begin
	always @(*) begin
		case(address)
			default : rdata = 55'b0000000000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 26) begin
	always @(*) begin
		case(address)
			default : rdata = 55'b0000000000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 27) begin
	always @(*) begin
		case(address)
			default : rdata = 55'b0000000000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 28) begin
	always @(*) begin
		case(address)
			default : rdata = 55'b0000000000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 29) begin
	always @(*) begin
		case(address)
			default : rdata = 55'b0000000000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 30) begin
	always @(*) begin
		case(address)
			default : rdata = 55'b0000000000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 31) begin
	always @(*) begin
		case(address)
			default : rdata = 55'b0000000000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 32) begin
	always @(*) begin
		case(address)
			default : rdata = 55'b0000000000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 33) begin
	always @(*) begin
		case(address)
			default : rdata = 55'b0000000000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 34) begin
	always @(*) begin
		case(address)
			default : rdata = 55'b0000000000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 35) begin
	always @(*) begin
		case(address)
			default : rdata = 55'b0000000000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 36) begin
	always @(*) begin
		case(address)
			default : rdata = 55'b0000000000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 37) begin
	always @(*) begin
		case(address)
			default : rdata = 55'b0000000000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 38) begin
	always @(*) begin
		case(address)
			default : rdata = 55'b0000000000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 39) begin
	always @(*) begin
		case(address)
			default : rdata = 55'b0000000000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 40) begin
	always @(*) begin
		case(address)
			default : rdata = 55'b0000000000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 41) begin
	always @(*) begin
		case(address)
			default : rdata = 55'b0000000000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 42) begin
	always @(*) begin
		case(address)
			default : rdata = 55'b0000000000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 43) begin
	always @(*) begin
		case(address)
			default : rdata = 55'b0000000000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 44) begin
	always @(*) begin
		case(address)
			default : rdata = 55'b0000000000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 45) begin
	always @(*) begin
		case(address)
			default : rdata = 55'b0000000000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 46) begin
	always @(*) begin
		case(address)
			default : rdata = 55'b0000000000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 47) begin
	always @(*) begin
		case(address)
			default : rdata = 55'b0000000000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 48) begin
	always @(*) begin
		case(address)
			default : rdata = 55'b0000000000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 49) begin
	always @(*) begin
		case(address)
			default : rdata = 55'b0000000000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 50) begin
	always @(*) begin
		case(address)
			default : rdata = 55'b0000000000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 51) begin
	always @(*) begin
		case(address)
			default : rdata = 55'b0000000000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 52) begin
	always @(*) begin
		case(address)
			default : rdata = 55'b0000000000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 53) begin
	always @(*) begin
		case(address)
			default : rdata = 55'b0000000000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 54) begin
	always @(*) begin
		case(address)
			default : rdata = 55'b0000000000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 55) begin
	always @(*) begin
		case(address)
			default : rdata = 55'b0000000000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 56) begin
	always @(*) begin
		case(address)
			default : rdata = 55'b0000000000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 57) begin
	always @(*) begin
		case(address)
			default : rdata = 55'b0000000000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 58) begin
	always @(*) begin
		case(address)
			default : rdata = 55'b0000000000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 59) begin
	always @(*) begin
		case(address)
			default : rdata = 55'b0000000000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 60) begin
	always @(*) begin
		case(address)
			default : rdata = 55'b0000000000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 61) begin
	always @(*) begin
		case(address)
			default : rdata = 55'b0000000000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 62) begin
	always @(*) begin
		case(address)
			default : rdata = 55'b0000000000000000000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 63) begin
	always @(*) begin
		case(address)
			default : rdata = 55'b0000000000000000000000000000000000000000000000000000000;
		endcase
	end
end

endgenerate
endmodule