module accelerator#(
    parameter INPUT_BITWIDTH = `INPUT_BITWIDTH,
    parameter BITWIDTH = `BITWIDTH,
    parameter SIZE = `SIZE
)(
input clk,
input rst_n,
%input%
%output%
);
%logic%
%stage%

endmodule;
