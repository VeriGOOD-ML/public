`timescale 1ns/1ps
module sigmoid#(

)(
	in,
	out
);

	parameter dataLen = 32;
	parameter indexLen =9;
	parameter fracLen = 16;

	input signed [dataLen - 1 : 0] in;
	output reg [dataLen - 1 : 0] out;
	reg [indexLen - 1 :0] index;

	always @(in)
	begin
		out = 0;

		if (in < -(8 << 16) begin
			out = 0;
		end else if (in > (8 << 16)) begin
			out = 1<<16;
		end else begin
		index[indexLen-1]	= in[dataLen-1];
		index[indexLen-2:0]	= in[fracLen+indexLen-5:fracLen-5];
		case(index)
            //
            9'd0= 32'b00000000000000001000000000000000;
            9'd1= 32'b00000000000000001000000111111111;
            9'd2= 32'b00000000000000001000001111111111;
            9'd3= 32'b00000000000000001000010111111110;
            9'd4= 32'b00000000000000001000011111111101;
            9'd5= 32'b00000000000000001000100111111010;
            9'd6= 32'b00000000000000001000101111110111;
            9'd7= 32'b00000000000000001000110111110001;
            9'd8= 32'b00000000000000001000111111101010;
            9'd9= 32'b00000000000000001001000111100001;
            9'd10= 32'b00000000000000001001001111010110;
            9'd11= 32'b00000000000000001001010111001001;
            9'd12= 32'b00000000000000001001011110111000;
            9'd13= 32'b00000000000000001001100110100101;
            9'd14= 32'b00000000000000001001101110001111;
            9'd15= 32'b00000000000000001001110101110110;
            9'd16= 32'b00000000000000001001111101011001;
            9'd17= 32'b00000000000000001010000100111000;
            9'd18= 32'b00000000000000001010001100010100;
            9'd19= 32'b00000000000000001010010011101011;
            9'd20= 32'b00000000000000001010011010111111;
            9'd21= 32'b00000000000000001010100010001110;
            9'd22= 32'b00000000000000001010101001011000;
            9'd23= 32'b00000000000000001010110000011101;
            9'd24= 32'b00000000000000001010110111011110;
            9'd25= 32'b00000000000000001010111110011010;
            9'd26= 32'b00000000000000001011000101010000;
            9'd27= 32'b00000000000000001011001100000010;
            9'd28= 32'b00000000000000001011010010101110;
            9'd29= 32'b00000000000000001011011001010100;
            9'd30= 32'b00000000000000001011011111110101;
            9'd31= 32'b00000000000000001011100110010001;
            9'd32= 32'b00000000000000001011101100100110;
            9'd33= 32'b00000000000000001011110010110110;
            9'd34= 32'b00000000000000001011111001000000;
            9'd35= 32'b00000000000000001011111111000100;
            9'd36= 32'b00000000000000001100000101000010;
            9'd37= 32'b00000000000000001100001010111010;
            9'd38= 32'b00000000000000001100010000101011;
            9'd39= 32'b00000000000000001100010110010111;
            9'd40= 32'b00000000000000001100011011111101;
            9'd41= 32'b00000000000000001100100001011100;
            9'd42= 32'b00000000000000001100100110110101;
            9'd43= 32'b00000000000000001100101100001000;
            9'd44= 32'b00000000000000001100110001010101;
            9'd45= 32'b00000000000000001100110110011100;
            9'd46= 32'b00000000000000001100111011011101;
            9'd47= 32'b00000000000000001101000000011000;
            9'd48= 32'b00000000000000001101000101001100;
            9'd49= 32'b00000000000000001101001001111010;
            9'd50= 32'b00000000000000001101001110100011;
            9'd51= 32'b00000000000000001101010011000101;
            9'd52= 32'b00000000000000001101010111100010;
            9'd53= 32'b00000000000000001101011011111000;
            9'd54= 32'b00000000000000001101100000001001;
            9'd55= 32'b00000000000000001101100100010100;
            9'd56= 32'b00000000000000001101101000011001;
            9'd57= 32'b00000000000000001101101100011001;
            9'd58= 32'b00000000000000001101110000010010;
            9'd59= 32'b00000000000000001101110100000111;
            9'd60= 32'b00000000000000001101110111110110;
            9'd61= 32'b00000000000000001101111011011111;
            9'd62= 32'b00000000000000001101111111000011;
            9'd63= 32'b00000000000000001110000010100010;
            9'd64= 32'b00000000000000001110000101111011;
            9'd65= 32'b00000000000000001110001001010000;
            9'd66= 32'b00000000000000001110001100011111;
            9'd67= 32'b00000000000000001110001111101010;
            9'd68= 32'b00000000000000001110010010101111;
            9'd69= 32'b00000000000000001110010101110000;
            9'd70= 32'b00000000000000001110011000101100;
            9'd71= 32'b00000000000000001110011011100100;
            9'd72= 32'b00000000000000001110011110010111;
            9'd73= 32'b00000000000000001110100001000101;
            9'd74= 32'b00000000000000001110100011101111;
            9'd75= 32'b00000000000000001110100110010101;
            9'd76= 32'b00000000000000001110101000110110;
            9'd77= 32'b00000000000000001110101011010100;
            9'd78= 32'b00000000000000001110101101101101;
            9'd79= 32'b00000000000000001110110000000011;
            9'd80= 32'b00000000000000001110110010010100;
            9'd81= 32'b00000000000000001110110100100010;
            9'd82= 32'b00000000000000001110110110101100;
            9'd83= 32'b00000000000000001110111000110010;
            9'd84= 32'b00000000000000001110111010110101;
            9'd85= 32'b00000000000000001110111100110100;
            9'd86= 32'b00000000000000001110111110110000;
            9'd87= 32'b00000000000000001111000000101000;
            9'd88= 32'b00000000000000001111000010011110;
            9'd89= 32'b00000000000000001111000100010000;
            9'd90= 32'b00000000000000001111000101111111;
            9'd91= 32'b00000000000000001111000111101011;
            9'd92= 32'b00000000000000001111001001010100;
            9'd93= 32'b00000000000000001111001010111010;
            9'd94= 32'b00000000000000001111001100011101;
            9'd95= 32'b00000000000000001111001101111110;
            9'd96= 32'b00000000000000001111001111011011;
            9'd97= 32'b00000000000000001111010000110111;
            9'd98= 32'b00000000000000001111010010001111;
            9'd99= 32'b00000000000000001111010011100101;
            9'd100= 32'b00000000000000001111010100111001;
            9'd101= 32'b00000000000000001111010110001011;
            9'd102= 32'b00000000000000001111010111011010;
            9'd103= 32'b00000000000000001111011000100111;
            9'd104= 32'b00000000000000001111011001110001;
            9'd105= 32'b00000000000000001111011010111010;
            9'd106= 32'b00000000000000001111011100000000;
            9'd107= 32'b00000000000000001111011101000101;
            9'd108= 32'b00000000000000001111011110000111;
            9'd109= 32'b00000000000000001111011111001000;
            9'd110= 32'b00000000000000001111100000000110;
            9'd111= 32'b00000000000000001111100001000011;
            9'd112= 32'b00000000000000001111100001111110;
            9'd113= 32'b00000000000000001111100010111000;
            9'd114= 32'b00000000000000001111100011110000;
            9'd115= 32'b00000000000000001111100100100110;
            9'd116= 32'b00000000000000001111100101011010;
            9'd117= 32'b00000000000000001111100110001101;
            9'd118= 32'b00000000000000001111100110111111;
            9'd119= 32'b00000000000000001111100111101111;
            9'd120= 32'b00000000000000001111101000011110;
            9'd121= 32'b00000000000000001111101001001011;
            9'd122= 32'b00000000000000001111101001110111;
            9'd123= 32'b00000000000000001111101010100010;
            9'd124= 32'b00000000000000001111101011001011;
            9'd125= 32'b00000000000000001111101011110011;
            9'd126= 32'b00000000000000001111101100011010;
            9'd127= 32'b00000000000000001111101101000000;
            9'd128= 32'b00000000000000001111101101100101;
            9'd129= 32'b00000000000000001111101110001000;
            9'd130= 32'b00000000000000001111101110101011;
            9'd131= 32'b00000000000000001111101111001101;
            9'd132= 32'b00000000000000001111101111101101;
            9'd133= 32'b00000000000000001111110000001101;
            9'd134= 32'b00000000000000001111110000101011;
            9'd135= 32'b00000000000000001111110001001001;
            9'd136= 32'b00000000000000001111110001100110;
            9'd137= 32'b00000000000000001111110010000010;
            9'd138= 32'b00000000000000001111110010011101;
            9'd139= 32'b00000000000000001111110010110111;
            9'd140= 32'b00000000000000001111110011010001;
            9'd141= 32'b00000000000000001111110011101010;
            9'd142= 32'b00000000000000001111110100000010;
            9'd143= 32'b00000000000000001111110100011001;
            9'd144= 32'b00000000000000001111110100101111;
            9'd145= 32'b00000000000000001111110101000101;
            9'd146= 32'b00000000000000001111110101011011;
            9'd147= 32'b00000000000000001111110101101111;
            9'd148= 32'b00000000000000001111110110000011;
            9'd149= 32'b00000000000000001111110110010111;
            9'd150= 32'b00000000000000001111110110101001;
            9'd151= 32'b00000000000000001111110110111100;
            9'd152= 32'b00000000000000001111110111001101;
            9'd153= 32'b00000000000000001111110111011111;
            9'd154= 32'b00000000000000001111110111101111;
            9'd155= 32'b00000000000000001111110111111111;
            9'd156= 32'b00000000000000001111111000001111;
            9'd157= 32'b00000000000000001111111000011110;
            9'd158= 32'b00000000000000001111111000101101;
            9'd159= 32'b00000000000000001111111000111011;
            9'd160= 32'b00000000000000001111111001001001;
            9'd161= 32'b00000000000000001111111001010110;
            9'd162= 32'b00000000000000001111111001100011;
            9'd163= 32'b00000000000000001111111001110000;
            9'd164= 32'b00000000000000001111111001111100;
            9'd165= 32'b00000000000000001111111010001000;
            9'd166= 32'b00000000000000001111111010010011;
            9'd167= 32'b00000000000000001111111010011111;
            9'd168= 32'b00000000000000001111111010101001;
            9'd169= 32'b00000000000000001111111010110100;
            9'd170= 32'b00000000000000001111111010111110;
            9'd171= 32'b00000000000000001111111011001000;
            9'd172= 32'b00000000000000001111111011010001;
            9'd173= 32'b00000000000000001111111011011011;
            9'd174= 32'b00000000000000001111111011100100;
            9'd175= 32'b00000000000000001111111011101100;
            9'd176= 32'b00000000000000001111111011110101;
            9'd177= 32'b00000000000000001111111011111101;
            9'd178= 32'b00000000000000001111111100000101;
            9'd179= 32'b00000000000000001111111100001101;
            9'd180= 32'b00000000000000001111111100010100;
            9'd181= 32'b00000000000000001111111100011011;
            9'd182= 32'b00000000000000001111111100100010;
            9'd183= 32'b00000000000000001111111100101001;
            9'd184= 32'b00000000000000001111111100110000;
            9'd185= 32'b00000000000000001111111100110110;
            9'd186= 32'b00000000000000001111111100111100;
            9'd187= 32'b00000000000000001111111101000010;
            9'd188= 32'b00000000000000001111111101001000;
            9'd189= 32'b00000000000000001111111101001110;
            9'd190= 32'b00000000000000001111111101010011;
            9'd191= 32'b00000000000000001111111101011000;
            9'd192= 32'b00000000000000001111111101011101;
            9'd193= 32'b00000000000000001111111101100010;
            9'd194= 32'b00000000000000001111111101100111;
            9'd195= 32'b00000000000000001111111101101100;
            9'd196= 32'b00000000000000001111111101110000;
            9'd197= 32'b00000000000000001111111101110101;
            9'd198= 32'b00000000000000001111111101111001;
            9'd199= 32'b00000000000000001111111101111101;
            9'd200= 32'b00000000000000001111111110000001;
            9'd201= 32'b00000000000000001111111110000101;
            9'd202= 32'b00000000000000001111111110001001;
            9'd203= 32'b00000000000000001111111110001101;
            9'd204= 32'b00000000000000001111111110010000;
            9'd205= 32'b00000000000000001111111110010011;
            9'd206= 32'b00000000000000001111111110010111;
            9'd207= 32'b00000000000000001111111110011010;
            9'd208= 32'b00000000000000001111111110011101;
            9'd209= 32'b00000000000000001111111110100000;
            9'd210= 32'b00000000000000001111111110100011;
            9'd211= 32'b00000000000000001111111110100110;
            9'd212= 32'b00000000000000001111111110101001;
            9'd213= 32'b00000000000000001111111110101011;
            9'd214= 32'b00000000000000001111111110101110;
            9'd215= 32'b00000000000000001111111110110000;
            9'd216= 32'b00000000000000001111111110110011;
            9'd217= 32'b00000000000000001111111110110101;
            9'd218= 32'b00000000000000001111111110110111;
            9'd219= 32'b00000000000000001111111110111010;
            9'd220= 32'b00000000000000001111111110111100;
            9'd221= 32'b00000000000000001111111110111110;
            9'd222= 32'b00000000000000001111111111000000;
            9'd223= 32'b00000000000000001111111111000010;
            9'd224= 32'b00000000000000001111111111000100;
            9'd225= 32'b00000000000000001111111111000110;
            9'd226= 32'b00000000000000001111111111000111;
            9'd227= 32'b00000000000000001111111111001001;
            9'd228= 32'b00000000000000001111111111001011;
            9'd229= 32'b00000000000000001111111111001100;
            9'd230= 32'b00000000000000001111111111001110;
            9'd231= 32'b00000000000000001111111111010000;
            9'd232= 32'b00000000000000001111111111010001;
            9'd233= 32'b00000000000000001111111111010010;
            9'd234= 32'b00000000000000001111111111010100;
            9'd235= 32'b00000000000000001111111111010101;
            9'd236= 32'b00000000000000001111111111010110;
            9'd237= 32'b00000000000000001111111111011000;
            9'd238= 32'b00000000000000001111111111011001;
            9'd239= 32'b00000000000000001111111111011010;
            9'd240= 32'b00000000000000001111111111011011;
            9'd241= 32'b00000000000000001111111111011100;
            9'd242= 32'b00000000000000001111111111011101;
            9'd243= 32'b00000000000000001111111111011111;
            9'd244= 32'b00000000000000001111111111100000;
            9'd245= 32'b00000000000000001111111111100001;
            9'd246= 32'b00000000000000001111111111100001;
            9'd247= 32'b00000000000000001111111111100010;
            9'd248= 32'b00000000000000001111111111100011;
            9'd249= 32'b00000000000000001111111111100100;
            9'd250= 32'b00000000000000001111111111100101;
            9'd251= 32'b00000000000000001111111111100110;
            9'd252= 32'b00000000000000001111111111100111;
            9'd253= 32'b00000000000000001111111111100111;
            9'd254= 32'b00000000000000001111111111101000;
            9'd255= 32'b00000000000000001111111111101001;
            9'd256= 32'b00000000000000000000000000010101;
            9'd257= 32'b00000000000000000000000000010110;
            9'd258= 32'b00000000000000000000000000010111;
            9'd259= 32'b00000000000000000000000000011000;
            9'd260= 32'b00000000000000000000000000011000;
            9'd261= 32'b00000000000000000000000000011001;
            9'd262= 32'b00000000000000000000000000011010;
            9'd263= 32'b00000000000000000000000000011011;
            9'd264= 32'b00000000000000000000000000011100;
            9'd265= 32'b00000000000000000000000000011101;
            9'd266= 32'b00000000000000000000000000011110;
            9'd267= 32'b00000000000000000000000000011110;
            9'd268= 32'b00000000000000000000000000011111;
            9'd269= 32'b00000000000000000000000000100000;
            9'd270= 32'b00000000000000000000000000100010;
            9'd271= 32'b00000000000000000000000000100011;
            9'd272= 32'b00000000000000000000000000100100;
            9'd273= 32'b00000000000000000000000000100101;
            9'd274= 32'b00000000000000000000000000100110;
            9'd275= 32'b00000000000000000000000000100111;
            9'd276= 32'b00000000000000000000000000101001;
            9'd277= 32'b00000000000000000000000000101010;
            9'd278= 32'b00000000000000000000000000101011;
            9'd279= 32'b00000000000000000000000000101101;
            9'd280= 32'b00000000000000000000000000101110;
            9'd281= 32'b00000000000000000000000000101111;
            9'd282= 32'b00000000000000000000000000110001;
            9'd283= 32'b00000000000000000000000000110011;
            9'd284= 32'b00000000000000000000000000110100;
            9'd285= 32'b00000000000000000000000000110110;
            9'd286= 32'b00000000000000000000000000111000;
            9'd287= 32'b00000000000000000000000000111001;
            9'd288= 32'b00000000000000000000000000111011;
            9'd289= 32'b00000000000000000000000000111101;
            9'd290= 32'b00000000000000000000000000111111;
            9'd291= 32'b00000000000000000000000001000001;
            9'd292= 32'b00000000000000000000000001000011;
            9'd293= 32'b00000000000000000000000001000101;
            9'd294= 32'b00000000000000000000000001001000;
            9'd295= 32'b00000000000000000000000001001010;
            9'd296= 32'b00000000000000000000000001001100;
            9'd297= 32'b00000000000000000000000001001111;
            9'd298= 32'b00000000000000000000000001010001;
            9'd299= 32'b00000000000000000000000001010100;
            9'd300= 32'b00000000000000000000000001010110;
            9'd301= 32'b00000000000000000000000001011001;
            9'd302= 32'b00000000000000000000000001011100;
            9'd303= 32'b00000000000000000000000001011111;
            9'd304= 32'b00000000000000000000000001100010;
            9'd305= 32'b00000000000000000000000001100101;
            9'd306= 32'b00000000000000000000000001101000;
            9'd307= 32'b00000000000000000000000001101100;
            9'd308= 32'b00000000000000000000000001101111;
            9'd309= 32'b00000000000000000000000001110010;
            9'd310= 32'b00000000000000000000000001110110;
            9'd311= 32'b00000000000000000000000001111010;
            9'd312= 32'b00000000000000000000000001111110;
            9'd313= 32'b00000000000000000000000010000010;
            9'd314= 32'b00000000000000000000000010000110;
            9'd315= 32'b00000000000000000000000010001010;
            9'd316= 32'b00000000000000000000000010001111;
            9'd317= 32'b00000000000000000000000010010011;
            9'd318= 32'b00000000000000000000000010011000;
            9'd319= 32'b00000000000000000000000010011101;
            9'd320= 32'b00000000000000000000000010100010;
            9'd321= 32'b00000000000000000000000010100111;
            9'd322= 32'b00000000000000000000000010101100;
            9'd323= 32'b00000000000000000000000010110001;
            9'd324= 32'b00000000000000000000000010110111;
            9'd325= 32'b00000000000000000000000010111101;
            9'd326= 32'b00000000000000000000000011000011;
            9'd327= 32'b00000000000000000000000011001001;
            9'd328= 32'b00000000000000000000000011001111;
            9'd329= 32'b00000000000000000000000011010110;
            9'd330= 32'b00000000000000000000000011011101;
            9'd331= 32'b00000000000000000000000011100100;
            9'd332= 32'b00000000000000000000000011101011;
            9'd333= 32'b00000000000000000000000011110010;
            9'd334= 32'b00000000000000000000000011111010;
            9'd335= 32'b00000000000000000000000100000010;
            9'd336= 32'b00000000000000000000000100001010;
            9'd337= 32'b00000000000000000000000100010011;
            9'd338= 32'b00000000000000000000000100011011;
            9'd339= 32'b00000000000000000000000100100100;
            9'd340= 32'b00000000000000000000000100101110;
            9'd341= 32'b00000000000000000000000100110111;
            9'd342= 32'b00000000000000000000000101000001;
            9'd343= 32'b00000000000000000000000101001011;
            9'd344= 32'b00000000000000000000000101010110;
            9'd345= 32'b00000000000000000000000101100000;
            9'd346= 32'b00000000000000000000000101101100;
            9'd347= 32'b00000000000000000000000101110111;
            9'd348= 32'b00000000000000000000000110000011;
            9'd349= 32'b00000000000000000000000110001111;
            9'd350= 32'b00000000000000000000000110011100;
            9'd351= 32'b00000000000000000000000110101001;
            9'd352= 32'b00000000000000000000000110110110;
            9'd353= 32'b00000000000000000000000111000100;
            9'd354= 32'b00000000000000000000000111010010;
            9'd355= 32'b00000000000000000000000111100001;
            9'd356= 32'b00000000000000000000000111110000;
            9'd357= 32'b00000000000000000000001000000000;
            9'd358= 32'b00000000000000000000001000010000;
            9'd359= 32'b00000000000000000000001000100000;
            9'd360= 32'b00000000000000000000001000110010;
            9'd361= 32'b00000000000000000000001001000011;
            9'd362= 32'b00000000000000000000001001010110;
            9'd363= 32'b00000000000000000000001001101000;
            9'd364= 32'b00000000000000000000001001111100;
            9'd365= 32'b00000000000000000000001010010000;
            9'd366= 32'b00000000000000000000001010100100;
            9'd367= 32'b00000000000000000000001010111010;
            9'd368= 32'b00000000000000000000001011010000;
            9'd369= 32'b00000000000000000000001011100110;
            9'd370= 32'b00000000000000000000001011111101;
            9'd371= 32'b00000000000000000000001100010101;
            9'd372= 32'b00000000000000000000001100101110;
            9'd373= 32'b00000000000000000000001101001000;
            9'd374= 32'b00000000000000000000001101100010;
            9'd375= 32'b00000000000000000000001101111101;
            9'd376= 32'b00000000000000000000001110011001;
            9'd377= 32'b00000000000000000000001110110110;
            9'd378= 32'b00000000000000000000001111010100;
            9'd379= 32'b00000000000000000000001111110010;
            9'd380= 32'b00000000000000000000010000010010;
            9'd381= 32'b00000000000000000000010000110010;
            9'd382= 32'b00000000000000000000010001010100;
            9'd383= 32'b00000000000000000000010001110111;
            9'd384= 32'b00000000000000000000010010011010;
            9'd385= 32'b00000000000000000000010010111111;
            9'd386= 32'b00000000000000000000010011100101;
            9'd387= 32'b00000000000000000000010100001100;
            9'd388= 32'b00000000000000000000010100110100;
            9'd389= 32'b00000000000000000000010101011101;
            9'd390= 32'b00000000000000000000010110001000;
            9'd391= 32'b00000000000000000000010110110100;
            9'd392= 32'b00000000000000000000010111100001;
            9'd393= 32'b00000000000000000000011000010000;
            9'd394= 32'b00000000000000000000011001000000;
            9'd395= 32'b00000000000000000000011001110010;
            9'd396= 32'b00000000000000000000011010100101;
            9'd397= 32'b00000000000000000000011011011001;
            9'd398= 32'b00000000000000000000011100001111;
            9'd399= 32'b00000000000000000000011101000111;
            9'd400= 32'b00000000000000000000011110000001;
            9'd401= 32'b00000000000000000000011110111100;
            9'd402= 32'b00000000000000000000011111111001;
            9'd403= 32'b00000000000000000000100000110111;
            9'd404= 32'b00000000000000000000100001111000;
            9'd405= 32'b00000000000000000000100010111010;
            9'd406= 32'b00000000000000000000100011111111;
            9'd407= 32'b00000000000000000000100101000101;
            9'd408= 32'b00000000000000000000100110001110;
            9'd409= 32'b00000000000000000000100111011000;
            9'd410= 32'b00000000000000000000101000100101;
            9'd411= 32'b00000000000000000000101001110100;
            9'd412= 32'b00000000000000000000101011000110;
            9'd413= 32'b00000000000000000000101100011010;
            9'd414= 32'b00000000000000000000101101110000;
            9'd415= 32'b00000000000000000000101111001000;
            9'd416= 32'b00000000000000000000110000100100;
            9'd417= 32'b00000000000000000000110010000001;
            9'd418= 32'b00000000000000000000110011100010;
            9'd419= 32'b00000000000000000000110101000101;
            9'd420= 32'b00000000000000000000110110101011;
            9'd421= 32'b00000000000000000000111000010100;
            9'd422= 32'b00000000000000000000111010000000;
            9'd423= 32'b00000000000000000000111011101111;
            9'd424= 32'b00000000000000000000111101100001;
            9'd425= 32'b00000000000000000000111111010111;
            9'd426= 32'b00000000000000000001000001001111;
            9'd427= 32'b00000000000000000001000011001011;
            9'd428= 32'b00000000000000000001000101001010;
            9'd429= 32'b00000000000000000001000111001101;
            9'd430= 32'b00000000000000000001001001010011;
            9'd431= 32'b00000000000000000001001011011101;
            9'd432= 32'b00000000000000000001001101101011;
            9'd433= 32'b00000000000000000001001111111100;
            9'd434= 32'b00000000000000000001010010010010;
            9'd435= 32'b00000000000000000001010100101011;
            9'd436= 32'b00000000000000000001010111001001;
            9'd437= 32'b00000000000000000001011001101010;
            9'd438= 32'b00000000000000000001011100010000;
            9'd439= 32'b00000000000000000001011110111010;
            9'd440= 32'b00000000000000000001100001101000;
            9'd441= 32'b00000000000000000001100100011011;
            9'd442= 32'b00000000000000000001100111010011;
            9'd443= 32'b00000000000000000001101010001111;
            9'd444= 32'b00000000000000000001101101010000;
            9'd445= 32'b00000000000000000001110000010101;
            9'd446= 32'b00000000000000000001110011100000;
            9'd447= 32'b00000000000000000001110110101111;
            9'd448= 32'b00000000000000000001111010000100;
            9'd449= 32'b00000000000000000001111101011101;
            9'd450= 32'b00000000000000000010000000111100;
            9'd451= 32'b00000000000000000010000100100000;
            9'd452= 32'b00000000000000000010001000001001;
            9'd453= 32'b00000000000000000010001011111000;
            9'd454= 32'b00000000000000000010001111101101;
            9'd455= 32'b00000000000000000010010011100110;
            9'd456= 32'b00000000000000000010010111100110;
            9'd457= 32'b00000000000000000010011011101011;
            9'd458= 32'b00000000000000000010011111110110;
            9'd459= 32'b00000000000000000010100100000111;
            9'd460= 32'b00000000000000000010101000011101;
            9'd461= 32'b00000000000000000010101100111010;
            9'd462= 32'b00000000000000000010110001011100;
            9'd463= 32'b00000000000000000010110110000101;
            9'd464= 32'b00000000000000000010111010110011;
            9'd465= 32'b00000000000000000010111111100111;
            9'd466= 32'b00000000000000000011000100100010;
            9'd467= 32'b00000000000000000011001001100011;
            9'd468= 32'b00000000000000000011001110101010;
            9'd469= 32'b00000000000000000011010011110111;
            9'd470= 32'b00000000000000000011011001001010;
            9'd471= 32'b00000000000000000011011110100011;
            9'd472= 32'b00000000000000000011100100000010;
            9'd473= 32'b00000000000000000011101001101000;
            9'd474= 32'b00000000000000000011101111010100;
            9'd475= 32'b00000000000000000011110101000101;
            9'd476= 32'b00000000000000000011111010111101;
            9'd477= 32'b00000000000000000100000000111011;
            9'd478= 32'b00000000000000000100000110111111;
            9'd479= 32'b00000000000000000100001101001001;
            9'd480= 32'b00000000000000000100010011011001;
            9'd481= 32'b00000000000000000100011001101110;
            9'd482= 32'b00000000000000000100100000001010;
            9'd483= 32'b00000000000000000100100110101011;
            9'd484= 32'b00000000000000000100101101010001;
            9'd485= 32'b00000000000000000100110011111101;
            9'd486= 32'b00000000000000000100111010101111;
            9'd487= 32'b00000000000000000101000001100101;
            9'd488= 32'b00000000000000000101001000100001;
            9'd489= 32'b00000000000000000101001111100010;
            9'd490= 32'b00000000000000000101010110100111;
            9'd491= 32'b00000000000000000101011101110001;
            9'd492= 32'b00000000000000000101100101000000;
            9'd493= 32'b00000000000000000101101100010100;
            9'd494= 32'b00000000000000000101110011101011;
            9'd495= 32'b00000000000000000101111011000111;
            9'd496= 32'b00000000000000000110000010100110;
            9'd497= 32'b00000000000000000110001010001001;
            9'd498= 32'b00000000000000000110010001110000;
            9'd499= 32'b00000000000000000110011001011010;
            9'd500= 32'b00000000000000000110100001000111;
            9'd501= 32'b00000000000000000110101000110110;
            9'd502= 32'b00000000000000000110110000101001;
            9'd503= 32'b00000000000000000110111000011110;
            9'd504= 32'b00000000000000000111000000010101;
            9'd505= 32'b00000000000000000111001000001110;
            9'd506= 32'b00000000000000000111010000001000;
            9'd507= 32'b00000000000000000111011000000101;
            9'd508= 32'b00000000000000000111100000000010;
            9'd509= 32'b00000000000000000111101000000001;
            9'd510= 32'b00000000000000000111110000000000;
            9'd511= 32'b00000000000000000111111000000000;
		endcase
		end
	end

endmodule
  