
`timescale 1ns/1ps
module instruction_memory #(
    parameter integer addrLen = 5,
    parameter integer dataLen = 32,
    parameter integer peId  = 1
)(
    input clk,
    input rstn,
    
    input stall,
    input start,
    input restart,
    
    output reg [dataLen - 1: 0] data_out
);
//--------------------------------------------------------------------------------------
//reg [dataLen - 1: 0] mem  [0: (1 << addrLen) - 1];
reg [addrLen-1:0]        address;
reg enable;
reg [dataLen - 1: 0] rdata;
wire end_of_instruction;
always @(posedge clk or negedge rstn)
    if(~rstn)
        enable <= 1'b0;
    else if(start)
        enable <= 1'b1;
    else if(end_of_instruction)
       enable <= 1'b0;
always @(posedge clk or negedge rstn) begin
    if(~rstn)
        address <= {addrLen{1'b0}};
    else begin
        if(end_of_instruction)
            address <= {addrLen{1'b0}};
        else if(~stall && enable )
            address <= address + {{addrLen-1{1'b0}},1'b1};   
    end     
end
always @(posedge clk or negedge rstn) begin
    if(~rstn)
        data_out <= {1'b1,{dataLen-1{1'b0}}};
    else if((~stall && enable && ~end_of_instruction)||(end_of_instruction && start))
       data_out <= rdata;
end
    
assign end_of_instruction = (data_out[dataLen-1:dataLen-5] == 5'b0);
/****************************************************************************/
generate
if(peId == 0) begin
	always @(*) begin
		case(address)
			// PEs: 7 -> 8
			// srcs: (3, 0)(122) 0 --> (122) 0:PENB, pass, PUNB
			6'd0 : rdata = 41'b11000110111111100000000000000001000000000;
			// PEs: 6 -> 16
			// srcs: (9, 1)(173) -4 --> (173) -4:PEGB6, pass, PUGB2
			6'd1 : rdata = 41'b11000111000011000000000000000000000001010;
			// PEs: 1 -> 40
			// srcs: (17, 2)(172) -6 --> (172) -6:PEGB1, pass, PUGB5
			6'd2 : rdata = 41'b11000111000000100000000000000000000001101;
			// PEs: 8 -> 0
			// srcs: (25, 3)(178) -4 --> (178) -4:PUGB1, pass, NI0
			6'd3 : rdata = 41'b11000111000000110000000000010000000000000;
			// PEs: 32 -> 1
			// srcs: (33, 4)(180) 2 --> (180) 2:PUGB4, pass, PENB
			6'd4 : rdata = 41'b11000111000010010000000000000000100000000;
			// PEs: 0 -> 1
			// srcs: (40, 5)(178) -4 --> (178) -4:NI0, pass, PENB
			6'd5 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 48 -> 0
			// srcs: (46, 7)(202) 9 --> (202) 9:PUGB6, pass, NI0
			6'd6 : rdata = 41'b11000111000011010000000000010000000000000;
			// PEs: 1 -> 40
			// srcs: (47, 6)(181) -2 --> (181) -2:PEGB1, pass, PUGB5
			6'd7 : rdata = 41'b11000111000000100000000000000000000001101;
			// PEs: 8 -> 1
			// srcs: (50, 8)(208) -3 --> (208) -3:PUGB1, pass, PENB
			6'd8 : rdata = 41'b11000111000000110000000000000000100000000;
			// PEs: 0 -> 1
			// srcs: (57, 9)(202) 9 --> (202) 9:NI0, pass, PENB
			6'd9 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 1 -> 8
			// srcs: (64, 10)(209) 6 --> (209) 6:PEGB1, pass, PUNB
			6'd10 : rdata = 41'b11000111000000100000000000000001000000000;
			// PEs: 48 -> 1
			// srcs: (101, 11)(224) 3 --> (224) 3:PUGB6, pass, PENB
			6'd11 : rdata = 41'b11000111000011010000000000000000100000000;
			// PEs: 48 -> 2
			// srcs: (105, 12)(224) 3 --> (224) 3:PUGB6, pass, PEGB2
			6'd12 : rdata = 41'b11000111000011010000000000000000010100000;
			// PEs: 48 -> 3
			// srcs: (106, 13)(224) 3 --> (224) 3:PUGB6, pass, PEGB3
			6'd13 : rdata = 41'b11000111000011010000000000000000010110000;
			// PEs: 48 -> 4
			// srcs: (107, 14)(224) 3 --> (224) 3:PUGB6, pass, PEGB4
			6'd14 : rdata = 41'b11000111000011010000000000000000011000000;
			// PEs: 48 -> 5
			// srcs: (108, 15)(224) 3 --> (224) 3:PUGB6, pass, PEGB5
			6'd15 : rdata = 41'b11000111000011010000000000000000011010000;
			// PEs: 48 -> 6
			// srcs: (109, 16)(224) 3 --> (224) 3:PUGB6, pass, PEGB6
			6'd16 : rdata = 41'b11000111000011010000000000000000011100000;
			// PEs: 48 -> 7
			// srcs: (111, 17)(224) 3 --> (224) 3:PUGB6, pass, PEGB7
			6'd17 : rdata = 41'b11000111000011010000000000000000011110000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 1) begin
	always @(*) begin
		case(address)
			// PEs: 1, 1 -> 2
			// srcs: (1, 0)(4) 2, (60) -2 --> (115) -4:ND0, NW0, *, PENB
			6'd0 : rdata = 41'b00011011000000000100000000000000100000000;
			// PEs: 4 -> 
			// srcs: (9, 1)(171) 0 --> (171) 0:PEGB4, pass, 
			6'd1 : rdata = 41'b11000111000010000000000000000000000000000;
			// PEs: 2, 1 -> 0
			// srcs: (12, 2)(170) -6, (171) 0 --> (172) -6:PEGB2, ALU, +, PEGB0
			6'd2 : rdata = 41'b00001111000001000011111111100000010000000;
			// PEs: 0 -> 
			// srcs: (35, 3)(180) 2 --> (180) 2:PENB, pass, 
			6'd3 : rdata = 41'b11000110111111100000000000000000000000000;
			// PEs: 0, 1 -> 0
			// srcs: (42, 4)(178) -4, (180) 2 --> (181) -2:PENB, ALU, +, PEGB0
			6'd4 : rdata = 41'b00001110111111100011111111100000010000000;
			// PEs: 0 -> 
			// srcs: (52, 5)(208) -3 --> (208) -3:PENB, pass, 
			6'd5 : rdata = 41'b11000110111111100000000000000000000000000;
			// PEs: 0, 1 -> 0
			// srcs: (59, 6)(202) 9, (208) -3 --> (209) 6:PENB, ALU, +, PEGB0
			6'd6 : rdata = 41'b00001110111111100011111111100000010000000;
			// PEs: 0, 1 -> 2
			// srcs: (104, 7)(224) 3, (4) 2 --> (225) 6:PENB, ND0, *, PENB
			6'd7 : rdata = 41'b00011110111111100110000000000000100000000;
			// PEs: 1, 2 -> 1
			// srcs: (113, 8)(60) -2, (280) 6 --> (335) -8:NW0, PEGB2, -, NW0
			6'd8 : rdata = 41'b00010010000000001110000010000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 2) begin
	always @(*) begin
		case(address)
			// PEs: 2, 2 -> 
			// srcs: (1, 0)(5) 2, (61) -1 --> (116) -2:ND0, NW0, *, 
			6'd0 : rdata = 41'b00011011000000000100000000000000000000000;
			// PEs: 1, 2 -> 1
			// srcs: (4, 1)(115) -4, (116) -2 --> (170) -6:PENB, ALU, +, PEGB1
			6'd1 : rdata = 41'b00001110111111100011111111100000010010000;
			// PEs: 2, 1 -> 1
			// srcs: (107, 3)(3) 1, (225) 6 --> (280) 6:NM0, PENB, *, PEGB1
			6'd2 : rdata = 41'b00011100000000001101111111000000010010000;
			// PEs: 0, 2 -> 3
			// srcs: (110, 2)(224) 3, (5) 2 --> (226) 6:PEGB0, ND0, *, PENB
			6'd3 : rdata = 41'b00011111000000000110000000000000100000000;
			// PEs: 2, 3 -> 2
			// srcs: (119, 4)(61) -1, (281) 6 --> (336) -7:NW0, PEGB3, -, NW0
			6'd4 : rdata = 41'b00010010000000001110000011000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 3) begin
	always @(*) begin
		case(address)
			// PEs: 3, 3 -> 4
			// srcs: (1, 0)(6) -1, (62) 0 --> (117) 0:ND0, NW0, *, PENB
			6'd0 : rdata = 41'b00011011000000000100000000000000100000000;
			// PEs: 0, 3 -> 3
			// srcs: (111, 1)(224) 3, (6) -1 --> (227) -3:PEGB0, ND0, *, NI0
			6'd1 : rdata = 41'b00011111000000000110000000010000000000000;
			// PEs: 3, 2 -> 2
			// srcs: (113, 2)(3) 1, (226) 6 --> (281) 6:NM0, PENB, *, PEGB2
			6'd2 : rdata = 41'b00011100000000001101111111000000010100000;
			// PEs: 3, 3 -> 
			// srcs: (114, 3)(3) 1, (227) -3 --> (282) -3:NM0, NI0, *, 
			6'd3 : rdata = 41'b00011100000000001010000000000000000000000;
			// PEs: 3, 3 -> 3
			// srcs: (117, 4)(62) 0, (282) -3 --> (337) 3:NW0, ALU, -, NW0
			6'd4 : rdata = 41'b00010010000000000011111111100100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 4) begin
	always @(*) begin
		case(address)
			// PEs: 4, 4 -> 
			// srcs: (1, 0)(7) -1, (63) 0 --> (118) 0:ND0, NW0, *, 
			6'd0 : rdata = 41'b00011011000000000100000000000000000000000;
			// PEs: 3, 4 -> 1
			// srcs: (4, 1)(117) 0, (118) 0 --> (171) 0:PENB, ALU, +, PEGB1
			6'd1 : rdata = 41'b00001110111111100011111111100000010010000;
			// PEs: 0, 4 -> 5
			// srcs: (112, 2)(224) 3, (7) -1 --> (228) -3:PEGB0, ND0, *, PENB
			6'd2 : rdata = 41'b00011111000000000110000000000000100000000;
			// PEs: 4, 5 -> 4
			// srcs: (121, 3)(63) 0, (283) -3 --> (338) 3:NW0, PEGB5, -, NW0
			6'd3 : rdata = 41'b00010010000000001110000101000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 5) begin
	always @(*) begin
		case(address)
			// PEs: 5, 5 -> 6
			// srcs: (1, 0)(8) -1, (64) 0 --> (119) 0:ND0, NW0, *, PENB
			6'd0 : rdata = 41'b00011011000000000100000000000000100000000;
			// PEs: 0, 5 -> 5
			// srcs: (113, 1)(224) 3, (8) -1 --> (229) -3:PEGB0, ND0, *, NI0
			6'd1 : rdata = 41'b00011111000000000110000000010000000000000;
			// PEs: 5, 4 -> 4
			// srcs: (115, 2)(3) 1, (228) -3 --> (283) -3:NM0, PENB, *, PEGB4
			6'd2 : rdata = 41'b00011100000000001101111111000000011000000;
			// PEs: 5, 5 -> 
			// srcs: (116, 3)(3) 1, (229) -3 --> (284) -3:NM0, NI0, *, 
			6'd3 : rdata = 41'b00011100000000001010000000000000000000000;
			// PEs: 5, 5 -> 5
			// srcs: (119, 4)(64) 0, (284) -3 --> (339) 3:NW0, ALU, -, NW0
			6'd4 : rdata = 41'b00010010000000000011111111100100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 6) begin
	always @(*) begin
		case(address)
			// PEs: 6, 6 -> 
			// srcs: (1, 0)(9) -2, (65) 2 --> (120) -4:ND0, NW0, *, 
			6'd0 : rdata = 41'b00011011000000000100000000000000000000000;
			// PEs: 5, 6 -> 0
			// srcs: (4, 1)(119) 0, (120) -4 --> (173) -4:PENB, ALU, +, PEGB0
			6'd1 : rdata = 41'b00001110111111100011111111100000010000000;
			// PEs: 0, 6 -> 7
			// srcs: (114, 2)(224) 3, (9) -2 --> (230) -6:PEGB0, ND0, *, PENB
			6'd2 : rdata = 41'b00011111000000000110000000000000100000000;
			// PEs: 6, 7 -> 6
			// srcs: (123, 3)(65) 2, (285) -6 --> (340) 8:NW0, PEGB7, -, NW0
			6'd3 : rdata = 41'b00010010000000001110000111000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 7) begin
	always @(*) begin
		case(address)
			// PEs: 7, 7 -> 0
			// srcs: (1, 0)(11) -1, (67) 0 --> (122) 0:ND0, NW0, *, PENB
			6'd0 : rdata = 41'b00011011000000000100000000000000100000000;
			// PEs: 0, 7 -> 7
			// srcs: (116, 1)(224) 3, (11) -1 --> (232) -3:PEGB0, ND0, *, NI0
			6'd1 : rdata = 41'b00011111000000000110000000010000000000000;
			// PEs: 7, 6 -> 6
			// srcs: (117, 2)(3) 1, (230) -6 --> (285) -6:NM0, PENB, *, PEGB6
			6'd2 : rdata = 41'b00011100000000001101111111000000011100000;
			// PEs: 7, 7 -> 
			// srcs: (119, 3)(3) 1, (232) -3 --> (287) -3:NM0, NI0, *, 
			6'd3 : rdata = 41'b00011100000000001010000000000000000000000;
			// PEs: 7, 7 -> 7
			// srcs: (122, 4)(67) 0, (287) -3 --> (342) 3:NW0, ALU, -, NW0
			6'd4 : rdata = 41'b00010010000000000011111111100100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 8) begin
	always @(*) begin
		case(address)
			// PEs: 0 -> 9
			// srcs: (5, 0)(122) 0 --> (122) 0:PUNB, pass, PENB
			6'd0 : rdata = 41'b11000110111111110000000000000000100000000;
			// PEs: 15 -> 16
			// srcs: (6, 2)(183) -6 --> (183) -6:PENB, pass, PUNB
			6'd1 : rdata = 41'b11000110111111100000000000000001000000000;
			// PEs: 13 -> 32
			// srcs: (9, 1)(179) 0 --> (179) 0:PEGB5, pass, PUGB4
			6'd2 : rdata = 41'b11000111000010100000000000000000000001100;
			// PEs: 40 -> 8
			// srcs: (18, 3)(206) 1 --> (206) 1:PUGB5, pass, NI0
			6'd3 : rdata = 41'b11000111000010110000000000010000000000000;
			// PEs: 56 -> 9
			// srcs: (19, 4)(156) 0 --> (156) 0:PUGB7, pass, PENB
			6'd4 : rdata = 41'b11000111000011110000000000000000100000000;
			// PEs: 10 -> 0
			// srcs: (20, 6)(178) -4 --> (178) -4:PEGB2, pass, PUGB0
			6'd5 : rdata = 41'b11000111000001000000000000000000000001000;
			// PEs: 8 -> 9
			// srcs: (25, 5)(206) 1 --> (206) 1:NI0, pass, PENB
			6'd6 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 32 -> 9
			// srcs: (26, 7)(205) -4 --> (205) -4:PUGB4, pass, PENB
			6'd7 : rdata = 41'b11000111000010010000000000000000100000000;
			// PEs: 9 -> 0
			// srcs: (45, 8)(208) -3 --> (208) -3:PEGB1, pass, PUGB0
			6'd8 : rdata = 41'b11000111000000100000000000000000000001000;
			// PEs: 16 -> 8
			// srcs: (48, 9)(215) 4 --> (215) 4:PUGB2, pass, NI0
			6'd9 : rdata = 41'b11000111000001010000000000010000000000000;
			// PEs: 56 -> 9
			// srcs: (49, 10)(220) 13 --> (220) 13:PUGB7, pass, PENB
			6'd10 : rdata = 41'b11000111000011110000000000000000100000000;
			// PEs: 8 -> 9
			// srcs: (55, 11)(215) 4 --> (215) 4:NI0, pass, PENB
			6'd11 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 0 -> 9
			// srcs: (66, 12)(209) 6 --> (209) 6:PUNB, pass, PENB
			6'd12 : rdata = 41'b11000110111111110000000000000000100000000;
			// PEs: 9 -> 48
			// srcs: (74, 13)(222) 23 --> (222) 23:PEGB1, pass, PUGB6
			6'd13 : rdata = 41'b11000111000000100000000000000000000001110;
			// PEs: 48 -> 9
			// srcs: (112, 14)(224) 3 --> (224) 3:PUGB6, pass, PENB
			6'd14 : rdata = 41'b11000111000011010000000000000000100000000;
			// PEs: 48 -> 10
			// srcs: (113, 15)(224) 3 --> (224) 3:PUGB6, pass, PEGB2
			6'd15 : rdata = 41'b11000111000011010000000000000000010100000;
			// PEs: 48 -> 11
			// srcs: (114, 16)(224) 3 --> (224) 3:PUGB6, pass, PEGB3
			6'd16 : rdata = 41'b11000111000011010000000000000000010110000;
			// PEs: 48 -> 12
			// srcs: (115, 17)(224) 3 --> (224) 3:PUGB6, pass, PEGB4
			6'd17 : rdata = 41'b11000111000011010000000000000000011000000;
			// PEs: 48 -> 13
			// srcs: (116, 18)(224) 3 --> (224) 3:PUGB6, pass, PEGB5
			6'd18 : rdata = 41'b11000111000011010000000000000000011010000;
			// PEs: 48 -> 14
			// srcs: (118, 19)(224) 3 --> (224) 3:PUGB6, pass, PEGB6
			6'd19 : rdata = 41'b11000111000011010000000000000000011100000;
			// PEs: 48 -> 15
			// srcs: (119, 20)(224) 3 --> (224) 3:PUGB6, pass, PEGB7
			6'd20 : rdata = 41'b11000111000011010000000000000000011110000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 9) begin
	always @(*) begin
		case(address)
			// PEs: 9, 9 -> 
			// srcs: (1, 0)(12) 1, (68) 2 --> (123) 2:ND0, NW0, *, 
			6'd0 : rdata = 41'b00011011000000000100000000000000000000000;
			// PEs: 8, 9 -> 10
			// srcs: (8, 1)(122) 0, (123) 2 --> (176) 2:PENB, ALU, +, PENB
			6'd1 : rdata = 41'b00001110111111100011111111100000100000000;
			// PEs: 8 -> 
			// srcs: (21, 2)(156) 0 --> (156) 0:PENB, pass, 
			6'd2 : rdata = 41'b11000110111111100000000000000000000000000;
			// PEs: 8, 9 -> 
			// srcs: (27, 3)(206) 1, (156) 0 --> (207) 1:PENB, ALU, +, 
			6'd3 : rdata = 41'b00001110111111100011111111100000000000000;
			// PEs: 8, 9 -> 8
			// srcs: (40, 4)(205) -4, (207) 1 --> (208) -3:PENB, ALU, +, PEGB0
			6'd4 : rdata = 41'b00001110111111100011111111100000010000000;
			// PEs: 8 -> 
			// srcs: (51, 5)(220) 13 --> (220) 13:PENB, pass, 
			6'd5 : rdata = 41'b11000110111111100000000000000000000000000;
			// PEs: 8, 9 -> 
			// srcs: (57, 6)(215) 4, (220) 13 --> (221) 17:PENB, ALU, +, 
			6'd6 : rdata = 41'b00001110111111100011111111100000000000000;
			// PEs: 8, 9 -> 8
			// srcs: (69, 7)(209) 6, (221) 17 --> (222) 23:PENB, ALU, +, PEGB0
			6'd7 : rdata = 41'b00001110111111100011111111100000010000000;
			// PEs: 8, 9 -> 10
			// srcs: (114, 8)(224) 3, (12) 1 --> (233) 3:PENB, ND0, *, PENB
			6'd8 : rdata = 41'b00011110111111100110000000000000100000000;
			// PEs: 9, 10 -> 9
			// srcs: (123, 9)(68) 2, (288) 3 --> (343) -1:NW0, PEGB2, -, NW0
			6'd9 : rdata = 41'b00010010000000001110000010000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 10) begin
	always @(*) begin
		case(address)
			// PEs: 10, 10 -> 11
			// srcs: (1, 0)(13) 0, (69) -1 --> (124) 0:ND0, NW0, *, PENB
			6'd0 : rdata = 41'b00011011000000000100000000000000100000000;
			// PEs: 9, 11 -> 8
			// srcs: (14, 1)(176) 2, (177) -6 --> (178) -4:PENB, PEGB3, +, PEGB0
			6'd1 : rdata = 41'b00001110111111101110000011000000010000000;
			// PEs: 10, 9 -> 9
			// srcs: (117, 3)(3) 1, (233) 3 --> (288) 3:NM0, PENB, *, PEGB1
			6'd2 : rdata = 41'b00011100000000001101111111000000010010000;
			// PEs: 8, 10 -> 11
			// srcs: (118, 2)(224) 3, (13) 0 --> (234) 0:PEGB0, ND0, *, PENB
			6'd3 : rdata = 41'b00011111000000000110000000000000100000000;
			// PEs: 10, 11 -> 10
			// srcs: (127, 4)(69) -1, (289) 0 --> (344) -1:NW0, PEGB3, -, NW0
			6'd4 : rdata = 41'b00010010000000001110000011000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 11) begin
	always @(*) begin
		case(address)
			// PEs: 11, 11 -> 
			// srcs: (1, 0)(14) -3, (70) 2 --> (125) -6:ND0, NW0, *, 
			6'd0 : rdata = 41'b00011011000000000100000000000000000000000;
			// PEs: 10, 11 -> 10
			// srcs: (4, 1)(124) 0, (125) -6 --> (177) -6:PENB, ALU, +, PEGB2
			6'd1 : rdata = 41'b00001110111111100011111111100000010100000;
			// PEs: 8, 11 -> 12
			// srcs: (119, 2)(224) 3, (14) -3 --> (235) -9:PEGB0, ND0, *, PENB
			6'd2 : rdata = 41'b00011111000000000110000000000000100000000;
			// PEs: 11, 10 -> 10
			// srcs: (121, 3)(3) 1, (234) 0 --> (289) 0:NM0, PENB, *, PEGB2
			6'd3 : rdata = 41'b00011100000000001101111111000000010100000;
			// PEs: 11, 12 -> 11
			// srcs: (128, 4)(70) 2, (290) -9 --> (345) 11:NW0, PEGB4, -, NW0
			6'd4 : rdata = 41'b00010010000000001110000100000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 12) begin
	always @(*) begin
		case(address)
			// PEs: 12, 12 -> 13
			// srcs: (1, 0)(15) 0, (71) 1 --> (126) 0:ND0, NW0, *, PENB
			6'd0 : rdata = 41'b00011011000000000100000000000000100000000;
			// PEs: 8, 12 -> 12
			// srcs: (120, 1)(224) 3, (15) 0 --> (236) 0:PEGB0, ND0, *, NI0
			6'd1 : rdata = 41'b00011111000000000110000000010000000000000;
			// PEs: 12, 11 -> 11
			// srcs: (122, 2)(3) 1, (235) -9 --> (290) -9:NM0, PENB, *, PEGB3
			6'd2 : rdata = 41'b00011100000000001101111111000000010110000;
			// PEs: 12, 12 -> 
			// srcs: (123, 3)(3) 1, (236) 0 --> (291) 0:NM0, NI0, *, 
			6'd3 : rdata = 41'b00011100000000001010000000000000000000000;
			// PEs: 12, 12 -> 12
			// srcs: (126, 4)(71) 1, (291) 0 --> (346) 1:NW0, ALU, -, NW0
			6'd4 : rdata = 41'b00010010000000000011111111100100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 13) begin
	always @(*) begin
		case(address)
			// PEs: 13, 13 -> 
			// srcs: (1, 0)(16) 1, (72) 0 --> (127) 0:ND0, NW0, *, 
			6'd0 : rdata = 41'b00011011000000000100000000000000000000000;
			// PEs: 12, 13 -> 8
			// srcs: (4, 1)(126) 0, (127) 0 --> (179) 0:PENB, ALU, +, PEGB0
			6'd1 : rdata = 41'b00001110111111100011111111100000010000000;
			// PEs: 8, 13 -> 14
			// srcs: (121, 2)(224) 3, (16) 1 --> (237) 3:PEGB0, ND0, *, PENB
			6'd2 : rdata = 41'b00011111000000000110000000000000100000000;
			// PEs: 13, 14 -> 13
			// srcs: (130, 3)(72) 0, (292) 3 --> (347) -3:NW0, PEGB6, -, NW0
			6'd3 : rdata = 41'b00010010000000001110000110000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 14) begin
	always @(*) begin
		case(address)
			// PEs: 14, 14 -> 15
			// srcs: (1, 0)(18) 0, (74) 1 --> (129) 0:ND0, NW0, *, PENB
			6'd0 : rdata = 41'b00011011000000000100000000000000100000000;
			// PEs: 8, 14 -> 14
			// srcs: (123, 1)(224) 3, (18) 0 --> (239) 0:PEGB0, ND0, *, NI0
			6'd1 : rdata = 41'b00011111000000000110000000010000000000000;
			// PEs: 14, 13 -> 13
			// srcs: (124, 2)(3) 1, (237) 3 --> (292) 3:NM0, PENB, *, PEGB5
			6'd2 : rdata = 41'b00011100000000001101111111000000011010000;
			// PEs: 14, 14 -> 
			// srcs: (126, 3)(3) 1, (239) 0 --> (294) 0:NM0, NI0, *, 
			6'd3 : rdata = 41'b00011100000000001010000000000000000000000;
			// PEs: 14, 14 -> 14
			// srcs: (129, 4)(74) 1, (294) 0 --> (349) 1:NW0, ALU, -, NW0
			6'd4 : rdata = 41'b00010010000000000011111111100100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 15) begin
	always @(*) begin
		case(address)
			// PEs: 15, 15 -> 
			// srcs: (1, 0)(19) 2, (75) -3 --> (130) -6:ND0, NW0, *, 
			6'd0 : rdata = 41'b00011011000000000100000000000000000000000;
			// PEs: 14, 15 -> 8
			// srcs: (4, 1)(129) 0, (130) -6 --> (183) -6:PENB, ALU, +, PENB
			6'd1 : rdata = 41'b00001110111111100011111111100000100000000;
			// PEs: 8, 15 -> 
			// srcs: (124, 2)(224) 3, (19) 2 --> (240) 6:PEGB0, ND0, *, 
			6'd2 : rdata = 41'b00011111000000000110000000000000000000000;
			// PEs: 15, 15 -> 
			// srcs: (127, 3)(3) 1, (240) 6 --> (295) 6:NM0, ALU, *, 
			6'd3 : rdata = 41'b00011100000000000011111111100000000000000;
			// PEs: 15, 15 -> 15
			// srcs: (130, 4)(75) -3, (295) 6 --> (350) -9:NW0, ALU, -, NW0
			6'd4 : rdata = 41'b00010010000000000011111111100100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 16) begin
	always @(*) begin
		case(address)
			// PEs: 23 -> 24
			// srcs: (3, 0)(138) 0 --> (138) 0:PENB, pass, PUNB
			6'd0 : rdata = 41'b11000110111111100000000000000001000000000;
			// PEs: 20 -> 24
			// srcs: (9, 5)(186) 0 --> (186) 0:PEGB4, pass, PUNB
			6'd1 : rdata = 41'b11000111000010000000000000000001000000000;
			// PEs: 22 -> 24
			// srcs: (10, 6)(189) 3 --> (189) 3:PEGB6, pass, PUNB
			6'd2 : rdata = 41'b11000111000011000000000000000001000000000;
			// PEs: 48 -> 16
			// srcs: (11, 2)(121) 1 --> (121) 1:PUGB6, pass, NI0
			6'd3 : rdata = 41'b11000111000011010000000000010000000000000;
			// PEs: 0 -> 17
			// srcs: (14, 1)(173) -4 --> (173) -4:PUGB0, pass, PENB
			6'd4 : rdata = 41'b11000111000000010000000000000000100000000;
			// PEs: 16 -> 17
			// srcs: (21, 3)(121) 1 --> (121) 1:NI0, pass, PENB
			6'd5 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 8 -> 17
			// srcs: (22, 4)(183) -6 --> (183) -6:PUNB, pass, PENB
			6'd6 : rdata = 41'b11000110111111110000000000000000100000000;
			// PEs: 40 -> 16
			// srcs: (23, 9)(212) -1 --> (212) -1:PUGB5, pass, NI0
			6'd7 : rdata = 41'b11000111000010110000000000010000000000000;
			// PEs: 17 -> 40
			// srcs: (28, 7)(174) -3 --> (174) -3:PEGB1, pass, PUGB5
			6'd8 : rdata = 41'b11000111000000100000000000000000000001101;
			// PEs: 17 -> 24
			// srcs: (29, 8)(185) -8 --> (185) -8:PEGB1, pass, PUNB
			6'd9 : rdata = 41'b11000111000000100000000000000001000000000;
			// PEs: 56 -> 17
			// srcs: (30, 10)(214) 5 --> (214) 5:PUGB7, pass, PENB
			6'd10 : rdata = 41'b11000111000011110000000000000000100000000;
			// PEs: 16 -> 17
			// srcs: (36, 11)(212) -1 --> (212) -1:NI0, pass, PENB
			6'd11 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 17 -> 8
			// srcs: (43, 12)(215) 4 --> (215) 4:PEGB1, pass, PUGB1
			6'd12 : rdata = 41'b11000111000000100000000000000000000001001;
			// PEs: 48 -> 17
			// srcs: (120, 13)(224) 3 --> (224) 3:PUGB6, pass, PENB
			6'd13 : rdata = 41'b11000111000011010000000000000000100000000;
			// PEs: 48 -> 18
			// srcs: (121, 14)(224) 3 --> (224) 3:PUGB6, pass, PEGB2
			6'd14 : rdata = 41'b11000111000011010000000000000000010100000;
			// PEs: 48 -> 19
			// srcs: (122, 15)(224) 3 --> (224) 3:PUGB6, pass, PEGB3
			6'd15 : rdata = 41'b11000111000011010000000000000000010110000;
			// PEs: 48 -> 20
			// srcs: (123, 16)(224) 3 --> (224) 3:PUGB6, pass, PEGB4
			6'd16 : rdata = 41'b11000111000011010000000000000000011000000;
			// PEs: 48 -> 21
			// srcs: (125, 17)(224) 3 --> (224) 3:PUGB6, pass, PEGB5
			6'd17 : rdata = 41'b11000111000011010000000000000000011010000;
			// PEs: 48 -> 22
			// srcs: (126, 18)(224) 3 --> (224) 3:PUGB6, pass, PEGB6
			6'd18 : rdata = 41'b11000111000011010000000000000000011100000;
			// PEs: 48 -> 23
			// srcs: (127, 19)(224) 3 --> (224) 3:PUGB6, pass, PEGB7
			6'd19 : rdata = 41'b11000111000011010000000000000000011110000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 17) begin
	always @(*) begin
		case(address)
			// PEs: 17, 17 -> 18
			// srcs: (1, 0)(20) -3, (76) 0 --> (131) 0:ND0, NW0, *, PENB
			6'd0 : rdata = 41'b00011011000000000100000000000000100000000;
			// PEs: 16 -> 
			// srcs: (16, 1)(173) -4 --> (173) -4:PENB, pass, 
			6'd1 : rdata = 41'b11000110111111100000000000000000000000000;
			// PEs: 17, 16 -> 16
			// srcs: (23, 2)(173) -4, (121) 1 --> (174) -3:ALU, PENB, +, PEGB0
			6'd2 : rdata = 41'b00001001111111111101111111000000010000000;
			// PEs: 16, 18 -> 16
			// srcs: (24, 3)(183) -6, (184) -2 --> (185) -8:PENB, PEGB2, +, PEGB0
			6'd3 : rdata = 41'b00001110111111101110000010000000010000000;
			// PEs: 16 -> 
			// srcs: (32, 4)(214) 5 --> (214) 5:PENB, pass, 
			6'd4 : rdata = 41'b11000110111111100000000000000000000000000;
			// PEs: 16, 17 -> 16
			// srcs: (38, 5)(212) -1, (214) 5 --> (215) 4:PENB, ALU, +, PEGB0
			6'd5 : rdata = 41'b00001110111111100011111111100000010000000;
			// PEs: 16, 17 -> 18
			// srcs: (122, 6)(224) 3, (20) -3 --> (241) -9:PENB, ND0, *, PENB
			6'd6 : rdata = 41'b00011110111111100110000000000000100000000;
			// PEs: 17, 18 -> 17
			// srcs: (131, 7)(76) 0, (296) -9 --> (351) 9:NW0, PEGB2, -, NW0
			6'd7 : rdata = 41'b00010010000000001110000010000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 18) begin
	always @(*) begin
		case(address)
			// PEs: 18, 18 -> 
			// srcs: (1, 0)(21) -1, (77) 2 --> (132) -2:ND0, NW0, *, 
			6'd0 : rdata = 41'b00011011000000000100000000000000000000000;
			// PEs: 17, 18 -> 17
			// srcs: (4, 1)(131) 0, (132) -2 --> (184) -2:PENB, ALU, +, PEGB1
			6'd1 : rdata = 41'b00001110111111100011111111100000010010000;
			// PEs: 18, 17 -> 17
			// srcs: (125, 3)(3) 1, (241) -9 --> (296) -9:NM0, PENB, *, PEGB1
			6'd2 : rdata = 41'b00011100000000001101111111000000010010000;
			// PEs: 16, 18 -> 19
			// srcs: (126, 2)(224) 3, (21) -1 --> (242) -3:PEGB0, ND0, *, PENB
			6'd3 : rdata = 41'b00011111000000000110000000000000100000000;
			// PEs: 18, 19 -> 18
			// srcs: (135, 4)(77) 2, (297) -3 --> (352) 5:NW0, PEGB3, -, NW0
			6'd4 : rdata = 41'b00010010000000001110000011000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 19) begin
	always @(*) begin
		case(address)
			// PEs: 19, 19 -> 20
			// srcs: (1, 0)(22) 1, (78) 0 --> (133) 0:ND0, NW0, *, PENB
			6'd0 : rdata = 41'b00011011000000000100000000000000100000000;
			// PEs: 16, 19 -> 19
			// srcs: (127, 1)(224) 3, (22) 1 --> (243) 3:PEGB0, ND0, *, NI0
			6'd1 : rdata = 41'b00011111000000000110000000010000000000000;
			// PEs: 19, 18 -> 18
			// srcs: (129, 2)(3) 1, (242) -3 --> (297) -3:NM0, PENB, *, PEGB2
			6'd2 : rdata = 41'b00011100000000001101111111000000010100000;
			// PEs: 19, 19 -> 
			// srcs: (130, 3)(3) 1, (243) 3 --> (298) 3:NM0, NI0, *, 
			6'd3 : rdata = 41'b00011100000000001010000000000000000000000;
			// PEs: 19, 19 -> 19
			// srcs: (133, 4)(78) 0, (298) 3 --> (353) -3:NW0, ALU, -, NW0
			6'd4 : rdata = 41'b00010010000000000011111111100100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 20) begin
	always @(*) begin
		case(address)
			// PEs: 20, 20 -> 
			// srcs: (1, 0)(23) 0, (79) 0 --> (134) 0:ND0, NW0, *, 
			6'd0 : rdata = 41'b00011011000000000100000000000000000000000;
			// PEs: 19, 20 -> 16
			// srcs: (4, 1)(133) 0, (134) 0 --> (186) 0:PENB, ALU, +, PEGB0
			6'd1 : rdata = 41'b00001110111111100011111111100000010000000;
			// PEs: 16, 20 -> 21
			// srcs: (128, 2)(224) 3, (23) 0 --> (244) 0:PEGB0, ND0, *, PENB
			6'd2 : rdata = 41'b00011111000000000110000000000000100000000;
			// PEs: 20, 21 -> 20
			// srcs: (137, 3)(79) 0, (299) 0 --> (354) 0:NW0, PEGB5, -, NW0
			6'd3 : rdata = 41'b00010010000000001110000101000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 21) begin
	always @(*) begin
		case(address)
			// PEs: 21, 21 -> 22
			// srcs: (1, 0)(25) -1, (81) 1 --> (136) -1:ND0, NW0, *, PENB
			6'd0 : rdata = 41'b00011011000000000100000000000000100000000;
			// PEs: 16, 21 -> 21
			// srcs: (130, 1)(224) 3, (25) -1 --> (246) -3:PEGB0, ND0, *, NI0
			6'd1 : rdata = 41'b00011111000000000110000000010000000000000;
			// PEs: 21, 20 -> 20
			// srcs: (131, 2)(3) 1, (244) 0 --> (299) 0:NM0, PENB, *, PEGB4
			6'd2 : rdata = 41'b00011100000000001101111111000000011000000;
			// PEs: 21, 21 -> 
			// srcs: (133, 3)(3) 1, (246) -3 --> (301) -3:NM0, NI0, *, 
			6'd3 : rdata = 41'b00011100000000001010000000000000000000000;
			// PEs: 21, 21 -> 21
			// srcs: (136, 4)(81) 1, (301) -3 --> (356) 4:NW0, ALU, -, NW0
			6'd4 : rdata = 41'b00010010000000000011111111100100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 22) begin
	always @(*) begin
		case(address)
			// PEs: 22, 22 -> 
			// srcs: (1, 0)(26) -2, (82) -2 --> (137) 4:ND0, NW0, *, 
			6'd0 : rdata = 41'b00011011000000000100000000000000000000000;
			// PEs: 21, 22 -> 16
			// srcs: (4, 1)(136) -1, (137) 4 --> (189) 3:PENB, ALU, +, PEGB0
			6'd1 : rdata = 41'b00001110111111100011111111100000010000000;
			// PEs: 16, 22 -> 23
			// srcs: (131, 2)(224) 3, (26) -2 --> (247) -6:PEGB0, ND0, *, PENB
			6'd2 : rdata = 41'b00011111000000000110000000000000100000000;
			// PEs: 22, 23 -> 22
			// srcs: (140, 3)(82) -2, (302) -6 --> (357) 4:NW0, PEGB7, -, NW0
			6'd3 : rdata = 41'b00010010000000001110000111000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 23) begin
	always @(*) begin
		case(address)
			// PEs: 23, 23 -> 16
			// srcs: (1, 0)(27) -3, (83) 0 --> (138) 0:ND0, NW0, *, PENB
			6'd0 : rdata = 41'b00011011000000000100000000000000100000000;
			// PEs: 16, 23 -> 23
			// srcs: (132, 1)(224) 3, (27) -3 --> (248) -9:PEGB0, ND0, *, NI0
			6'd1 : rdata = 41'b00011111000000000110000000010000000000000;
			// PEs: 23, 22 -> 22
			// srcs: (134, 2)(3) 1, (247) -6 --> (302) -6:NM0, PENB, *, PEGB6
			6'd2 : rdata = 41'b00011100000000001101111111000000011100000;
			// PEs: 23, 23 -> 
			// srcs: (135, 3)(3) 1, (248) -9 --> (303) -9:NM0, NI0, *, 
			6'd3 : rdata = 41'b00011100000000001010000000000000000000000;
			// PEs: 23, 23 -> 23
			// srcs: (138, 4)(83) 0, (303) -9 --> (358) 9:NW0, ALU, -, NW0
			6'd4 : rdata = 41'b00010010000000000011111111100100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 24) begin
	always @(*) begin
		case(address)
			// PEs: 16 -> 25
			// srcs: (5, 0)(138) 0 --> (138) 0:PUNB, pass, PENB
			6'd0 : rdata = 41'b11000110111111110000000000000000100000000;
			// PEs: 27 -> 48
			// srcs: (9, 5)(192) -1 --> (192) -1:PEGB3, pass, PUGB6
			6'd1 : rdata = 41'b11000111000001100000000000000000000001110;
			// PEs: 16 -> 24
			// srcs: (11, 1)(186) 0 --> (186) 0:PUNB, pass, NI0
			6'd2 : rdata = 41'b11000110111111110000000000010000000000000;
			// PEs: 48 -> 25
			// srcs: (12, 2)(135) -4 --> (135) -4:PUGB6, pass, PENB
			6'd3 : rdata = 41'b11000111000011010000000000000000100000000;
			// PEs: 26 -> 48
			// srcs: (17, 8)(199) 9 --> (199) 9:PEGB2, pass, PUGB6
			6'd4 : rdata = 41'b11000111000001000000000000000000000001110;
			// PEs: 24 -> 25
			// srcs: (18, 3)(186) 0 --> (186) 0:NI0, pass, PENB
			6'd5 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 16 -> 25
			// srcs: (19, 4)(189) 3 --> (189) 3:PUNB, pass, PENB
			6'd6 : rdata = 41'b11000110111111110000000000000000100000000;
			// PEs: 25 -> 32
			// srcs: (26, 7)(191) 0 --> (191) 0:PEGB1, pass, PUNB
			6'd7 : rdata = 41'b11000111000000100000000000000001000000000;
			// PEs: 16 -> 25
			// srcs: (31, 6)(185) -8 --> (185) -8:PUNB, pass, PENB
			6'd8 : rdata = 41'b11000110111111110000000000000000100000000;
			// PEs: 25 -> 32
			// srcs: (39, 9)(188) -12 --> (188) -12:PEGB1, pass, PUNB
			6'd9 : rdata = 41'b11000111000000100000000000000001000000000;
			// PEs: 48 -> 25
			// srcs: (128, 10)(224) 3 --> (224) 3:PUGB6, pass, PENB
			6'd10 : rdata = 41'b11000111000011010000000000000000100000000;
			// PEs: 48 -> 26
			// srcs: (129, 11)(224) 3 --> (224) 3:PUGB6, pass, PEGB2
			6'd11 : rdata = 41'b11000111000011010000000000000000010100000;
			// PEs: 48 -> 27
			// srcs: (130, 12)(224) 3 --> (224) 3:PUGB6, pass, PEGB3
			6'd12 : rdata = 41'b11000111000011010000000000000000010110000;
			// PEs: 48 -> 28
			// srcs: (132, 13)(224) 3 --> (224) 3:PUGB6, pass, PEGB4
			6'd13 : rdata = 41'b11000111000011010000000000000000011000000;
			// PEs: 48 -> 29
			// srcs: (133, 14)(224) 3 --> (224) 3:PUGB6, pass, PEGB5
			6'd14 : rdata = 41'b11000111000011010000000000000000011010000;
			// PEs: 48 -> 30
			// srcs: (134, 15)(224) 3 --> (224) 3:PUGB6, pass, PEGB6
			6'd15 : rdata = 41'b11000111000011010000000000000000011100000;
			// PEs: 48 -> 31
			// srcs: (135, 16)(224) 3 --> (224) 3:PUGB6, pass, PEGB7
			6'd16 : rdata = 41'b11000111000011010000000000000000011110000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 25) begin
	always @(*) begin
		case(address)
			// PEs: 25, 25 -> 
			// srcs: (1, 0)(28) 1, (84) -3 --> (139) -3:ND0, NW0, *, 
			6'd0 : rdata = 41'b00011011000000000100000000000000000000000;
			// PEs: 24, 25 -> 25
			// srcs: (8, 1)(138) 0, (139) -3 --> (190) -3:PENB, ALU, +, NI0
			6'd1 : rdata = 41'b00001110111111100011111111110000000000000;
			// PEs: 24 -> 
			// srcs: (14, 2)(135) -4 --> (135) -4:PENB, pass, 
			6'd2 : rdata = 41'b11000110111111100000000000000000000000000;
			// PEs: 24, 25 -> 25
			// srcs: (20, 3)(186) 0, (135) -4 --> (187) -4:PENB, ALU, +, NI1
			6'd3 : rdata = 41'b00001110111111100011111111111000000000000;
			// PEs: 24, 25 -> 24
			// srcs: (21, 4)(189) 3, (190) -3 --> (191) 0:PENB, NI0, +, PEGB0
			6'd4 : rdata = 41'b00001110111111101010000000000000010000000;
			// PEs: 24, 25 -> 24
			// srcs: (34, 5)(185) -8, (187) -4 --> (188) -12:PENB, NI1, +, PEGB0
			6'd5 : rdata = 41'b00001110111111101010000000100000010000000;
			// PEs: 24, 25 -> 26
			// srcs: (130, 6)(224) 3, (28) 1 --> (249) 3:PENB, ND0, *, PENB
			6'd6 : rdata = 41'b00011110111111100110000000000000100000000;
			// PEs: 25, 26 -> 25
			// srcs: (139, 7)(84) -3, (304) 3 --> (359) -6:NW0, PEGB2, -, NW0
			6'd7 : rdata = 41'b00010010000000001110000010000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 26) begin
	always @(*) begin
		case(address)
			// PEs: 26, 26 -> 27
			// srcs: (1, 0)(29) 0, (85) -3 --> (140) 0:ND0, NW0, *, PENB
			6'd0 : rdata = 41'b00011011000000000100000000000000100000000;
			// PEs: 31 -> 
			// srcs: (9, 1)(198) 10 --> (198) 10:PEGB7, pass, 
			6'd1 : rdata = 41'b11000111000011100000000000000000000000000;
			// PEs: 29, 26 -> 24
			// srcs: (12, 2)(197) -1, (198) 10 --> (199) 9:PEGB5, ALU, +, PEGB0
			6'd2 : rdata = 41'b00001111000010100011111111100000010000000;
			// PEs: 26, 25 -> 25
			// srcs: (133, 4)(3) 1, (249) 3 --> (304) 3:NM0, PENB, *, PEGB1
			6'd3 : rdata = 41'b00011100000000001101111111000000010010000;
			// PEs: 24, 26 -> 27
			// srcs: (134, 3)(224) 3, (29) 0 --> (250) 0:PEGB0, ND0, *, PENB
			6'd4 : rdata = 41'b00011111000000000110000000000000100000000;
			// PEs: 26, 27 -> 26
			// srcs: (143, 5)(85) -3, (305) 0 --> (360) -3:NW0, PEGB3, -, NW0
			6'd5 : rdata = 41'b00010010000000001110000011000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 27) begin
	always @(*) begin
		case(address)
			// PEs: 27, 27 -> 
			// srcs: (1, 0)(30) 1, (86) -1 --> (141) -1:ND0, NW0, *, 
			6'd0 : rdata = 41'b00011011000000000100000000000000000000000;
			// PEs: 26, 27 -> 24
			// srcs: (4, 1)(140) 0, (141) -1 --> (192) -1:PENB, ALU, +, PEGB0
			6'd1 : rdata = 41'b00001110111111100011111111100000010000000;
			// PEs: 24, 27 -> 28
			// srcs: (135, 2)(224) 3, (30) 1 --> (251) 3:PEGB0, ND0, *, PENB
			6'd2 : rdata = 41'b00011111000000000110000000000000100000000;
			// PEs: 27, 26 -> 26
			// srcs: (137, 3)(3) 1, (250) 0 --> (305) 0:NM0, PENB, *, PEGB2
			6'd3 : rdata = 41'b00011100000000001101111111000000010100000;
			// PEs: 27, 28 -> 27
			// srcs: (144, 4)(86) -1, (306) 3 --> (361) -4:NW0, PEGB4, -, NW0
			6'd4 : rdata = 41'b00010010000000001110000100000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 28) begin
	always @(*) begin
		case(address)
			// PEs: 28, 28 -> 29
			// srcs: (1, 0)(32) 0, (88) 2 --> (143) 0:ND0, NW0, *, PENB
			6'd0 : rdata = 41'b00011011000000000100000000000000100000000;
			// PEs: 24, 28 -> 28
			// srcs: (137, 1)(224) 3, (32) 0 --> (253) 0:PEGB0, ND0, *, NI0
			6'd1 : rdata = 41'b00011111000000000110000000010000000000000;
			// PEs: 28, 27 -> 27
			// srcs: (138, 2)(3) 1, (251) 3 --> (306) 3:NM0, PENB, *, PEGB3
			6'd2 : rdata = 41'b00011100000000001101111111000000010110000;
			// PEs: 28, 28 -> 
			// srcs: (140, 3)(3) 1, (253) 0 --> (308) 0:NM0, NI0, *, 
			6'd3 : rdata = 41'b00011100000000001010000000000000000000000;
			// PEs: 28, 28 -> 28
			// srcs: (143, 4)(88) 2, (308) 0 --> (363) 2:NW0, ALU, -, NW0
			6'd4 : rdata = 41'b00010010000000000011111111100100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 29) begin
	always @(*) begin
		case(address)
			// PEs: 29, 29 -> 
			// srcs: (1, 0)(33) 1, (89) -1 --> (144) -1:ND0, NW0, *, 
			6'd0 : rdata = 41'b00011011000000000100000000000000000000000;
			// PEs: 28, 29 -> 26
			// srcs: (4, 1)(143) 0, (144) -1 --> (197) -1:PENB, ALU, +, PEGB2
			6'd1 : rdata = 41'b00001110111111100011111111100000010100000;
			// PEs: 24, 29 -> 30
			// srcs: (138, 2)(224) 3, (33) 1 --> (254) 3:PEGB0, ND0, *, PENB
			6'd2 : rdata = 41'b00011111000000000110000000000000100000000;
			// PEs: 29, 30 -> 29
			// srcs: (147, 3)(89) -1, (309) 3 --> (364) -4:NW0, PEGB6, -, NW0
			6'd3 : rdata = 41'b00010010000000001110000110000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 30) begin
	always @(*) begin
		case(address)
			// PEs: 30, 30 -> 31
			// srcs: (1, 0)(34) -1, (90) -1 --> (145) 1:ND0, NW0, *, PENB
			6'd0 : rdata = 41'b00011011000000000100000000000000100000000;
			// PEs: 24, 30 -> 30
			// srcs: (139, 1)(224) 3, (34) -1 --> (255) -3:PEGB0, ND0, *, NI0
			6'd1 : rdata = 41'b00011111000000000110000000010000000000000;
			// PEs: 30, 29 -> 29
			// srcs: (141, 2)(3) 1, (254) 3 --> (309) 3:NM0, PENB, *, PEGB5
			6'd2 : rdata = 41'b00011100000000001101111111000000011010000;
			// PEs: 30, 30 -> 
			// srcs: (142, 3)(3) 1, (255) -3 --> (310) -3:NM0, NI0, *, 
			6'd3 : rdata = 41'b00011100000000001010000000000000000000000;
			// PEs: 30, 30 -> 30
			// srcs: (145, 4)(90) -1, (310) -3 --> (365) 2:NW0, ALU, -, NW0
			6'd4 : rdata = 41'b00010010000000000011111111100100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 31) begin
	always @(*) begin
		case(address)
			// PEs: 31, 31 -> 
			// srcs: (1, 0)(35) -3, (91) -3 --> (146) 9:ND0, NW0, *, 
			6'd0 : rdata = 41'b00011011000000000100000000000000000000000;
			// PEs: 30, 31 -> 26
			// srcs: (4, 1)(145) 1, (146) 9 --> (198) 10:PENB, ALU, +, PEGB2
			6'd1 : rdata = 41'b00001110111111100011111111100000010100000;
			// PEs: 24, 31 -> 
			// srcs: (140, 2)(224) 3, (35) -3 --> (256) -9:PEGB0, ND0, *, 
			6'd2 : rdata = 41'b00011111000000000110000000000000000000000;
			// PEs: 31, 31 -> 
			// srcs: (143, 3)(3) 1, (256) -9 --> (311) -9:NM0, ALU, *, 
			6'd3 : rdata = 41'b00011100000000000011111111100000000000000;
			// PEs: 31, 31 -> 31
			// srcs: (146, 4)(91) -3, (311) -9 --> (366) 6:NW0, ALU, -, NW0
			6'd4 : rdata = 41'b00010010000000000011111111100100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 32) begin
	always @(*) begin
		case(address)
			// PEs: 39 -> 40
			// srcs: (3, 0)(154) -2 --> (154) -2:PENB, pass, PUNB
			6'd0 : rdata = 41'b11000110111111100000000000000001000000000;
			// PEs: 34 -> 56
			// srcs: (9, 4)(200) -2 --> (200) -2:PEGB2, pass, PUGB7
			6'd1 : rdata = 41'b11000111000001000000000000000000000001111;
			// PEs: 48 -> 32
			// srcs: (12, 2)(128) 2 --> (128) 2:PUGB6, pass, NI0
			6'd2 : rdata = 41'b11000111000011010000000000010000000000000;
			// PEs: 8 -> 33
			// srcs: (14, 1)(179) 0 --> (179) 0:PUGB1, pass, PENB
			6'd3 : rdata = 41'b11000111000000110000000000000000100000000;
			// PEs: 35 -> 8
			// srcs: (17, 9)(205) -4 --> (205) -4:PEGB3, pass, PUGB1
			6'd4 : rdata = 41'b11000111000001100000000000000000000001001;
			// PEs: 32 -> 33
			// srcs: (21, 3)(128) 2 --> (128) 2:NI0, pass, PENB
			6'd5 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 33 -> 0
			// srcs: (28, 5)(180) 2 --> (180) 2:PEGB1, pass, PUGB0
			6'd6 : rdata = 41'b11000111000000100000000000000000000001000;
			// PEs: 24 -> 32
			// srcs: (29, 6)(191) 0 --> (191) 0:PUNB, pass, NI0
			6'd7 : rdata = 41'b11000110111111110000000000010000000000000;
			// PEs: 48 -> 33
			// srcs: (33, 7)(193) 3 --> (193) 3:PUGB6, pass, PENB
			6'd8 : rdata = 41'b11000111000011010000000000000000100000000;
			// PEs: 32 -> 33
			// srcs: (40, 8)(191) 0 --> (191) 0:NI0, pass, PENB
			6'd9 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 24 -> 33
			// srcs: (41, 10)(188) -12 --> (188) -12:PUNB, pass, PENB
			6'd10 : rdata = 41'b11000110111111110000000000000000100000000;
			// PEs: 33 -> 40
			// srcs: (57, 11)(195) -9 --> (195) -9:PEGB1, pass, PUNB
			6'd11 : rdata = 41'b11000111000000100000000000000001000000000;
			// PEs: 48 -> 33
			// srcs: (136, 12)(224) 3 --> (224) 3:PUGB6, pass, PENB
			6'd12 : rdata = 41'b11000111000011010000000000000000100000000;
			// PEs: 48 -> 34
			// srcs: (137, 13)(224) 3 --> (224) 3:PUGB6, pass, PEGB2
			6'd13 : rdata = 41'b11000111000011010000000000000000010100000;
			// PEs: 48 -> 35
			// srcs: (139, 14)(224) 3 --> (224) 3:PUGB6, pass, PEGB3
			6'd14 : rdata = 41'b11000111000011010000000000000000010110000;
			// PEs: 48 -> 36
			// srcs: (140, 15)(224) 3 --> (224) 3:PUGB6, pass, PEGB4
			6'd15 : rdata = 41'b11000111000011010000000000000000011000000;
			// PEs: 48 -> 37
			// srcs: (141, 16)(224) 3 --> (224) 3:PUGB6, pass, PEGB5
			6'd16 : rdata = 41'b11000111000011010000000000000000011010000;
			// PEs: 48 -> 38
			// srcs: (142, 17)(224) 3 --> (224) 3:PUGB6, pass, PEGB6
			6'd17 : rdata = 41'b11000111000011010000000000000000011100000;
			// PEs: 48 -> 39
			// srcs: (143, 18)(224) 3 --> (224) 3:PUGB6, pass, PEGB7
			6'd18 : rdata = 41'b11000111000011010000000000000000011110000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 33) begin
	always @(*) begin
		case(address)
			// PEs: 33, 33 -> 34
			// srcs: (1, 0)(36) 1, (92) -2 --> (147) -2:ND0, NW0, *, PENB
			6'd0 : rdata = 41'b00011011000000000100000000000000100000000;
			// PEs: 32 -> 
			// srcs: (16, 1)(179) 0 --> (179) 0:PENB, pass, 
			6'd1 : rdata = 41'b11000110111111100000000000000000000000000;
			// PEs: 33, 32 -> 32
			// srcs: (23, 2)(179) 0, (128) 2 --> (180) 2:ALU, PENB, +, PEGB0
			6'd2 : rdata = 41'b00001001111111111101111111000000010000000;
			// PEs: 32 -> 
			// srcs: (35, 3)(193) 3 --> (193) 3:PENB, pass, 
			6'd3 : rdata = 41'b11000110111111100000000000000000000000000;
			// PEs: 32, 33 -> 
			// srcs: (42, 4)(191) 0, (193) 3 --> (194) 3:PENB, ALU, +, 
			6'd4 : rdata = 41'b00001110111111100011111111100000000000000;
			// PEs: 32, 33 -> 32
			// srcs: (52, 5)(188) -12, (194) 3 --> (195) -9:PENB, ALU, +, PEGB0
			6'd5 : rdata = 41'b00001110111111100011111111100000010000000;
			// PEs: 32, 33 -> 34
			// srcs: (138, 6)(224) 3, (36) 1 --> (257) 3:PENB, ND0, *, PENB
			6'd6 : rdata = 41'b00011110111111100110000000000000100000000;
			// PEs: 33, 34 -> 33
			// srcs: (147, 7)(92) -2, (312) 3 --> (367) -5:NW0, PEGB2, -, NW0
			6'd7 : rdata = 41'b00010010000000001110000010000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 34) begin
	always @(*) begin
		case(address)
			// PEs: 34, 34 -> 
			// srcs: (1, 0)(37) 0, (93) 1 --> (148) 0:ND0, NW0, *, 
			6'd0 : rdata = 41'b00011011000000000100000000000000000000000;
			// PEs: 33, 34 -> 32
			// srcs: (4, 1)(147) -2, (148) 0 --> (200) -2:PENB, ALU, +, PEGB0
			6'd1 : rdata = 41'b00001110111111100011111111100000010000000;
			// PEs: 34, 33 -> 33
			// srcs: (141, 3)(3) 1, (257) 3 --> (312) 3:NM0, PENB, *, PEGB1
			6'd2 : rdata = 41'b00011100000000001101111111000000010010000;
			// PEs: 32, 34 -> 
			// srcs: (142, 2)(224) 3, (37) 0 --> (258) 0:PEGB0, ND0, *, 
			6'd3 : rdata = 41'b00011111000000000110000000000000000000000;
			// PEs: 34, 34 -> 
			// srcs: (145, 4)(3) 1, (258) 0 --> (313) 0:NM0, ALU, *, 
			6'd4 : rdata = 41'b00011100000000000011111111100000000000000;
			// PEs: 34, 34 -> 34
			// srcs: (148, 5)(93) 1, (313) 0 --> (368) 1:NW0, ALU, -, NW0
			6'd5 : rdata = 41'b00010010000000000011111111100100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 35) begin
	always @(*) begin
		case(address)
			// PEs: 35, 35 -> 36
			// srcs: (1, 0)(39) 2, (95) -1 --> (150) -2:ND0, NW0, *, PENB
			6'd0 : rdata = 41'b00011011000000000100000000000000100000000;
			// PEs: 38 -> 
			// srcs: (9, 1)(204) -2 --> (204) -2:PEGB6, pass, 
			6'd1 : rdata = 41'b11000111000011000000000000000000000000000;
			// PEs: 36, 35 -> 32
			// srcs: (12, 2)(203) -2, (204) -2 --> (205) -4:PEGB4, ALU, +, PEGB0
			6'd2 : rdata = 41'b00001111000010000011111111100000010000000;
			// PEs: 32, 35 -> 36
			// srcs: (144, 3)(224) 3, (39) 2 --> (260) 6:PEGB0, ND0, *, PENB
			6'd3 : rdata = 41'b00011111000000000110000000000000100000000;
			// PEs: 35, 36 -> 35
			// srcs: (153, 4)(95) -1, (315) 6 --> (370) -7:NW0, PEGB4, -, NW0
			6'd4 : rdata = 41'b00010010000000001110000100000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 36) begin
	always @(*) begin
		case(address)
			// PEs: 36, 36 -> 
			// srcs: (1, 0)(40) 0, (96) -1 --> (151) 0:ND0, NW0, *, 
			6'd0 : rdata = 41'b00011011000000000100000000000000000000000;
			// PEs: 35, 36 -> 35
			// srcs: (4, 1)(150) -2, (151) 0 --> (203) -2:PENB, ALU, +, PEGB3
			6'd1 : rdata = 41'b00001110111111100011111111100000010110000;
			// PEs: 32, 36 -> 37
			// srcs: (145, 2)(224) 3, (40) 0 --> (261) 0:PEGB0, ND0, *, PENB
			6'd2 : rdata = 41'b00011111000000000110000000000000100000000;
			// PEs: 36, 35 -> 35
			// srcs: (147, 3)(3) 1, (260) 6 --> (315) 6:NM0, PENB, *, PEGB3
			6'd3 : rdata = 41'b00011100000000001101111111000000010110000;
			// PEs: 36, 37 -> 36
			// srcs: (154, 4)(96) -1, (316) 0 --> (371) -1:NW0, PEGB5, -, NW0
			6'd4 : rdata = 41'b00010010000000001110000101000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 37) begin
	always @(*) begin
		case(address)
			// PEs: 37, 37 -> 38
			// srcs: (1, 0)(41) 1, (97) -2 --> (152) -2:ND0, NW0, *, PENB
			6'd0 : rdata = 41'b00011011000000000100000000000000100000000;
			// PEs: 32, 37 -> 37
			// srcs: (146, 1)(224) 3, (41) 1 --> (262) 3:PEGB0, ND0, *, NI0
			6'd1 : rdata = 41'b00011111000000000110000000010000000000000;
			// PEs: 37, 36 -> 36
			// srcs: (148, 2)(3) 1, (261) 0 --> (316) 0:NM0, PENB, *, PEGB4
			6'd2 : rdata = 41'b00011100000000001101111111000000011000000;
			// PEs: 37, 37 -> 
			// srcs: (149, 3)(3) 1, (262) 3 --> (317) 3:NM0, NI0, *, 
			6'd3 : rdata = 41'b00011100000000001010000000000000000000000;
			// PEs: 37, 37 -> 37
			// srcs: (152, 4)(97) -2, (317) 3 --> (372) -5:NW0, ALU, -, NW0
			6'd4 : rdata = 41'b00010010000000000011111111100100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 38) begin
	always @(*) begin
		case(address)
			// PEs: 38, 38 -> 
			// srcs: (1, 0)(42) 0, (98) -3 --> (153) 0:ND0, NW0, *, 
			6'd0 : rdata = 41'b00011011000000000100000000000000000000000;
			// PEs: 37, 38 -> 35
			// srcs: (4, 1)(152) -2, (153) 0 --> (204) -2:PENB, ALU, +, PEGB3
			6'd1 : rdata = 41'b00001110111111100011111111100000010110000;
			// PEs: 32, 38 -> 39
			// srcs: (147, 2)(224) 3, (42) 0 --> (263) 0:PEGB0, ND0, *, PENB
			6'd2 : rdata = 41'b00011111000000000110000000000000100000000;
			// PEs: 38, 39 -> 38
			// srcs: (156, 3)(98) -3, (318) 0 --> (373) -3:NW0, PEGB7, -, NW0
			6'd3 : rdata = 41'b00010010000000001110000111000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 39) begin
	always @(*) begin
		case(address)
			// PEs: 39, 39 -> 32
			// srcs: (1, 0)(43) -1, (99) 2 --> (154) -2:ND0, NW0, *, PENB
			6'd0 : rdata = 41'b00011011000000000100000000000000100000000;
			// PEs: 32, 39 -> 39
			// srcs: (148, 1)(224) 3, (43) -1 --> (264) -3:PEGB0, ND0, *, NI0
			6'd1 : rdata = 41'b00011111000000000110000000010000000000000;
			// PEs: 39, 38 -> 38
			// srcs: (150, 2)(3) 1, (263) 0 --> (318) 0:NM0, PENB, *, PEGB6
			6'd2 : rdata = 41'b00011100000000001101111111000000011100000;
			// PEs: 39, 39 -> 
			// srcs: (151, 3)(3) 1, (264) -3 --> (319) -3:NM0, NI0, *, 
			6'd3 : rdata = 41'b00011100000000001010000000000000000000000;
			// PEs: 39, 39 -> 39
			// srcs: (154, 4)(99) 2, (319) -3 --> (374) 5:NW0, ALU, -, NW0
			6'd4 : rdata = 41'b00010010000000000011111111100100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 40) begin
	always @(*) begin
		case(address)
			// PEs: 32 -> 41
			// srcs: (5, 0)(154) -2 --> (154) -2:PUNB, pass, PENB
			6'd0 : rdata = 41'b11000110111111110000000000000000100000000;
			// PEs: 47 -> 56
			// srcs: (6, 2)(213) 3 --> (213) 3:PENB, pass, PUGB7
			6'd1 : rdata = 41'b11000110111111100000000000000000000001111;
			// PEs: 41 -> 8
			// srcs: (13, 1)(206) 1 --> (206) 1:PEGB1, pass, PUGB1
			6'd2 : rdata = 41'b11000111000000100000000000000000000001001;
			// PEs: 42 -> 16
			// srcs: (17, 6)(212) -1 --> (212) -1:PEGB2, pass, PUGB2
			6'd3 : rdata = 41'b11000111000001000000000000000000000001010;
			// PEs: 0 -> 40
			// srcs: (22, 3)(172) -6 --> (172) -6:PUGB0, pass, NI0
			6'd4 : rdata = 41'b11000111000000010000000000010000000000000;
			// PEs: 16 -> 41
			// srcs: (33, 4)(174) -3 --> (174) -3:PUGB2, pass, PENB
			6'd5 : rdata = 41'b11000111000001010000000000000000100000000;
			// PEs: 40 -> 41
			// srcs: (40, 5)(172) -6 --> (172) -6:NI0, pass, PENB
			6'd6 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 0 -> 41
			// srcs: (52, 7)(181) -2 --> (181) -2:PUGB0, pass, PENB
			6'd7 : rdata = 41'b11000111000000010000000000000000100000000;
			// PEs: 32 -> 41
			// srcs: (59, 8)(195) -9 --> (195) -9:PUNB, pass, PENB
			6'd8 : rdata = 41'b11000110111111110000000000000000100000000;
			// PEs: 41 -> 48
			// srcs: (70, 9)(196) -20 --> (196) -20:PEGB1, pass, PUNB
			6'd9 : rdata = 41'b11000111000000100000000000000001000000000;
			// PEs: 48 -> 41
			// srcs: (144, 10)(224) 3 --> (224) 3:PUGB6, pass, PENB
			6'd10 : rdata = 41'b11000111000011010000000000000000100000000;
			// PEs: 48 -> 42
			// srcs: (146, 11)(224) 3 --> (224) 3:PUGB6, pass, PEGB2
			6'd11 : rdata = 41'b11000111000011010000000000000000010100000;
			// PEs: 48 -> 43
			// srcs: (147, 12)(224) 3 --> (224) 3:PUGB6, pass, PEGB3
			6'd12 : rdata = 41'b11000111000011010000000000000000010110000;
			// PEs: 48 -> 44
			// srcs: (148, 13)(224) 3 --> (224) 3:PUGB6, pass, PEGB4
			6'd13 : rdata = 41'b11000111000011010000000000000000011000000;
			// PEs: 48 -> 45
			// srcs: (149, 14)(224) 3 --> (224) 3:PUGB6, pass, PEGB5
			6'd14 : rdata = 41'b11000111000011010000000000000000011010000;
			// PEs: 48 -> 46
			// srcs: (150, 15)(224) 3 --> (224) 3:PUGB6, pass, PEGB6
			6'd15 : rdata = 41'b11000111000011010000000000000000011100000;
			// PEs: 48 -> 47
			// srcs: (151, 16)(224) 3 --> (224) 3:PUGB6, pass, PEGB7
			6'd16 : rdata = 41'b11000111000011010000000000000000011110000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 41) begin
	always @(*) begin
		case(address)
			// PEs: 41, 41 -> 
			// srcs: (1, 0)(44) -3, (100) -1 --> (155) 3:ND0, NW0, *, 
			6'd0 : rdata = 41'b00011011000000000100000000000000000000000;
			// PEs: 40, 41 -> 40
			// srcs: (8, 1)(154) -2, (155) 3 --> (206) 1:PENB, ALU, +, PEGB0
			6'd1 : rdata = 41'b00001110111111100011111111100000010000000;
			// PEs: 40 -> 
			// srcs: (35, 2)(174) -3 --> (174) -3:PENB, pass, 
			6'd2 : rdata = 41'b11000110111111100000000000000000000000000;
			// PEs: 40, 41 -> 
			// srcs: (42, 3)(172) -6, (174) -3 --> (175) -9:PENB, ALU, +, 
			6'd3 : rdata = 41'b00001110111111100011111111100000000000000;
			// PEs: 41, 40 -> 
			// srcs: (55, 4)(175) -9, (181) -2 --> (182) -11:ALU, PENB, +, 
			6'd4 : rdata = 41'b00001001111111111101111111000000000000000;
			// PEs: 41, 40 -> 40
			// srcs: (65, 5)(182) -11, (195) -9 --> (196) -20:ALU, PENB, +, PEGB0
			6'd5 : rdata = 41'b00001001111111111101111111000000010000000;
			// PEs: 40, 41 -> 42
			// srcs: (146, 6)(224) 3, (44) -3 --> (265) -9:PENB, ND0, *, PENB
			6'd6 : rdata = 41'b00011110111111100110000000000000100000000;
			// PEs: 41, 42 -> 41
			// srcs: (155, 7)(100) -1, (320) -9 --> (375) 8:NW0, PEGB2, -, NW0
			6'd7 : rdata = 41'b00010010000000001110000010000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 42) begin
	always @(*) begin
		case(address)
			// PEs: 42, 42 -> 43
			// srcs: (1, 0)(46) 2, (102) -3 --> (157) -6:ND0, NW0, *, PENB
			6'd0 : rdata = 41'b00011011000000000100000000000000100000000;
			// PEs: 45 -> 
			// srcs: (9, 1)(211) -1 --> (211) -1:PEGB5, pass, 
			6'd1 : rdata = 41'b11000111000010100000000000000000000000000;
			// PEs: 43, 42 -> 40
			// srcs: (12, 2)(210) 0, (211) -1 --> (212) -1:PEGB3, ALU, +, PEGB0
			6'd2 : rdata = 41'b00001111000001100011111111100000010000000;
			// PEs: 42, 41 -> 41
			// srcs: (149, 4)(3) 1, (265) -9 --> (320) -9:NM0, PENB, *, PEGB1
			6'd3 : rdata = 41'b00011100000000001101111111000000010010000;
			// PEs: 40, 42 -> 43
			// srcs: (151, 3)(224) 3, (46) 2 --> (267) 6:PEGB0, ND0, *, PENB
			6'd4 : rdata = 41'b00011111000000000110000000000000100000000;
			// PEs: 42, 43 -> 42
			// srcs: (160, 5)(102) -3, (322) 6 --> (377) -9:NW0, PEGB3, -, NW0
			6'd5 : rdata = 41'b00010010000000001110000011000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 43) begin
	always @(*) begin
		case(address)
			// PEs: 43, 43 -> 
			// srcs: (1, 0)(47) -2, (103) -3 --> (158) 6:ND0, NW0, *, 
			6'd0 : rdata = 41'b00011011000000000100000000000000000000000;
			// PEs: 42, 43 -> 42
			// srcs: (4, 1)(157) -6, (158) 6 --> (210) 0:PENB, ALU, +, PEGB2
			6'd1 : rdata = 41'b00001110111111100011111111100000010100000;
			// PEs: 40, 43 -> 44
			// srcs: (152, 2)(224) 3, (47) -2 --> (268) -6:PEGB0, ND0, *, PENB
			6'd2 : rdata = 41'b00011111000000000110000000000000100000000;
			// PEs: 43, 42 -> 42
			// srcs: (154, 3)(3) 1, (267) 6 --> (322) 6:NM0, PENB, *, PEGB2
			6'd3 : rdata = 41'b00011100000000001101111111000000010100000;
			// PEs: 43, 44 -> 43
			// srcs: (161, 4)(103) -3, (323) -6 --> (378) 3:NW0, PEGB4, -, NW0
			6'd4 : rdata = 41'b00010010000000001110000100000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 44) begin
	always @(*) begin
		case(address)
			// PEs: 44, 44 -> 45
			// srcs: (1, 0)(48) -3, (104) 1 --> (159) -3:ND0, NW0, *, PENB
			6'd0 : rdata = 41'b00011011000000000100000000000000100000000;
			// PEs: 40, 44 -> 44
			// srcs: (153, 1)(224) 3, (48) -3 --> (269) -9:PEGB0, ND0, *, NI0
			6'd1 : rdata = 41'b00011111000000000110000000010000000000000;
			// PEs: 44, 43 -> 43
			// srcs: (155, 2)(3) 1, (268) -6 --> (323) -6:NM0, PENB, *, PEGB3
			6'd2 : rdata = 41'b00011100000000001101111111000000010110000;
			// PEs: 44, 44 -> 
			// srcs: (156, 3)(3) 1, (269) -9 --> (324) -9:NM0, NI0, *, 
			6'd3 : rdata = 41'b00011100000000001010000000000000000000000;
			// PEs: 44, 44 -> 44
			// srcs: (159, 4)(104) 1, (324) -9 --> (379) 10:NW0, ALU, -, NW0
			6'd4 : rdata = 41'b00010010000000000011111111100100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 45) begin
	always @(*) begin
		case(address)
			// PEs: 45, 45 -> 
			// srcs: (1, 0)(49) -2, (105) -1 --> (160) 2:ND0, NW0, *, 
			6'd0 : rdata = 41'b00011011000000000100000000000000000000000;
			// PEs: 44, 45 -> 42
			// srcs: (4, 1)(159) -3, (160) 2 --> (211) -1:PENB, ALU, +, PEGB2
			6'd1 : rdata = 41'b00001110111111100011111111100000010100000;
			// PEs: 40, 45 -> 46
			// srcs: (154, 2)(224) 3, (49) -2 --> (270) -6:PEGB0, ND0, *, PENB
			6'd2 : rdata = 41'b00011111000000000110000000000000100000000;
			// PEs: 45, 46 -> 45
			// srcs: (163, 3)(105) -1, (325) -6 --> (380) 5:NW0, PEGB6, -, NW0
			6'd3 : rdata = 41'b00010010000000001110000110000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 46) begin
	always @(*) begin
		case(address)
			// PEs: 46, 46 -> 47
			// srcs: (1, 0)(50) -3, (106) -1 --> (161) 3:ND0, NW0, *, PENB
			6'd0 : rdata = 41'b00011011000000000100000000000000100000000;
			// PEs: 40, 46 -> 46
			// srcs: (155, 1)(224) 3, (50) -3 --> (271) -9:PEGB0, ND0, *, NI0
			6'd1 : rdata = 41'b00011111000000000110000000010000000000000;
			// PEs: 46, 45 -> 45
			// srcs: (157, 2)(3) 1, (270) -6 --> (325) -6:NM0, PENB, *, PEGB5
			6'd2 : rdata = 41'b00011100000000001101111111000000011010000;
			// PEs: 46, 46 -> 
			// srcs: (158, 3)(3) 1, (271) -9 --> (326) -9:NM0, NI0, *, 
			6'd3 : rdata = 41'b00011100000000001010000000000000000000000;
			// PEs: 46, 46 -> 46
			// srcs: (161, 4)(106) -1, (326) -9 --> (381) 8:NW0, ALU, -, NW0
			6'd4 : rdata = 41'b00010010000000000011111111100100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 47) begin
	always @(*) begin
		case(address)
			// PEs: 47, 47 -> 
			// srcs: (1, 0)(51) 0, (107) 1 --> (162) 0:ND0, NW0, *, 
			6'd0 : rdata = 41'b00011011000000000100000000000000000000000;
			// PEs: 46, 47 -> 40
			// srcs: (4, 1)(161) 3, (162) 0 --> (213) 3:PENB, ALU, +, PENB
			6'd1 : rdata = 41'b00001110111111100011111111100000100000000;
			// PEs: 40, 47 -> 
			// srcs: (156, 2)(224) 3, (51) 0 --> (272) 0:PEGB0, ND0, *, 
			6'd2 : rdata = 41'b00011111000000000110000000000000000000000;
			// PEs: 47, 47 -> 
			// srcs: (159, 3)(3) 1, (272) 0 --> (327) 0:NM0, ALU, *, 
			6'd3 : rdata = 41'b00011100000000000011111111100000000000000;
			// PEs: 47, 47 -> 47
			// srcs: (162, 4)(107) 1, (327) 0 --> (382) 1:NW0, ALU, -, NW0
			6'd4 : rdata = 41'b00010010000000000011111111100100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 48) begin
	always @(*) begin
		case(address)
			// PEs: 55 -> 24
			// srcs: (3, 2)(135) -4 --> (135) -4:PENB, pass, PUGB3
			6'd0 : rdata = 41'b11000110111111100000000000000000000001011;
			// PEs: 53 -> 16
			// srcs: (6, 0)(121) 1 --> (121) 1:PEGB5, pass, PUGB2
			6'd1 : rdata = 41'b11000111000010100000000000000000000001010;
			// PEs: 54 -> 32
			// srcs: (7, 1)(128) 2 --> (128) 2:PEGB6, pass, PUGB4
			6'd2 : rdata = 41'b11000111000011000000000000000000000001100;
			// PEs: 50 -> 56
			// srcs: (9, 6)(216) 9 --> (216) 9:PEGB2, pass, PUNB
			6'd3 : rdata = 41'b11000111000001000000000000000001000000000;
			// PEs: 52 -> 56
			// srcs: (10, 7)(218) 2 --> (218) 2:PEGB4, pass, PUNB
			6'd4 : rdata = 41'b11000111000010000000000000000001000000000;
			// PEs: 56 -> 48
			// srcs: (11, 4)(142) 4 --> (142) 4:PUGB7, pass, NI0
			6'd5 : rdata = 41'b11000111000011110000000000010000000000000;
			// PEs: 24 -> 49
			// srcs: (14, 3)(192) -1 --> (192) -1:PUGB3, pass, PENB
			6'd6 : rdata = 41'b11000111000001110000000000000000100000000;
			// PEs: 48 -> 49
			// srcs: (21, 5)(142) 4 --> (142) 4:NI0, pass, PENB
			6'd7 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 24 -> 48
			// srcs: (22, 9)(199) 9 --> (199) 9:PUGB3, pass, NI0
			6'd8 : rdata = 41'b11000111000001110000000000010000000000000;
			// PEs: 56 -> 49
			// srcs: (27, 10)(201) 0 --> (201) 0:PUGB7, pass, PENB
			6'd9 : rdata = 41'b11000111000011110000000000000000100000000;
			// PEs: 49 -> 32
			// srcs: (28, 8)(193) 3 --> (193) 3:PEGB1, pass, PUGB4
			6'd10 : rdata = 41'b11000111000000100000000000000000000001100;
			// PEs: 48 -> 49
			// srcs: (34, 11)(199) 9 --> (199) 9:NI0, pass, PENB
			6'd11 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 49 -> 0
			// srcs: (41, 12)(202) 9 --> (202) 9:PEGB1, pass, PUGB0
			6'd12 : rdata = 41'b11000111000000100000000000000000000001000;
			// PEs: 40 -> 48
			// srcs: (72, 13)(196) -20 --> (196) -20:PUNB, pass, NI0
			6'd13 : rdata = 41'b11000110111111110000000000010000000000000;
			// PEs: 8 -> 49
			// srcs: (79, 14)(222) 23 --> (222) 23:PUGB1, pass, PENB
			6'd14 : rdata = 41'b11000111000000110000000000000000100000000;
			// PEs: 48 -> 49
			// srcs: (86, 15)(196) -20 --> (196) -20:NI0, pass, PENB
			6'd15 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 50 -> 0
			// srcs: (96, 16)(224) 3 --> (224) 3:PEGB2, pass, PUGB0
			6'd16 : rdata = 41'b11000111000001000000000000000000000001000;
			// PEs: 50 -> 0
			// srcs: (100, 17)(224) 3 --> (224) 3:PEGB2, pass, PUGB0
			6'd17 : rdata = 41'b11000111000001000000000000000000000001000;
			// PEs: 50 -> 0
			// srcs: (101, 18)(224) 3 --> (224) 3:PEGB2, pass, PUGB0
			6'd18 : rdata = 41'b11000111000001000000000000000000000001000;
			// PEs: 50 -> 0
			// srcs: (102, 19)(224) 3 --> (224) 3:PEGB2, pass, PUGB0
			6'd19 : rdata = 41'b11000111000001000000000000000000000001000;
			// PEs: 50 -> 0
			// srcs: (103, 20)(224) 3 --> (224) 3:PEGB2, pass, PUGB0
			6'd20 : rdata = 41'b11000111000001000000000000000000000001000;
			// PEs: 50 -> 0
			// srcs: (104, 21)(224) 3 --> (224) 3:PEGB2, pass, PUGB0
			6'd21 : rdata = 41'b11000111000001000000000000000000000001000;
			// PEs: 50 -> 0
			// srcs: (106, 22)(224) 3 --> (224) 3:PEGB2, pass, PUGB0
			6'd22 : rdata = 41'b11000111000001000000000000000000000001000;
			// PEs: 50 -> 8
			// srcs: (107, 23)(224) 3 --> (224) 3:PEGB2, pass, PUGB1
			6'd23 : rdata = 41'b11000111000001000000000000000000000001001;
			// PEs: 50 -> 8
			// srcs: (108, 24)(224) 3 --> (224) 3:PEGB2, pass, PUGB1
			6'd24 : rdata = 41'b11000111000001000000000000000000000001001;
			// PEs: 50 -> 8
			// srcs: (109, 25)(224) 3 --> (224) 3:PEGB2, pass, PUGB1
			6'd25 : rdata = 41'b11000111000001000000000000000000000001001;
			// PEs: 50 -> 8
			// srcs: (110, 26)(224) 3 --> (224) 3:PEGB2, pass, PUGB1
			6'd26 : rdata = 41'b11000111000001000000000000000000000001001;
			// PEs: 50 -> 8
			// srcs: (111, 27)(224) 3 --> (224) 3:PEGB2, pass, PUGB1
			6'd27 : rdata = 41'b11000111000001000000000000000000000001001;
			// PEs: 50 -> 8
			// srcs: (113, 28)(224) 3 --> (224) 3:PEGB2, pass, PUGB1
			6'd28 : rdata = 41'b11000111000001000000000000000000000001001;
			// PEs: 50 -> 8
			// srcs: (114, 29)(224) 3 --> (224) 3:PEGB2, pass, PUGB1
			6'd29 : rdata = 41'b11000111000001000000000000000000000001001;
			// PEs: 50 -> 16
			// srcs: (115, 30)(224) 3 --> (224) 3:PEGB2, pass, PUGB2
			6'd30 : rdata = 41'b11000111000001000000000000000000000001010;
			// PEs: 50 -> 16
			// srcs: (116, 31)(224) 3 --> (224) 3:PEGB2, pass, PUGB2
			6'd31 : rdata = 41'b11000111000001000000000000000000000001010;
			// PEs: 50 -> 16
			// srcs: (117, 32)(224) 3 --> (224) 3:PEGB2, pass, PUGB2
			6'd32 : rdata = 41'b11000111000001000000000000000000000001010;
			// PEs: 50 -> 16
			// srcs: (118, 33)(224) 3 --> (224) 3:PEGB2, pass, PUGB2
			6'd33 : rdata = 41'b11000111000001000000000000000000000001010;
			// PEs: 50 -> 16
			// srcs: (120, 34)(224) 3 --> (224) 3:PEGB2, pass, PUGB2
			6'd34 : rdata = 41'b11000111000001000000000000000000000001010;
			// PEs: 50 -> 16
			// srcs: (121, 35)(224) 3 --> (224) 3:PEGB2, pass, PUGB2
			6'd35 : rdata = 41'b11000111000001000000000000000000000001010;
			// PEs: 50 -> 16
			// srcs: (122, 36)(224) 3 --> (224) 3:PEGB2, pass, PUGB2
			6'd36 : rdata = 41'b11000111000001000000000000000000000001010;
			// PEs: 50 -> 24
			// srcs: (123, 37)(224) 3 --> (224) 3:PEGB2, pass, PUGB3
			6'd37 : rdata = 41'b11000111000001000000000000000000000001011;
			// PEs: 50 -> 24
			// srcs: (124, 38)(224) 3 --> (224) 3:PEGB2, pass, PUGB3
			6'd38 : rdata = 41'b11000111000001000000000000000000000001011;
			// PEs: 50 -> 24
			// srcs: (125, 39)(224) 3 --> (224) 3:PEGB2, pass, PUGB3
			6'd39 : rdata = 41'b11000111000001000000000000000000000001011;
			// PEs: 50 -> 56
			// srcs: (126, 40)(224) 3 --> (224) 3:PEGB2, pass, PUNB
			6'd40 : rdata = 41'b11000111000001000000000000000001000000000;
			// PEs: 50 -> 24
			// srcs: (127, 41)(224) 3 --> (224) 3:PEGB2, pass, PUGB3
			6'd41 : rdata = 41'b11000111000001000000000000000000000001011;
			// PEs: 50 -> 24
			// srcs: (128, 42)(224) 3 --> (224) 3:PEGB2, pass, PUGB3
			6'd42 : rdata = 41'b11000111000001000000000000000000000001011;
			// PEs: 50 -> 24
			// srcs: (129, 43)(224) 3 --> (224) 3:PEGB2, pass, PUGB3
			6'd43 : rdata = 41'b11000111000001000000000000000000000001011;
			// PEs: 50 -> 24
			// srcs: (130, 44)(224) 3 --> (224) 3:PEGB2, pass, PUGB3
			6'd44 : rdata = 41'b11000111000001000000000000000000000001011;
			// PEs: 50 -> 32
			// srcs: (131, 45)(224) 3 --> (224) 3:PEGB2, pass, PUGB4
			6'd45 : rdata = 41'b11000111000001000000000000000000000001100;
			// PEs: 50 -> 32
			// srcs: (132, 46)(224) 3 --> (224) 3:PEGB2, pass, PUGB4
			6'd46 : rdata = 41'b11000111000001000000000000000000000001100;
			// PEs: 50 -> 56
			// srcs: (133, 47)(224) 3 --> (224) 3:PEGB2, pass, PUNB
			6'd47 : rdata = 41'b11000111000001000000000000000001000000000;
			// PEs: 50 -> 32
			// srcs: (134, 48)(224) 3 --> (224) 3:PEGB2, pass, PUGB4
			6'd48 : rdata = 41'b11000111000001000000000000000000000001100;
			// PEs: 50 -> 32
			// srcs: (135, 49)(224) 3 --> (224) 3:PEGB2, pass, PUGB4
			6'd49 : rdata = 41'b11000111000001000000000000000000000001100;
			// PEs: 50 -> 32
			// srcs: (136, 50)(224) 3 --> (224) 3:PEGB2, pass, PUGB4
			6'd50 : rdata = 41'b11000111000001000000000000000000000001100;
			// PEs: 50 -> 32
			// srcs: (137, 51)(224) 3 --> (224) 3:PEGB2, pass, PUGB4
			6'd51 : rdata = 41'b11000111000001000000000000000000000001100;
			// PEs: 50 -> 32
			// srcs: (138, 52)(224) 3 --> (224) 3:PEGB2, pass, PUGB4
			6'd52 : rdata = 41'b11000111000001000000000000000000000001100;
			// PEs: 50 -> 40
			// srcs: (139, 53)(224) 3 --> (224) 3:PEGB2, pass, PUGB5
			6'd53 : rdata = 41'b11000111000001000000000000000000000001101;
			// PEs: 50 -> 56
			// srcs: (140, 54)(224) 3 --> (224) 3:PEGB2, pass, PUNB
			6'd54 : rdata = 41'b11000111000001000000000000000001000000000;
			// PEs: 50 -> 40
			// srcs: (141, 55)(224) 3 --> (224) 3:PEGB2, pass, PUGB5
			6'd55 : rdata = 41'b11000111000001000000000000000000000001101;
			// PEs: 50 -> 40
			// srcs: (142, 56)(224) 3 --> (224) 3:PEGB2, pass, PUGB5
			6'd56 : rdata = 41'b11000111000001000000000000000000000001101;
			// PEs: 50 -> 40
			// srcs: (143, 57)(224) 3 --> (224) 3:PEGB2, pass, PUGB5
			6'd57 : rdata = 41'b11000111000001000000000000000000000001101;
			// PEs: 50 -> 40
			// srcs: (144, 58)(224) 3 --> (224) 3:PEGB2, pass, PUGB5
			6'd58 : rdata = 41'b11000111000001000000000000000000000001101;
			// PEs: 50 -> 40
			// srcs: (145, 59)(224) 3 --> (224) 3:PEGB2, pass, PUGB5
			6'd59 : rdata = 41'b11000111000001000000000000000000000001101;
			// PEs: 50 -> 40
			// srcs: (146, 60)(224) 3 --> (224) 3:PEGB2, pass, PUGB5
			6'd60 : rdata = 41'b11000111000001000000000000000000000001101;
			// PEs: 50 -> 56
			// srcs: (147, 61)(224) 3 --> (224) 3:PEGB2, pass, PUNB
			6'd61 : rdata = 41'b11000111000001000000000000000001000000000;
			// PEs: 50 -> 56
			// srcs: (150, 62)(224) 3 --> (224) 3:PEGB2, pass, PUNB
			6'd62 : rdata = 41'b11000111000001000000000000000001000000000;
			// PEs: 50 -> 56
			// srcs: (152, 63)(224) 3 --> (224) 3:PEGB2, pass, PUNB
			6'd63 : rdata = 41'b11000111000001000000000000000001000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 49) begin
	always @(*) begin
		case(address)
			// PEs: 49, 49 -> 50
			// srcs: (1, 0)(53) -3, (109) -3 --> (164) 9:ND0, NW0, *, PENB
			6'd0 : rdata = 41'b00011011000000000100000000000000100000000;
			// PEs: 48 -> 
			// srcs: (16, 1)(192) -1 --> (192) -1:PENB, pass, 
			6'd1 : rdata = 41'b11000110111111100000000000000000000000000;
			// PEs: 49, 48 -> 48
			// srcs: (23, 2)(192) -1, (142) 4 --> (193) 3:ALU, PENB, +, PEGB0
			6'd2 : rdata = 41'b00001001111111111101111111000000010000000;
			// PEs: 48 -> 
			// srcs: (29, 3)(201) 0 --> (201) 0:PENB, pass, 
			6'd3 : rdata = 41'b11000110111111100000000000000000000000000;
			// PEs: 48, 49 -> 48
			// srcs: (36, 4)(199) 9, (201) 0 --> (202) 9:PENB, ALU, +, PEGB0
			6'd4 : rdata = 41'b00001110111111100011111111100000010000000;
			// PEs: 48 -> 
			// srcs: (81, 5)(222) 23 --> (222) 23:PENB, pass, 
			6'd5 : rdata = 41'b11000110111111100000000000000000000000000;
			// PEs: 48, 49 -> 50
			// srcs: (88, 6)(196) -20, (222) 23 --> (223) 3:PENB, ALU, +, PENB
			6'd6 : rdata = 41'b00001110111111100011111111100000100000000;
			// PEs: 50, 49 -> 
			// srcs: (148, 7)(224) 3, (53) -3 --> (274) -9:PEGB2, ND0, *, 
			6'd7 : rdata = 41'b00011111000001000110000000000000000000000;
			// PEs: 49, 49 -> 
			// srcs: (151, 8)(3) 1, (274) -9 --> (329) -9:NM0, ALU, *, 
			6'd8 : rdata = 41'b00011100000000000011111111100000000000000;
			// PEs: 49, 49 -> 49
			// srcs: (154, 9)(109) -3, (329) -9 --> (384) 6:NW0, ALU, -, NW0
			6'd9 : rdata = 41'b00010010000000000011111111100100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 50) begin
	always @(*) begin
		case(address)
			// PEs: 50, 50 -> 
			// srcs: (1, 0)(54) 2, (110) 0 --> (165) 0:ND0, NW0, *, 
			6'd0 : rdata = 41'b00011011000000000100000000000000000000000;
			// PEs: 49, 50 -> 48
			// srcs: (4, 1)(164) 9, (165) 0 --> (216) 9:PENB, ALU, +, PEGB0
			6'd1 : rdata = 41'b00001110111111100011111111100000010000000;
			// PEs: 49, 50 -> 51, 48, 50
			// srcs: (91, 2)(223) 3, (59) 0 --> (224) 3:PENB, ND1, -, NI0, PENB, PEGB0
			6'd2 : rdata = 41'b00010110111111100110000000110000110000000;
			// PEs: 50 -> 48
			// srcs: (93, 3)(224) 3 --> (224) 3:ALU, pass, PEGB0
			6'd3 : rdata = 41'b11000001111111110000000000000000010000000;
			// PEs: 50 -> 48
			// srcs: (94, 4)(224) 3 --> (224) 3:NI0, pass, PEGB0
			6'd4 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 50 -> 48
			// srcs: (95, 5)(224) 3 --> (224) 3:NI0, pass, PEGB0
			6'd5 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 50 -> 48
			// srcs: (96, 6)(224) 3 --> (224) 3:NI0, pass, PEGB0
			6'd6 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 50 -> 48
			// srcs: (97, 7)(224) 3 --> (224) 3:NI0, pass, PEGB0
			6'd7 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 50 -> 53
			// srcs: (98, 8)(224) 3 --> (224) 3:NI0, pass, PEGB5
			6'd8 : rdata = 41'b11000101000000000000000000000000011010000;
			// PEs: 50 -> 48
			// srcs: (99, 9)(224) 3 --> (224) 3:NI0, pass, PEGB0
			6'd9 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 50 -> 48
			// srcs: (100, 10)(224) 3 --> (224) 3:NI0, pass, PEGB0
			6'd10 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 50 -> 48
			// srcs: (101, 11)(224) 3 --> (224) 3:NI0, pass, PEGB0
			6'd11 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 50 -> 48
			// srcs: (102, 12)(224) 3 --> (224) 3:NI0, pass, PEGB0
			6'd12 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 50 -> 48
			// srcs: (103, 13)(224) 3 --> (224) 3:NI0, pass, PEGB0
			6'd13 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 50 -> 48
			// srcs: (104, 14)(224) 3 --> (224) 3:NI0, pass, PEGB0
			6'd14 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 50 -> 54
			// srcs: (105, 15)(224) 3 --> (224) 3:NI0, pass, PEGB6
			6'd15 : rdata = 41'b11000101000000000000000000000000011100000;
			// PEs: 50 -> 48
			// srcs: (106, 16)(224) 3 --> (224) 3:NI0, pass, PEGB0
			6'd16 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 50 -> 48
			// srcs: (107, 17)(224) 3 --> (224) 3:NI0, pass, PEGB0
			6'd17 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 50 -> 48
			// srcs: (108, 18)(224) 3 --> (224) 3:NI0, pass, PEGB0
			6'd18 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 50 -> 48
			// srcs: (109, 19)(224) 3 --> (224) 3:NI0, pass, PEGB0
			6'd19 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 50 -> 48
			// srcs: (110, 20)(224) 3 --> (224) 3:NI0, pass, PEGB0
			6'd20 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 50 -> 48
			// srcs: (111, 21)(224) 3 --> (224) 3:NI0, pass, PEGB0
			6'd21 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 50 -> 55
			// srcs: (112, 22)(224) 3 --> (224) 3:NI0, pass, PEGB7
			6'd22 : rdata = 41'b11000101000000000000000000000000011110000;
			// PEs: 50 -> 48
			// srcs: (113, 23)(224) 3 --> (224) 3:NI0, pass, PEGB0
			6'd23 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 50 -> 48
			// srcs: (114, 24)(224) 3 --> (224) 3:NI0, pass, PEGB0
			6'd24 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 50 -> 48
			// srcs: (115, 25)(224) 3 --> (224) 3:NI0, pass, PEGB0
			6'd25 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 50 -> 48
			// srcs: (116, 26)(224) 3 --> (224) 3:NI0, pass, PEGB0
			6'd26 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 50 -> 48
			// srcs: (117, 27)(224) 3 --> (224) 3:NI0, pass, PEGB0
			6'd27 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 50 -> 48
			// srcs: (118, 28)(224) 3 --> (224) 3:NI0, pass, PEGB0
			6'd28 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 50 -> 48
			// srcs: (119, 29)(224) 3 --> (224) 3:NI0, pass, PEGB0
			6'd29 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 50 -> 48
			// srcs: (120, 30)(224) 3 --> (224) 3:NI0, pass, PEGB0
			6'd30 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 50 -> 48
			// srcs: (121, 31)(224) 3 --> (224) 3:NI0, pass, PEGB0
			6'd31 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 50 -> 48
			// srcs: (122, 32)(224) 3 --> (224) 3:NI0, pass, PEGB0
			6'd32 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 50 -> 48
			// srcs: (123, 33)(224) 3 --> (224) 3:NI0, pass, PEGB0
			6'd33 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 50 -> 48
			// srcs: (124, 34)(224) 3 --> (224) 3:NI0, pass, PEGB0
			6'd34 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 50 -> 48
			// srcs: (125, 35)(224) 3 --> (224) 3:NI0, pass, PEGB0
			6'd35 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 50 -> 48
			// srcs: (126, 36)(224) 3 --> (224) 3:NI0, pass, PEGB0
			6'd36 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 50 -> 48
			// srcs: (127, 37)(224) 3 --> (224) 3:NI0, pass, PEGB0
			6'd37 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 50 -> 48
			// srcs: (128, 38)(224) 3 --> (224) 3:NI0, pass, PEGB0
			6'd38 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 50 -> 48
			// srcs: (129, 39)(224) 3 --> (224) 3:NI0, pass, PEGB0
			6'd39 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 50 -> 48
			// srcs: (130, 40)(224) 3 --> (224) 3:NI0, pass, PEGB0
			6'd40 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 50 -> 48
			// srcs: (131, 41)(224) 3 --> (224) 3:NI0, pass, PEGB0
			6'd41 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 50 -> 48
			// srcs: (132, 42)(224) 3 --> (224) 3:NI0, pass, PEGB0
			6'd42 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 50 -> 48
			// srcs: (133, 43)(224) 3 --> (224) 3:NI0, pass, PEGB0
			6'd43 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 50 -> 48
			// srcs: (134, 44)(224) 3 --> (224) 3:NI0, pass, PEGB0
			6'd44 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 50 -> 48
			// srcs: (135, 45)(224) 3 --> (224) 3:NI0, pass, PEGB0
			6'd45 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 50 -> 48
			// srcs: (136, 46)(224) 3 --> (224) 3:NI0, pass, PEGB0
			6'd46 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 50 -> 48
			// srcs: (137, 47)(224) 3 --> (224) 3:NI0, pass, PEGB0
			6'd47 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 50 -> 48
			// srcs: (138, 48)(224) 3 --> (224) 3:NI0, pass, PEGB0
			6'd48 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 50 -> 48
			// srcs: (139, 49)(224) 3 --> (224) 3:NI0, pass, PEGB0
			6'd49 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 50 -> 48
			// srcs: (140, 50)(224) 3 --> (224) 3:NI0, pass, PEGB0
			6'd50 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 50 -> 49
			// srcs: (141, 51)(224) 3 --> (224) 3:NI0, pass, PEGB1
			6'd51 : rdata = 41'b11000101000000000000000000000000010010000;
			// PEs: 50, 50 -> 51
			// srcs: (142, 52)(224) 3, (54) 2 --> (275) 6:NI0, ND0, *, PENB
			6'd52 : rdata = 41'b00011101000000000110000000000000100000000;
			// PEs: 50 -> 48
			// srcs: (143, 53)(224) 3 --> (224) 3:NI0, pass, PEGB0
			6'd53 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 50 -> 52
			// srcs: (144, 54)(224) 3 --> (224) 3:NI0, pass, PEGB4
			6'd54 : rdata = 41'b11000101000000000000000000000000011000000;
			// PEs: 50 -> 48
			// srcs: (145, 55)(224) 3 --> (224) 3:NI0, pass, PEGB0
			6'd55 : rdata = 41'b11000101000000000000000000000000010000000;
			// PEs: 50, 51 -> 50
			// srcs: (151, 56)(110) 0, (330) 6 --> (385) -6:NW0, PEGB3, -, NW0
			6'd56 : rdata = 41'b00010010000000001110000011000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 51) begin
	always @(*) begin
		case(address)
			// PEs: 51, 51 -> 52
			// srcs: (1, 0)(56) 2, (112) 1 --> (167) 2:ND0, NW0, *, PENB
			6'd0 : rdata = 41'b00011011000000000100000000000000100000000;
			// PEs: 50, 51 -> 
			// srcs: (94, 1)(224) 3, (56) 2 --> (277) 6:PENB, ND0, *, 
			6'd1 : rdata = 41'b00011110111111100110000000000000000000000;
			// PEs: 51, 51 -> 
			// srcs: (97, 3)(3) 1, (277) 6 --> (332) 6:NM0, ALU, *, 
			6'd2 : rdata = 41'b00011100000000000011111111100000000000000;
			// PEs: 51, 51 -> 51
			// srcs: (100, 4)(112) 1, (332) 6 --> (387) -5:NW0, ALU, -, NW0
			6'd3 : rdata = 41'b00010010000000000011111111100100000000000;
			// PEs: 51, 50 -> 50
			// srcs: (145, 2)(3) 1, (275) 6 --> (330) 6:NM0, PENB, *, PEGB2
			6'd4 : rdata = 41'b00011100000000001101111111000000010100000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 52) begin
	always @(*) begin
		case(address)
			// PEs: 52, 52 -> 
			// srcs: (1, 0)(57) 0, (113) 1 --> (168) 0:ND0, NW0, *, 
			6'd0 : rdata = 41'b00011011000000000100000000000000000000000;
			// PEs: 51, 52 -> 48
			// srcs: (4, 1)(167) 2, (168) 0 --> (218) 2:PENB, ALU, +, PEGB0
			6'd1 : rdata = 41'b00001110111111100011111111100000010000000;
			// PEs: 50, 52 -> 
			// srcs: (151, 2)(224) 3, (57) 0 --> (278) 0:PEGB2, ND0, *, 
			6'd2 : rdata = 41'b00011111000001000110000000000000000000000;
			// PEs: 52, 52 -> 
			// srcs: (154, 3)(3) 1, (278) 0 --> (333) 0:NM0, ALU, *, 
			6'd3 : rdata = 41'b00011100000000000011111111100000000000000;
			// PEs: 52, 52 -> 52
			// srcs: (157, 4)(113) 1, (333) 0 --> (388) 1:NW0, ALU, -, NW0
			6'd4 : rdata = 41'b00010010000000000011111111100100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 53) begin
	always @(*) begin
		case(address)
			// PEs: 53, 53 -> 48
			// srcs: (1, 0)(10) -1, (66) -1 --> (121) 1:ND0, NW0, *, PEGB0
			6'd0 : rdata = 41'b00011011000000000100000000000000010000000;
			// PEs: 50, 53 -> 
			// srcs: (105, 1)(224) 3, (10) -1 --> (231) -3:PEGB2, ND0, *, 
			6'd1 : rdata = 41'b00011111000001000110000000000000000000000;
			// PEs: 53, 53 -> 
			// srcs: (108, 2)(3) 1, (231) -3 --> (286) -3:NM0, ALU, *, 
			6'd2 : rdata = 41'b00011100000000000011111111100000000000000;
			// PEs: 53, 53 -> 53
			// srcs: (111, 3)(66) -1, (286) -3 --> (341) 2:NW0, ALU, -, NW0
			6'd3 : rdata = 41'b00010010000000000011111111100100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 54) begin
	always @(*) begin
		case(address)
			// PEs: 54, 54 -> 48
			// srcs: (1, 0)(17) -2, (73) -1 --> (128) 2:ND0, NW0, *, PEGB0
			6'd0 : rdata = 41'b00011011000000000100000000000000010000000;
			// PEs: 50, 54 -> 
			// srcs: (112, 1)(224) 3, (17) -2 --> (238) -6:PEGB2, ND0, *, 
			6'd1 : rdata = 41'b00011111000001000110000000000000000000000;
			// PEs: 54, 54 -> 
			// srcs: (115, 2)(3) 1, (238) -6 --> (293) -6:NM0, ALU, *, 
			6'd2 : rdata = 41'b00011100000000000011111111100000000000000;
			// PEs: 54, 54 -> 54
			// srcs: (118, 3)(73) -1, (293) -6 --> (348) 5:NW0, ALU, -, NW0
			6'd3 : rdata = 41'b00010010000000000011111111100100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 55) begin
	always @(*) begin
		case(address)
			// PEs: 55, 55 -> 48
			// srcs: (1, 0)(24) -2, (80) 2 --> (135) -4:ND0, NW0, *, PENB
			6'd0 : rdata = 41'b00011011000000000100000000000000100000000;
			// PEs: 50, 55 -> 
			// srcs: (119, 1)(224) 3, (24) -2 --> (245) -6:PEGB2, ND0, *, 
			6'd1 : rdata = 41'b00011111000001000110000000000000000000000;
			// PEs: 55, 55 -> 
			// srcs: (122, 2)(3) 1, (245) -6 --> (300) -6:NM0, ALU, *, 
			6'd2 : rdata = 41'b00011100000000000011111111100000000000000;
			// PEs: 55, 55 -> 55
			// srcs: (125, 3)(80) 2, (300) -6 --> (355) 8:NW0, ALU, -, NW0
			6'd3 : rdata = 41'b00010010000000000011111111100100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 56) begin
	always @(*) begin
		case(address)
			// PEs: 57 -> 48
			// srcs: (6, 0)(142) 4 --> (142) 4:PEGB1, pass, PUGB6
			6'd0 : rdata = 41'b11000111000000100000000000000000000001110;
			// PEs: 59 -> 8
			// srcs: (7, 2)(156) 0 --> (156) 0:PEGB3, pass, PUGB1
			6'd1 : rdata = 41'b11000111000001100000000000000000000001001;
			// PEs: 32 -> 57
			// srcs: (14, 1)(200) -2 --> (200) -2:PUGB4, pass, PENB
			6'd2 : rdata = 41'b11000111000010010000000000000000100000000;
			// PEs: 40 -> 57
			// srcs: (15, 3)(213) 3 --> (213) 3:PUGB5, pass, PENB
			6'd3 : rdata = 41'b11000111000010110000000000000000100000000;
			// PEs: 48 -> 57
			// srcs: (16, 4)(216) 9 --> (216) 9:PUNB, pass, PENB
			6'd4 : rdata = 41'b11000110111111110000000000000000100000000;
			// PEs: 48 -> 57
			// srcs: (17, 5)(218) 2 --> (218) 2:PUNB, pass, PENB
			6'd5 : rdata = 41'b11000110111111110000000000000000100000000;
			// PEs: 57 -> 48
			// srcs: (22, 6)(201) 0 --> (201) 0:PEGB1, pass, PUGB6
			6'd6 : rdata = 41'b11000111000000100000000000000000000001110;
			// PEs: 57 -> 16
			// srcs: (23, 7)(214) 5 --> (214) 5:PEGB1, pass, PUGB2
			6'd7 : rdata = 41'b11000111000000100000000000000000000001010;
			// PEs: 58 -> 8
			// srcs: (34, 8)(220) 13 --> (220) 13:PEGB2, pass, PUGB1
			6'd8 : rdata = 41'b11000111000001000000000000000000000001001;
			// PEs: 48 -> 57
			// srcs: (128, 9)(224) 3 --> (224) 3:PUNB, pass, PENB
			6'd9 : rdata = 41'b11000110111111110000000000000000100000000;
			// PEs: 48 -> 58
			// srcs: (135, 10)(224) 3 --> (224) 3:PUNB, pass, PEGB2
			6'd10 : rdata = 41'b11000110111111110000000000000000010100000;
			// PEs: 48 -> 59
			// srcs: (142, 11)(224) 3 --> (224) 3:PUNB, pass, PEGB3
			6'd11 : rdata = 41'b11000110111111110000000000000000010110000;
			// PEs: 48 -> 60
			// srcs: (149, 12)(224) 3 --> (224) 3:PUNB, pass, PEGB4
			6'd12 : rdata = 41'b11000110111111110000000000000000011000000;
			// PEs: 48 -> 61
			// srcs: (152, 13)(224) 3 --> (224) 3:PUNB, pass, PEGB5
			6'd13 : rdata = 41'b11000110111111110000000000000000011010000;
			// PEs: 48 -> 62
			// srcs: (154, 14)(224) 3 --> (224) 3:PUNB, pass, PEGB6
			6'd14 : rdata = 41'b11000110111111110000000000000000011100000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 57) begin
	always @(*) begin
		case(address)
			// PEs: 57, 57 -> 56
			// srcs: (1, 0)(31) 2, (87) 2 --> (142) 4:ND0, NW0, *, PEGB0
			6'd0 : rdata = 41'b00011011000000000100000000000000010000000;
			// PEs: 56, 58 -> 56
			// srcs: (17, 1)(200) -2, (149) 2 --> (201) 0:PENB, PEGB2, +, PEGB0
			6'd1 : rdata = 41'b00001110111111101110000010000000010000000;
			// PEs: 56, 60 -> 56
			// srcs: (18, 2)(213) 3, (163) 2 --> (214) 5:PENB, PEGB4, +, PEGB0
			6'd2 : rdata = 41'b00001110111111101110000100000000010000000;
			// PEs: 56, 61 -> 57
			// srcs: (19, 3)(216) 9, (166) 2 --> (217) 11:PENB, PEGB5, +, NI0
			6'd3 : rdata = 41'b00001110111111101110000101010000000000000;
			// PEs: 56, 62 -> 58
			// srcs: (20, 4)(218) 2, (169) 0 --> (219) 2:PENB, PEGB6, +, PENB
			6'd4 : rdata = 41'b00001110111111101110000110000000100000000;
			// PEs: 57 -> 58
			// srcs: (27, 5)(217) 11 --> (217) 11:NI0, pass, PENB
			6'd5 : rdata = 41'b11000101000000000000000000000000100000000;
			// PEs: 56, 57 -> 58
			// srcs: (130, 6)(224) 3, (31) 2 --> (252) 6:PENB, ND0, *, PENB
			6'd6 : rdata = 41'b00011110111111100110000000000000100000000;
			// PEs: 57, 58 -> 57
			// srcs: (139, 7)(87) 2, (307) 6 --> (362) -4:NW0, PEGB2, -, NW0
			6'd7 : rdata = 41'b00010010000000001110000010000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 58) begin
	always @(*) begin
		case(address)
			// PEs: 58, 58 -> 57
			// srcs: (1, 0)(38) -2, (94) -1 --> (149) 2:ND0, NW0, *, PEGB1
			6'd0 : rdata = 41'b00011011000000000100000000000000010010000;
			// PEs: 57 -> 
			// srcs: (22, 1)(219) 2 --> (219) 2:PENB, pass, 
			6'd1 : rdata = 41'b11000110111111100000000000000000000000000;
			// PEs: 57, 58 -> 56
			// srcs: (29, 2)(217) 11, (219) 2 --> (220) 13:PENB, ALU, +, PEGB0
			6'd2 : rdata = 41'b00001110111111100011111111100000010000000;
			// PEs: 58, 57 -> 57
			// srcs: (133, 4)(3) 1, (252) 6 --> (307) 6:NM0, PENB, *, PEGB1
			6'd3 : rdata = 41'b00011100000000001101111111000000010010000;
			// PEs: 56, 58 -> 59
			// srcs: (140, 3)(224) 3, (38) -2 --> (259) -6:PEGB0, ND0, *, PENB
			6'd4 : rdata = 41'b00011111000000000110000000000000100000000;
			// PEs: 58, 59 -> 58
			// srcs: (149, 5)(94) -1, (314) -6 --> (369) 5:NW0, PEGB3, -, NW0
			6'd5 : rdata = 41'b00010010000000001110000011000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 59) begin
	always @(*) begin
		case(address)
			// PEs: 59, 59 -> 56
			// srcs: (1, 0)(45) 0, (101) -1 --> (156) 0:ND0, NW0, *, PEGB0
			6'd0 : rdata = 41'b00011011000000000100000000000000010000000;
			// PEs: 59, 58 -> 58
			// srcs: (143, 2)(3) 1, (259) -6 --> (314) -6:NM0, PENB, *, PEGB2
			6'd1 : rdata = 41'b00011100000000001101111111000000010100000;
			// PEs: 56, 59 -> 60
			// srcs: (147, 1)(224) 3, (45) 0 --> (266) 0:PEGB0, ND0, *, PENB
			6'd2 : rdata = 41'b00011111000000000110000000000000100000000;
			// PEs: 59, 60 -> 59
			// srcs: (156, 3)(101) -1, (321) 0 --> (376) -1:NW0, PEGB4, -, NW0
			6'd3 : rdata = 41'b00010010000000001110000100000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 60) begin
	always @(*) begin
		case(address)
			// PEs: 60, 60 -> 57
			// srcs: (1, 0)(52) 1, (108) 2 --> (163) 2:ND0, NW0, *, PEGB1
			6'd0 : rdata = 41'b00011011000000000100000000000000010010000;
			// PEs: 60, 59 -> 59
			// srcs: (150, 2)(3) 1, (266) 0 --> (321) 0:NM0, PENB, *, PEGB3
			6'd1 : rdata = 41'b00011100000000001101111111000000010110000;
			// PEs: 56, 60 -> 
			// srcs: (154, 1)(224) 3, (52) 1 --> (273) 3:PEGB0, ND0, *, 
			6'd2 : rdata = 41'b00011111000000000110000000000000000000000;
			// PEs: 60, 60 -> 
			// srcs: (157, 3)(3) 1, (273) 3 --> (328) 3:NM0, ALU, *, 
			6'd3 : rdata = 41'b00011100000000000011111111100000000000000;
			// PEs: 60, 60 -> 60
			// srcs: (160, 4)(108) 2, (328) 3 --> (383) -1:NW0, ALU, -, NW0
			6'd4 : rdata = 41'b00010010000000000011111111100100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 61) begin
	always @(*) begin
		case(address)
			// PEs: 61, 61 -> 57
			// srcs: (1, 0)(55) -2, (111) -1 --> (166) 2:ND0, NW0, *, PEGB1
			6'd0 : rdata = 41'b00011011000000000100000000000000010010000;
			// PEs: 56, 61 -> 
			// srcs: (157, 1)(224) 3, (55) -2 --> (276) -6:PEGB0, ND0, *, 
			6'd1 : rdata = 41'b00011111000000000110000000000000000000000;
			// PEs: 61, 61 -> 
			// srcs: (160, 2)(3) 1, (276) -6 --> (331) -6:NM0, ALU, *, 
			6'd2 : rdata = 41'b00011100000000000011111111100000000000000;
			// PEs: 61, 61 -> 61
			// srcs: (163, 3)(111) -1, (331) -6 --> (386) 5:NW0, ALU, -, NW0
			6'd3 : rdata = 41'b00010010000000000011111111100100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 62) begin
	always @(*) begin
		case(address)
			// PEs: 62, 62 -> 57
			// srcs: (1, 0)(58) 0, (114) 1 --> (169) 0:ND0, NW0, *, PEGB1
			6'd0 : rdata = 41'b00011011000000000100000000000000010010000;
			// PEs: 56, 62 -> 63
			// srcs: (159, 1)(224) 3, (58) 0 --> (279) 0:PEGB0, ND0, *, PENB
			6'd1 : rdata = 41'b00011111000000000110000000000000100000000;
			// PEs: 62, 63 -> 62
			// srcs: (168, 2)(114) 1, (334) 0 --> (389) 1:NW0, PEGB7, -, NW0
			6'd2 : rdata = 41'b00010010000000001110000111000100000000000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

if(peId == 63) begin
	always @(*) begin
		case(address)
			// PEs: 63, 62 -> 62
			// srcs: (162, 0)(3) 1, (279) 0 --> (334) 0:NM0, PENB, *, PEGB6
			6'd0 : rdata = 41'b00011100000000001101111111000000011100000;
			default : rdata = 41'b00000000000000000000000000000000000000000;
		endcase
	end
end

endgenerate
/*****************************************************************************/
endmodule
